magic
tech sky130A
magscale 1 2
timestamp 1667783412
<< metal1 >>
rect 102042 700748 102048 700800
rect 102100 700788 102106 700800
rect 105446 700788 105452 700800
rect 102100 700760 105452 700788
rect 102100 700748 102106 700760
rect 105446 700748 105452 700760
rect 105504 700748 105510 700800
rect 200022 700748 200028 700800
rect 200080 700788 200086 700800
rect 202782 700788 202788 700800
rect 200080 700760 202788 700788
rect 200080 700748 200086 700760
rect 202782 700748 202788 700760
rect 202840 700748 202846 700800
rect 314470 700748 314476 700800
rect 314528 700788 314534 700800
rect 316310 700788 316316 700800
rect 314528 700760 316316 700788
rect 314528 700748 314534 700760
rect 316310 700748 316316 700760
rect 316368 700748 316374 700800
rect 53006 700544 53012 700596
rect 53064 700584 53070 700596
rect 56778 700584 56784 700596
rect 53064 700556 56784 700584
rect 53064 700544 53070 700556
rect 56778 700544 56784 700556
rect 56836 700544 56842 700596
rect 151078 700544 151084 700596
rect 151136 700584 151142 700596
rect 154114 700584 154120 700596
rect 151136 700556 154120 700584
rect 151136 700544 151142 700556
rect 154114 700544 154120 700556
rect 154172 700544 154178 700596
rect 412450 700408 412456 700460
rect 412508 700448 412514 700460
rect 413646 700448 413652 700460
rect 412508 700420 413652 700448
rect 412508 700408 412514 700420
rect 413646 700408 413652 700420
rect 413704 700408 413710 700460
rect 363506 700340 363512 700392
rect 363564 700380 363570 700392
rect 364978 700380 364984 700392
rect 363564 700352 364984 700380
rect 363564 700340 363570 700352
rect 364978 700340 364984 700352
rect 365036 700340 365042 700392
rect 20346 700204 20352 700256
rect 20404 700244 20410 700256
rect 24302 700244 24308 700256
rect 20404 700216 24308 700244
rect 20404 700204 20410 700216
rect 24302 700204 24308 700216
rect 24360 700204 24366 700256
rect 36722 700204 36728 700256
rect 36780 700244 36786 700256
rect 40494 700244 40500 700256
rect 36780 700216 40500 700244
rect 36780 700204 36786 700216
rect 40494 700204 40500 700216
rect 40552 700204 40558 700256
rect 69382 700204 69388 700256
rect 69440 700244 69446 700256
rect 72970 700244 72976 700256
rect 69440 700216 72976 700244
rect 69440 700204 69446 700216
rect 72970 700204 72976 700216
rect 73028 700204 73034 700256
rect 85758 700204 85764 700256
rect 85816 700244 85822 700256
rect 89162 700244 89168 700256
rect 85816 700216 89168 700244
rect 85816 700204 85822 700216
rect 89162 700204 89168 700216
rect 89220 700204 89226 700256
rect 134702 700204 134708 700256
rect 134760 700244 134766 700256
rect 137830 700244 137836 700256
rect 134760 700216 137836 700244
rect 134760 700204 134766 700216
rect 137830 700204 137836 700216
rect 137888 700204 137894 700256
rect 167362 700204 167368 700256
rect 167420 700244 167426 700256
rect 170306 700244 170312 700256
rect 167420 700216 170312 700244
rect 167420 700204 167426 700216
rect 170306 700204 170312 700216
rect 170364 700204 170370 700256
rect 183738 700204 183744 700256
rect 183796 700244 183802 700256
rect 186498 700244 186504 700256
rect 183796 700216 186504 700244
rect 183796 700204 183802 700216
rect 186498 700204 186504 700216
rect 186556 700204 186562 700256
rect 232774 700204 232780 700256
rect 232832 700244 232838 700256
rect 235166 700244 235172 700256
rect 232832 700216 235172 700244
rect 232832 700204 232838 700216
rect 235166 700204 235172 700216
rect 235224 700204 235230 700256
rect 249058 700204 249064 700256
rect 249116 700244 249122 700256
rect 251450 700244 251456 700256
rect 249116 700216 251456 700244
rect 249116 700204 249122 700216
rect 251450 700204 251456 700216
rect 251508 700204 251514 700256
rect 265434 700204 265440 700256
rect 265492 700244 265498 700256
rect 267642 700244 267648 700256
rect 265492 700216 267648 700244
rect 265492 700204 265498 700216
rect 267642 700204 267648 700216
rect 267700 700204 267706 700256
rect 281810 700204 281816 700256
rect 281868 700244 281874 700256
rect 283834 700244 283840 700256
rect 281868 700216 283840 700244
rect 281868 700204 281874 700216
rect 283834 700204 283840 700216
rect 283892 700204 283898 700256
rect 330754 700204 330760 700256
rect 330812 700244 330818 700256
rect 332502 700244 332508 700256
rect 330812 700216 332508 700244
rect 330812 700204 330818 700216
rect 332502 700204 332508 700216
rect 332560 700204 332566 700256
rect 347130 700204 347136 700256
rect 347188 700244 347194 700256
rect 348786 700244 348792 700256
rect 347188 700216 348792 700244
rect 347188 700204 347194 700216
rect 348786 700204 348792 700216
rect 348844 700204 348850 700256
rect 396166 700204 396172 700256
rect 396224 700244 396230 700256
rect 397454 700244 397460 700256
rect 396224 700216 397460 700244
rect 396224 700204 396230 700216
rect 397454 700204 397460 700216
rect 397512 700204 397518 700256
rect 428826 700204 428832 700256
rect 428884 700244 428890 700256
rect 429838 700244 429844 700256
rect 428884 700216 429844 700244
rect 428884 700204 428890 700216
rect 429838 700204 429844 700216
rect 429896 700204 429902 700256
rect 445202 700204 445208 700256
rect 445260 700244 445266 700256
rect 446122 700244 446128 700256
rect 445260 700216 446128 700244
rect 445260 700204 445266 700216
rect 446122 700204 446128 700216
rect 446180 700204 446186 700256
rect 461486 700204 461492 700256
rect 461544 700244 461550 700256
rect 462314 700244 462320 700256
rect 461544 700216 462320 700244
rect 461544 700204 461550 700216
rect 462314 700204 462320 700216
rect 462372 700204 462378 700256
rect 118418 700136 118424 700188
rect 118476 700176 118482 700188
rect 121638 700176 121644 700188
rect 118476 700148 121644 700176
rect 118476 700136 118482 700148
rect 121638 700136 121644 700148
rect 121696 700136 121702 700188
rect 216398 700136 216404 700188
rect 216456 700176 216462 700188
rect 218974 700176 218980 700188
rect 216456 700148 218980 700176
rect 216456 700136 216462 700148
rect 218974 700136 218980 700148
rect 219032 700136 219038 700188
rect 298002 700136 298008 700188
rect 298060 700176 298066 700188
rect 300118 700176 300124 700188
rect 298060 700148 300124 700176
rect 298060 700136 298066 700148
rect 300118 700136 300124 700148
rect 300176 700136 300182 700188
rect 477862 700136 477868 700188
rect 477920 700176 477926 700188
rect 478506 700176 478512 700188
rect 477920 700148 478512 700176
rect 477920 700136 477926 700148
rect 478506 700136 478512 700148
rect 478564 700136 478570 700188
rect 494238 700136 494244 700188
rect 494296 700176 494302 700188
rect 494790 700176 494796 700188
rect 494296 700148 494796 700176
rect 494296 700136 494302 700148
rect 494790 700136 494796 700148
rect 494848 700136 494854 700188
rect 379790 699864 379796 699916
rect 379848 699904 379854 699916
rect 381170 699904 381176 699916
rect 379848 699876 381176 699904
rect 379848 699864 379854 699876
rect 381170 699864 381176 699876
rect 381228 699864 381234 699916
rect 576762 698232 576768 698284
rect 576820 698272 576826 698284
rect 580166 698272 580172 698284
rect 576820 698244 580172 698272
rect 576820 698232 576826 698244
rect 580166 698232 580172 698244
rect 580224 698232 580230 698284
rect 4014 698164 4020 698216
rect 4072 698204 4078 698216
rect 8110 698204 8116 698216
rect 4072 698176 8116 698204
rect 4072 698164 4078 698176
rect 8110 698164 8116 698176
rect 8168 698164 8174 698216
rect 578326 644512 578332 644564
rect 578384 644552 578390 644564
rect 580902 644552 580908 644564
rect 578384 644524 580908 644552
rect 578384 644512 578390 644524
rect 580902 644512 580908 644524
rect 580960 644512 580966 644564
rect 578878 257796 578884 257848
rect 578936 257836 578942 257848
rect 580902 257836 580908 257848
rect 578936 257808 580908 257836
rect 578936 257796 578942 257808
rect 580902 257796 580908 257808
rect 580960 257796 580966 257848
rect 578510 151444 578516 151496
rect 578568 151484 578574 151496
rect 580902 151484 580908 151496
rect 578568 151456 580908 151484
rect 578568 151444 578574 151456
rect 580902 151444 580908 151456
rect 580960 151444 580966 151496
rect 578326 44956 578332 45008
rect 578384 44996 578390 45008
rect 579982 44996 579988 45008
rect 578384 44968 579988 44996
rect 578384 44956 578390 44968
rect 579982 44956 579988 44968
rect 580040 44956 580046 45008
rect 576854 5516 576860 5568
rect 576912 5556 576918 5568
rect 579614 5556 579620 5568
rect 576912 5528 579620 5556
rect 576912 5516 576918 5528
rect 579614 5516 579620 5528
rect 579672 5516 579678 5568
rect 11146 3884 11152 3936
rect 11204 3924 11210 3936
rect 14502 3924 14508 3936
rect 11204 3896 14508 3924
rect 11204 3884 11210 3896
rect 14502 3884 14508 3896
rect 14560 3884 14566 3936
rect 14734 3884 14740 3936
rect 14792 3924 14798 3936
rect 17998 3924 18004 3936
rect 14792 3896 18004 3924
rect 14792 3884 14798 3896
rect 17998 3884 18004 3896
rect 18056 3884 18062 3936
rect 20622 3884 20628 3936
rect 20680 3924 20686 3936
rect 23794 3924 23800 3936
rect 20680 3896 23800 3924
rect 20680 3884 20686 3896
rect 23794 3884 23800 3896
rect 23852 3884 23858 3936
rect 24210 3884 24216 3936
rect 24268 3924 24274 3936
rect 27290 3924 27296 3936
rect 24268 3896 27296 3924
rect 24268 3884 24274 3896
rect 27290 3884 27296 3896
rect 27348 3884 27354 3936
rect 27706 3884 27712 3936
rect 27764 3924 27770 3936
rect 30694 3924 30700 3936
rect 27764 3896 30700 3924
rect 27764 3884 27770 3896
rect 30694 3884 30700 3896
rect 30752 3884 30758 3936
rect 32398 3884 32404 3936
rect 32456 3924 32462 3936
rect 35386 3924 35392 3936
rect 32456 3896 35392 3924
rect 32456 3884 32462 3896
rect 35386 3884 35392 3896
rect 35444 3884 35450 3936
rect 38378 3884 38384 3936
rect 38436 3924 38442 3936
rect 41182 3924 41188 3936
rect 38436 3896 41188 3924
rect 38436 3884 38442 3896
rect 41182 3884 41188 3896
rect 41240 3884 41246 3936
rect 43070 3884 43076 3936
rect 43128 3924 43134 3936
rect 45782 3924 45788 3936
rect 43128 3896 45788 3924
rect 43128 3884 43134 3896
rect 45782 3884 45788 3896
rect 45840 3884 45846 3936
rect 46658 3884 46664 3936
rect 46716 3924 46722 3936
rect 49278 3924 49284 3936
rect 46716 3896 49284 3924
rect 46716 3884 46722 3896
rect 49278 3884 49284 3896
rect 49336 3884 49342 3936
rect 50154 3884 50160 3936
rect 50212 3924 50218 3936
rect 52774 3924 52780 3936
rect 50212 3896 52780 3924
rect 50212 3884 50218 3896
rect 52774 3884 52780 3896
rect 52832 3884 52838 3936
rect 56042 3884 56048 3936
rect 56100 3924 56106 3936
rect 58570 3924 58576 3936
rect 56100 3896 58576 3924
rect 56100 3884 56106 3896
rect 58570 3884 58576 3896
rect 58628 3884 58634 3936
rect 72602 3884 72608 3936
rect 72660 3924 72666 3936
rect 74854 3924 74860 3936
rect 72660 3896 74860 3924
rect 72660 3884 72666 3896
rect 74854 3884 74860 3896
rect 74912 3884 74918 3936
rect 247630 3884 247636 3936
rect 247688 3924 247694 3936
rect 248598 3924 248604 3936
rect 247688 3896 248604 3924
rect 247688 3884 247694 3896
rect 248598 3884 248604 3896
rect 248656 3884 248662 3936
rect 285902 3884 285908 3936
rect 285960 3924 285966 3936
rect 287790 3924 287796 3936
rect 285960 3896 287796 3924
rect 285960 3884 285966 3896
rect 287790 3884 287796 3896
rect 287848 3884 287854 3936
rect 1670 3816 1676 3868
rect 1728 3856 1734 3868
rect 5210 3856 5216 3868
rect 1728 3828 5216 3856
rect 1728 3816 1734 3828
rect 5210 3816 5216 3828
rect 5268 3816 5274 3868
rect 13538 3816 13544 3868
rect 13596 3856 13602 3868
rect 16802 3856 16808 3868
rect 13596 3828 16808 3856
rect 13596 3816 13602 3828
rect 16802 3816 16808 3828
rect 16860 3816 16866 3868
rect 19426 3816 19432 3868
rect 19484 3856 19490 3868
rect 22598 3856 22604 3868
rect 19484 3828 22604 3856
rect 19484 3816 19490 3828
rect 22598 3816 22604 3828
rect 22656 3816 22662 3868
rect 23014 3816 23020 3868
rect 23072 3856 23078 3868
rect 26094 3856 26100 3868
rect 23072 3828 26100 3856
rect 23072 3816 23078 3828
rect 26094 3816 26100 3828
rect 26152 3816 26158 3868
rect 26510 3816 26516 3868
rect 26568 3856 26574 3868
rect 29590 3856 29596 3868
rect 26568 3828 29596 3856
rect 26568 3816 26574 3828
rect 29590 3816 29596 3828
rect 29648 3816 29654 3868
rect 30098 3816 30104 3868
rect 30156 3856 30162 3868
rect 33086 3856 33092 3868
rect 30156 3828 33092 3856
rect 30156 3816 30162 3828
rect 33086 3816 33092 3828
rect 33144 3816 33150 3868
rect 33594 3816 33600 3868
rect 33652 3856 33658 3868
rect 36582 3856 36588 3868
rect 33652 3828 36588 3856
rect 33652 3816 33658 3828
rect 36582 3816 36588 3828
rect 36640 3816 36646 3868
rect 37182 3816 37188 3868
rect 37240 3856 37246 3868
rect 39986 3856 39992 3868
rect 37240 3828 39992 3856
rect 37240 3816 37246 3828
rect 39986 3816 39992 3828
rect 40044 3816 40050 3868
rect 41874 3816 41880 3868
rect 41932 3856 41938 3868
rect 44678 3856 44684 3868
rect 41932 3828 44684 3856
rect 41932 3816 41938 3828
rect 44678 3816 44684 3828
rect 44736 3816 44742 3868
rect 45462 3816 45468 3868
rect 45520 3856 45526 3868
rect 48174 3856 48180 3868
rect 45520 3828 48180 3856
rect 45520 3816 45526 3828
rect 48174 3816 48180 3828
rect 48232 3816 48238 3868
rect 48958 3816 48964 3868
rect 49016 3856 49022 3868
rect 51578 3856 51584 3868
rect 49016 3828 51584 3856
rect 49016 3816 49022 3828
rect 51578 3816 51584 3828
rect 51636 3816 51642 3868
rect 53742 3816 53748 3868
rect 53800 3856 53806 3868
rect 56270 3856 56276 3868
rect 53800 3828 56276 3856
rect 53800 3816 53806 3828
rect 56270 3816 56276 3828
rect 56328 3816 56334 3868
rect 57238 3816 57244 3868
rect 57296 3856 57302 3868
rect 59766 3856 59772 3868
rect 57296 3828 59772 3856
rect 57296 3816 57302 3828
rect 59766 3816 59772 3828
rect 59824 3816 59830 3868
rect 71498 3816 71504 3868
rect 71556 3856 71562 3868
rect 73658 3856 73664 3868
rect 71556 3828 73664 3856
rect 71556 3816 71562 3828
rect 73658 3816 73664 3828
rect 73716 3816 73722 3868
rect 78582 3816 78588 3868
rect 78640 3856 78646 3868
rect 80650 3856 80656 3868
rect 78640 3828 80656 3856
rect 78640 3816 78646 3828
rect 80650 3816 80656 3828
rect 80708 3816 80714 3868
rect 80882 3816 80888 3868
rect 80940 3856 80946 3868
rect 82950 3856 82956 3868
rect 80940 3828 82956 3856
rect 80940 3816 80946 3828
rect 82950 3816 82956 3828
rect 83008 3816 83014 3868
rect 87966 3816 87972 3868
rect 88024 3856 88030 3868
rect 89942 3856 89948 3868
rect 88024 3828 89948 3856
rect 88024 3816 88030 3828
rect 89942 3816 89948 3828
rect 90000 3816 90006 3868
rect 96246 3816 96252 3868
rect 96304 3856 96310 3868
rect 98038 3856 98044 3868
rect 96304 3828 98044 3856
rect 96304 3816 96310 3828
rect 98038 3816 98044 3828
rect 98096 3816 98102 3868
rect 244134 3816 244140 3868
rect 244192 3856 244198 3868
rect 245194 3856 245200 3868
rect 244192 3828 245200 3856
rect 244192 3816 244198 3828
rect 245194 3816 245200 3828
rect 245252 3816 245258 3868
rect 256922 3816 256928 3868
rect 256980 3856 256986 3868
rect 258258 3856 258264 3868
rect 256980 3828 258264 3856
rect 256980 3816 256986 3828
rect 258258 3816 258264 3828
rect 258316 3816 258322 3868
rect 259222 3816 259228 3868
rect 259280 3856 259286 3868
rect 260650 3856 260656 3868
rect 259280 3828 260656 3856
rect 259280 3816 259286 3828
rect 260650 3816 260656 3828
rect 260708 3816 260714 3868
rect 261614 3816 261620 3868
rect 261672 3856 261678 3868
rect 262950 3856 262956 3868
rect 261672 3828 262956 3856
rect 261672 3816 261678 3828
rect 262950 3816 262956 3828
rect 263008 3816 263014 3868
rect 263914 3816 263920 3868
rect 263972 3856 263978 3868
rect 265342 3856 265348 3868
rect 263972 3828 265348 3856
rect 263972 3816 263978 3828
rect 265342 3816 265348 3828
rect 265400 3816 265406 3868
rect 268514 3816 268520 3868
rect 268572 3856 268578 3868
rect 270034 3856 270040 3868
rect 268572 3828 270040 3856
rect 268572 3816 268578 3828
rect 270034 3816 270040 3828
rect 270092 3816 270098 3868
rect 270814 3816 270820 3868
rect 270872 3856 270878 3868
rect 272426 3856 272432 3868
rect 270872 3828 272432 3856
rect 270872 3816 270878 3828
rect 272426 3816 272432 3828
rect 272484 3816 272490 3868
rect 275506 3816 275512 3868
rect 275564 3856 275570 3868
rect 277118 3856 277124 3868
rect 275564 3828 277124 3856
rect 275564 3816 275570 3828
rect 277118 3816 277124 3828
rect 277176 3816 277182 3868
rect 277806 3816 277812 3868
rect 277864 3856 277870 3868
rect 279510 3856 279516 3868
rect 277864 3828 279516 3856
rect 277864 3816 277870 3828
rect 279510 3816 279516 3828
rect 279568 3816 279574 3868
rect 284798 3816 284804 3868
rect 284856 3856 284862 3868
rect 286594 3856 286600 3868
rect 284856 3828 286600 3856
rect 284856 3816 284862 3828
rect 286594 3816 286600 3828
rect 286652 3816 286658 3868
rect 292894 3816 292900 3868
rect 292952 3856 292958 3868
rect 294874 3856 294880 3868
rect 292952 3828 294880 3856
rect 292952 3816 292958 3828
rect 294874 3816 294880 3828
rect 294932 3816 294938 3868
rect 299886 3816 299892 3868
rect 299944 3856 299950 3868
rect 301958 3856 301964 3868
rect 299944 3828 301964 3856
rect 299944 3816 299950 3828
rect 301958 3816 301964 3828
rect 302016 3816 302022 3868
rect 306786 3816 306792 3868
rect 306844 3856 306850 3868
rect 309042 3856 309048 3868
rect 306844 3828 309048 3856
rect 306844 3816 306850 3828
rect 309042 3816 309048 3828
rect 309100 3816 309106 3868
rect 566 3748 572 3800
rect 624 3788 630 3800
rect 4106 3788 4112 3800
rect 624 3760 4112 3788
rect 624 3748 630 3760
rect 4106 3748 4112 3760
rect 4164 3748 4170 3800
rect 7650 3748 7656 3800
rect 7708 3788 7714 3800
rect 11006 3788 11012 3800
rect 7708 3760 11012 3788
rect 7708 3748 7714 3760
rect 11006 3748 11012 3760
rect 11064 3748 11070 3800
rect 12342 3748 12348 3800
rect 12400 3788 12406 3800
rect 15698 3788 15704 3800
rect 12400 3760 15704 3788
rect 12400 3748 12406 3760
rect 15698 3748 15704 3760
rect 15756 3748 15762 3800
rect 15930 3748 15936 3800
rect 15988 3788 15994 3800
rect 19102 3788 19108 3800
rect 15988 3760 19108 3788
rect 15988 3748 15994 3760
rect 19102 3748 19108 3760
rect 19160 3748 19166 3800
rect 21818 3748 21824 3800
rect 21876 3788 21882 3800
rect 24898 3788 24904 3800
rect 21876 3760 24904 3788
rect 21876 3748 21882 3760
rect 24898 3748 24904 3760
rect 24956 3748 24962 3800
rect 25314 3748 25320 3800
rect 25372 3788 25378 3800
rect 28394 3788 28400 3800
rect 25372 3760 28400 3788
rect 25372 3748 25378 3760
rect 28394 3748 28400 3760
rect 28452 3748 28458 3800
rect 31294 3748 31300 3800
rect 31352 3788 31358 3800
rect 34190 3788 34196 3800
rect 31352 3760 34196 3788
rect 31352 3748 31358 3760
rect 34190 3748 34196 3760
rect 34248 3748 34254 3800
rect 34790 3748 34796 3800
rect 34848 3788 34854 3800
rect 37686 3788 37692 3800
rect 34848 3760 37692 3788
rect 34848 3748 34854 3760
rect 37686 3748 37692 3760
rect 37744 3748 37750 3800
rect 40678 3748 40684 3800
rect 40736 3788 40742 3800
rect 43482 3788 43488 3800
rect 40736 3760 43488 3788
rect 40736 3748 40742 3760
rect 43482 3748 43488 3760
rect 43540 3748 43546 3800
rect 44266 3748 44272 3800
rect 44324 3788 44330 3800
rect 46978 3788 46984 3800
rect 44324 3760 46984 3788
rect 44324 3748 44330 3760
rect 46978 3748 46984 3760
rect 47036 3748 47042 3800
rect 47854 3748 47860 3800
rect 47912 3788 47918 3800
rect 50474 3788 50480 3800
rect 47912 3760 50480 3788
rect 47912 3748 47918 3760
rect 50474 3748 50480 3760
rect 50532 3748 50538 3800
rect 51350 3748 51356 3800
rect 51408 3788 51414 3800
rect 53970 3788 53976 3800
rect 51408 3760 53976 3788
rect 51408 3748 51414 3760
rect 53970 3748 53976 3760
rect 54028 3748 54034 3800
rect 54938 3748 54944 3800
rect 54996 3788 55002 3800
rect 57374 3788 57380 3800
rect 54996 3760 57380 3788
rect 54996 3748 55002 3760
rect 57374 3748 57380 3760
rect 57432 3748 57438 3800
rect 58434 3748 58440 3800
rect 58492 3788 58498 3800
rect 60870 3788 60876 3800
rect 58492 3760 60876 3788
rect 58492 3748 58498 3760
rect 60870 3748 60876 3760
rect 60928 3748 60934 3800
rect 64322 3748 64328 3800
rect 64380 3788 64386 3800
rect 66666 3788 66672 3800
rect 64380 3760 66672 3788
rect 64380 3748 64386 3760
rect 66666 3748 66672 3760
rect 66724 3748 66730 3800
rect 67082 3748 67088 3800
rect 67140 3788 67146 3800
rect 69058 3788 69064 3800
rect 67140 3760 69064 3788
rect 67140 3748 67146 3760
rect 69058 3748 69064 3760
rect 69116 3748 69122 3800
rect 70302 3748 70308 3800
rect 70360 3788 70366 3800
rect 72462 3788 72468 3800
rect 70360 3760 72468 3788
rect 70360 3748 70366 3760
rect 72462 3748 72468 3760
rect 72520 3748 72526 3800
rect 73798 3748 73804 3800
rect 73856 3788 73862 3800
rect 75958 3788 75964 3800
rect 73856 3760 75964 3788
rect 73856 3748 73862 3760
rect 75958 3748 75964 3760
rect 76016 3748 76022 3800
rect 79686 3748 79692 3800
rect 79744 3788 79750 3800
rect 81754 3788 81760 3800
rect 79744 3760 81760 3788
rect 79744 3748 79750 3760
rect 81754 3748 81760 3760
rect 81812 3748 81818 3800
rect 86862 3748 86868 3800
rect 86920 3788 86926 3800
rect 88746 3788 88752 3800
rect 86920 3760 88752 3788
rect 86920 3748 86926 3760
rect 88746 3748 88752 3760
rect 88804 3748 88810 3800
rect 95142 3748 95148 3800
rect 95200 3788 95206 3800
rect 96842 3788 96848 3800
rect 95200 3760 96848 3788
rect 95200 3748 95206 3760
rect 96842 3748 96848 3760
rect 96900 3748 96906 3800
rect 103330 3748 103336 3800
rect 103388 3788 103394 3800
rect 104938 3788 104944 3800
rect 103388 3760 104944 3788
rect 103388 3748 103394 3760
rect 104938 3748 104944 3760
rect 104996 3748 105002 3800
rect 216350 3748 216356 3800
rect 216408 3788 216414 3800
rect 216858 3788 216864 3800
rect 216408 3760 216864 3788
rect 216408 3748 216414 3760
rect 216858 3748 216864 3760
rect 216916 3748 216922 3800
rect 222146 3748 222152 3800
rect 222204 3788 222210 3800
rect 222746 3788 222752 3800
rect 222204 3760 222752 3788
rect 222204 3748 222210 3760
rect 222746 3748 222752 3760
rect 222804 3748 222810 3800
rect 224446 3748 224452 3800
rect 224504 3788 224510 3800
rect 225138 3788 225144 3800
rect 224504 3760 225144 3788
rect 224504 3748 224510 3760
rect 225138 3748 225144 3760
rect 225196 3748 225202 3800
rect 230242 3748 230248 3800
rect 230300 3788 230306 3800
rect 231026 3788 231032 3800
rect 230300 3760 231032 3788
rect 230300 3748 230306 3760
rect 231026 3748 231032 3760
rect 231084 3748 231090 3800
rect 231438 3748 231444 3800
rect 231496 3788 231502 3800
rect 232222 3788 232228 3800
rect 231496 3760 232228 3788
rect 231496 3748 231502 3760
rect 232222 3748 232228 3760
rect 232280 3748 232286 3800
rect 232542 3748 232548 3800
rect 232600 3788 232606 3800
rect 233418 3788 233424 3800
rect 232600 3760 233424 3788
rect 232600 3748 232606 3760
rect 233418 3748 233424 3760
rect 233476 3748 233482 3800
rect 233738 3748 233744 3800
rect 233796 3788 233802 3800
rect 234614 3788 234620 3800
rect 233796 3760 234620 3788
rect 233796 3748 233802 3760
rect 234614 3748 234620 3760
rect 234672 3748 234678 3800
rect 237234 3748 237240 3800
rect 237292 3788 237298 3800
rect 238110 3788 238116 3800
rect 237292 3760 238116 3788
rect 237292 3748 237298 3760
rect 238110 3748 238116 3760
rect 238168 3748 238174 3800
rect 238338 3748 238344 3800
rect 238396 3788 238402 3800
rect 239306 3788 239312 3800
rect 238396 3760 239312 3788
rect 238396 3748 238402 3760
rect 239306 3748 239312 3760
rect 239364 3748 239370 3800
rect 239534 3748 239540 3800
rect 239592 3788 239598 3800
rect 240502 3788 240508 3800
rect 239592 3760 240508 3788
rect 239592 3748 239598 3760
rect 240502 3748 240508 3760
rect 240560 3748 240566 3800
rect 240730 3748 240736 3800
rect 240788 3788 240794 3800
rect 241698 3788 241704 3800
rect 240788 3760 241704 3788
rect 240788 3748 240794 3760
rect 241698 3748 241704 3760
rect 241756 3748 241762 3800
rect 241834 3748 241840 3800
rect 241892 3788 241898 3800
rect 242894 3788 242900 3800
rect 241892 3760 242900 3788
rect 241892 3748 241898 3760
rect 242894 3748 242900 3760
rect 242952 3748 242958 3800
rect 245330 3748 245336 3800
rect 245388 3788 245394 3800
rect 246390 3788 246396 3800
rect 245388 3760 246396 3788
rect 245388 3748 245394 3760
rect 246390 3748 246396 3760
rect 246448 3748 246454 3800
rect 246526 3748 246532 3800
rect 246584 3788 246590 3800
rect 247586 3788 247592 3800
rect 246584 3760 247592 3788
rect 246584 3748 246590 3760
rect 247586 3748 247592 3760
rect 247644 3748 247650 3800
rect 250022 3748 250028 3800
rect 250080 3788 250086 3800
rect 251174 3788 251180 3800
rect 250080 3760 251180 3788
rect 250080 3748 250086 3760
rect 251174 3748 251180 3760
rect 251232 3748 251238 3800
rect 252322 3748 252328 3800
rect 252380 3788 252386 3800
rect 253474 3788 253480 3800
rect 252380 3760 253480 3788
rect 252380 3748 252386 3760
rect 253474 3748 253480 3760
rect 253532 3748 253538 3800
rect 255818 3748 255824 3800
rect 255876 3788 255882 3800
rect 257062 3788 257068 3800
rect 255876 3760 257068 3788
rect 255876 3748 255882 3760
rect 257062 3748 257068 3760
rect 257120 3748 257126 3800
rect 258118 3748 258124 3800
rect 258176 3788 258182 3800
rect 259454 3788 259460 3800
rect 258176 3760 259460 3788
rect 258176 3748 258182 3760
rect 259454 3748 259460 3760
rect 259512 3748 259518 3800
rect 260418 3748 260424 3800
rect 260476 3788 260482 3800
rect 261754 3788 261760 3800
rect 260476 3760 261760 3788
rect 260476 3748 260482 3760
rect 261754 3748 261760 3760
rect 261812 3748 261818 3800
rect 262718 3748 262724 3800
rect 262776 3788 262782 3800
rect 264146 3788 264152 3800
rect 262776 3760 264152 3788
rect 262776 3748 262782 3760
rect 264146 3748 264152 3760
rect 264204 3748 264210 3800
rect 265018 3748 265024 3800
rect 265076 3788 265082 3800
rect 266538 3788 266544 3800
rect 265076 3760 266544 3788
rect 265076 3748 265082 3760
rect 266538 3748 266544 3760
rect 266596 3748 266602 3800
rect 267410 3748 267416 3800
rect 267468 3788 267474 3800
rect 268838 3788 268844 3800
rect 267468 3760 268844 3788
rect 267468 3748 267474 3760
rect 268838 3748 268844 3760
rect 268896 3748 268902 3800
rect 269710 3748 269716 3800
rect 269768 3788 269774 3800
rect 271230 3788 271236 3800
rect 269768 3760 271236 3788
rect 269768 3748 269774 3760
rect 271230 3748 271236 3760
rect 271288 3748 271294 3800
rect 272010 3748 272016 3800
rect 272068 3788 272074 3800
rect 273622 3788 273628 3800
rect 272068 3760 273628 3788
rect 272068 3748 272074 3760
rect 273622 3748 273628 3760
rect 273680 3748 273686 3800
rect 276702 3748 276708 3800
rect 276760 3788 276766 3800
rect 278314 3788 278320 3800
rect 276760 3760 278320 3788
rect 276760 3748 276766 3760
rect 278314 3748 278320 3760
rect 278372 3748 278378 3800
rect 279002 3748 279008 3800
rect 279060 3788 279066 3800
rect 280706 3788 280712 3800
rect 279060 3760 280712 3788
rect 279060 3748 279066 3760
rect 280706 3748 280712 3760
rect 280764 3748 280770 3800
rect 283602 3748 283608 3800
rect 283660 3788 283666 3800
rect 285398 3788 285404 3800
rect 283660 3760 285404 3788
rect 283660 3748 283666 3760
rect 285398 3748 285404 3760
rect 285456 3748 285462 3800
rect 287098 3748 287104 3800
rect 287156 3788 287162 3800
rect 288986 3788 288992 3800
rect 287156 3760 288992 3788
rect 287156 3748 287162 3760
rect 288986 3748 288992 3760
rect 289044 3748 289050 3800
rect 291698 3748 291704 3800
rect 291756 3788 291762 3800
rect 293678 3788 293684 3800
rect 291756 3760 293684 3788
rect 291756 3748 291762 3760
rect 293678 3748 293684 3760
rect 293736 3748 293742 3800
rect 294090 3748 294096 3800
rect 294148 3788 294154 3800
rect 296070 3788 296076 3800
rect 294148 3760 296076 3788
rect 294148 3748 294154 3760
rect 296070 3748 296076 3760
rect 296128 3748 296134 3800
rect 298690 3748 298696 3800
rect 298748 3788 298754 3800
rect 300762 3788 300768 3800
rect 298748 3760 300768 3788
rect 298748 3748 298754 3760
rect 300762 3748 300768 3760
rect 300820 3748 300826 3800
rect 300990 3748 300996 3800
rect 301048 3788 301054 3800
rect 303154 3788 303160 3800
rect 301048 3760 303160 3788
rect 301048 3748 301054 3760
rect 303154 3748 303160 3760
rect 303212 3748 303218 3800
rect 307982 3748 307988 3800
rect 308040 3788 308046 3800
rect 310238 3788 310244 3800
rect 308040 3760 310244 3788
rect 308040 3748 308046 3760
rect 310238 3748 310244 3760
rect 310296 3748 310302 3800
rect 316078 3748 316084 3800
rect 316136 3788 316142 3800
rect 318518 3788 318524 3800
rect 316136 3760 318524 3788
rect 316136 3748 316142 3760
rect 318518 3748 318524 3760
rect 318576 3748 318582 3800
rect 323070 3748 323076 3800
rect 323128 3788 323134 3800
rect 325602 3788 325608 3800
rect 323128 3760 325608 3788
rect 323128 3748 323134 3760
rect 325602 3748 325608 3760
rect 325660 3748 325666 3800
rect 6454 3000 6460 3052
rect 6512 3040 6518 3052
rect 9858 3040 9864 3052
rect 6512 3012 9864 3040
rect 6512 3000 6518 3012
rect 9858 3000 9864 3012
rect 9916 3000 9922 3052
rect 63218 3000 63224 3052
rect 63276 3040 63282 3052
rect 65518 3040 65524 3052
rect 63276 3012 65524 3040
rect 63276 3000 63282 3012
rect 65518 3000 65524 3012
rect 65576 3000 65582 3052
rect 18230 2864 18236 2916
rect 18288 2904 18294 2916
rect 21450 2904 21456 2916
rect 18288 2876 21456 2904
rect 18288 2864 18294 2876
rect 21450 2864 21456 2876
rect 21508 2864 21514 2916
rect 253382 2864 253388 2916
rect 253440 2904 253446 2916
rect 254670 2904 254676 2916
rect 253440 2876 254676 2904
rect 253440 2864 253446 2876
rect 254670 2864 254676 2876
rect 254728 2864 254734 2916
rect 4062 2796 4068 2848
rect 4120 2836 4126 2848
rect 7466 2836 7472 2848
rect 4120 2808 7472 2836
rect 4120 2796 4126 2808
rect 7466 2796 7472 2808
rect 7524 2796 7530 2848
rect 9950 2796 9956 2848
rect 10008 2836 10014 2848
rect 13262 2836 13268 2848
rect 10008 2808 13268 2836
rect 10008 2796 10014 2808
rect 13262 2796 13268 2808
rect 13320 2796 13326 2848
rect 17034 2796 17040 2848
rect 17092 2836 17098 2848
rect 20254 2836 20260 2848
rect 17092 2808 20260 2836
rect 17092 2796 17098 2808
rect 20254 2796 20260 2808
rect 20312 2796 20318 2848
rect 28902 2796 28908 2848
rect 28960 2836 28966 2848
rect 31846 2836 31852 2848
rect 28960 2808 31852 2836
rect 28960 2796 28966 2808
rect 31846 2796 31852 2808
rect 31904 2796 31910 2848
rect 35986 2796 35992 2848
rect 36044 2836 36050 2848
rect 38838 2836 38844 2848
rect 36044 2808 38844 2836
rect 36044 2796 36050 2808
rect 38838 2796 38844 2808
rect 38896 2796 38902 2848
rect 39574 2796 39580 2848
rect 39632 2836 39638 2848
rect 42334 2836 42340 2848
rect 39632 2808 42340 2836
rect 39632 2796 39638 2808
rect 42334 2796 42340 2808
rect 42392 2796 42398 2848
rect 62022 2796 62028 2848
rect 62080 2836 62086 2848
rect 64414 2836 64420 2848
rect 62080 2808 64420 2836
rect 62080 2796 62086 2808
rect 64414 2796 64420 2808
rect 64472 2796 64478 2848
rect 65518 2796 65524 2848
rect 65576 2836 65582 2848
rect 67818 2836 67824 2848
rect 65576 2808 67824 2836
rect 65576 2796 65582 2808
rect 67818 2796 67824 2808
rect 67876 2796 67882 2848
rect 248874 2796 248880 2848
rect 248932 2836 248938 2848
rect 249978 2836 249984 2848
rect 248932 2808 249984 2836
rect 248932 2796 248938 2808
rect 249978 2796 249984 2808
rect 250036 2796 250042 2848
rect 251082 2796 251088 2848
rect 251140 2836 251146 2848
rect 252370 2836 252376 2848
rect 251140 2808 252376 2836
rect 251140 2796 251146 2808
rect 252370 2796 252376 2808
rect 252428 2796 252434 2848
rect 254578 2796 254584 2848
rect 254636 2836 254642 2848
rect 255866 2836 255872 2848
rect 254636 2808 255872 2836
rect 254636 2796 254642 2808
rect 255866 2796 255872 2808
rect 255924 2796 255930 2848
rect 309226 2796 309232 2848
rect 309284 2836 309290 2848
rect 311434 2836 311440 2848
rect 309284 2808 311440 2836
rect 309284 2796 309290 2808
rect 311434 2796 311440 2808
rect 311492 2796 311498 2848
rect 315022 2796 315028 2848
rect 315080 2836 315086 2848
rect 317322 2836 317328 2848
rect 315080 2808 317328 2836
rect 315080 2796 315086 2808
rect 317322 2796 317328 2808
rect 317380 2796 317386 2848
rect 411162 2796 411168 2848
rect 411220 2836 411226 2848
rect 415486 2836 415492 2848
rect 411220 2808 415492 2836
rect 411220 2796 411226 2808
rect 415486 2796 415492 2808
rect 415544 2796 415550 2848
rect 440142 2796 440148 2848
rect 440200 2836 440206 2848
rect 445018 2836 445024 2848
rect 440200 2808 445024 2836
rect 440200 2796 440206 2808
rect 445018 2796 445024 2808
rect 445076 2796 445082 2848
rect 449526 2796 449532 2848
rect 449584 2836 449590 2848
rect 454494 2836 454500 2848
rect 449584 2808 454500 2836
rect 449584 2796 449590 2808
rect 454494 2796 454500 2808
rect 454552 2796 454558 2848
rect 478506 2796 478512 2848
rect 478564 2836 478570 2848
rect 484026 2836 484032 2848
rect 478564 2808 484032 2836
rect 478564 2796 478570 2808
rect 484026 2796 484032 2808
rect 484084 2796 484090 2848
rect 3234 1300 3240 1352
rect 3292 1340 3298 1352
rect 6362 1340 6368 1352
rect 3292 1312 6368 1340
rect 3292 1300 3298 1312
rect 6362 1300 6368 1312
rect 6420 1300 6426 1352
rect 60826 1300 60832 1352
rect 60884 1340 60890 1352
rect 63310 1340 63316 1352
rect 60884 1312 63316 1340
rect 60884 1300 60890 1312
rect 63310 1300 63316 1312
rect 63368 1300 63374 1352
rect 67910 1300 67916 1352
rect 67968 1340 67974 1352
rect 70118 1340 70124 1352
rect 67968 1312 70124 1340
rect 67968 1300 67974 1312
rect 70118 1300 70124 1312
rect 70176 1300 70182 1352
rect 76190 1300 76196 1352
rect 76248 1340 76254 1352
rect 78214 1340 78220 1352
rect 76248 1312 78220 1340
rect 76248 1300 76254 1312
rect 78214 1300 78220 1312
rect 78272 1300 78278 1352
rect 83274 1300 83280 1352
rect 83332 1340 83338 1352
rect 85206 1340 85212 1352
rect 83332 1312 85212 1340
rect 83332 1300 83338 1312
rect 85206 1300 85212 1312
rect 85264 1300 85270 1352
rect 85666 1300 85672 1352
rect 85724 1340 85730 1352
rect 87506 1340 87512 1352
rect 85724 1312 87512 1340
rect 85724 1300 85730 1312
rect 87506 1300 87512 1312
rect 87564 1300 87570 1352
rect 89162 1300 89168 1352
rect 89220 1340 89226 1352
rect 91002 1340 91008 1352
rect 89220 1312 91008 1340
rect 89220 1300 89226 1312
rect 91002 1300 91008 1312
rect 91060 1300 91066 1352
rect 91554 1300 91560 1352
rect 91612 1340 91618 1352
rect 93302 1340 93308 1352
rect 91612 1312 93308 1340
rect 91612 1300 91618 1312
rect 93302 1300 93308 1312
rect 93360 1300 93366 1352
rect 93946 1300 93952 1352
rect 94004 1340 94010 1352
rect 95694 1340 95700 1352
rect 94004 1312 95700 1340
rect 94004 1300 94010 1312
rect 95694 1300 95700 1312
rect 95752 1300 95758 1352
rect 97442 1300 97448 1352
rect 97500 1340 97506 1352
rect 99098 1340 99104 1352
rect 97500 1312 99104 1340
rect 97500 1300 97506 1312
rect 99098 1300 99104 1312
rect 99156 1300 99162 1352
rect 101030 1300 101036 1352
rect 101088 1340 101094 1352
rect 102594 1340 102600 1352
rect 101088 1312 102600 1340
rect 101088 1300 101094 1312
rect 102594 1300 102600 1312
rect 102652 1300 102658 1352
rect 104526 1300 104532 1352
rect 104584 1340 104590 1352
rect 106090 1340 106096 1352
rect 104584 1312 106096 1340
rect 104584 1300 104590 1312
rect 106090 1300 106096 1312
rect 106148 1300 106154 1352
rect 106918 1300 106924 1352
rect 106976 1340 106982 1352
rect 108390 1340 108396 1352
rect 106976 1312 108396 1340
rect 106976 1300 106982 1312
rect 108390 1300 108396 1312
rect 108448 1300 108454 1352
rect 109310 1300 109316 1352
rect 109368 1340 109374 1352
rect 110690 1340 110696 1352
rect 109368 1312 110696 1340
rect 109368 1300 109374 1312
rect 110690 1300 110696 1312
rect 110748 1300 110754 1352
rect 112806 1300 112812 1352
rect 112864 1340 112870 1352
rect 114186 1340 114192 1352
rect 112864 1312 114192 1340
rect 112864 1300 112870 1312
rect 114186 1300 114192 1312
rect 114244 1300 114250 1352
rect 116394 1300 116400 1352
rect 116452 1340 116458 1352
rect 117682 1340 117688 1352
rect 116452 1312 117688 1340
rect 116452 1300 116458 1312
rect 117682 1300 117688 1312
rect 117740 1300 117746 1352
rect 119890 1300 119896 1352
rect 119948 1340 119954 1352
rect 121178 1340 121184 1352
rect 119948 1312 121184 1340
rect 119948 1300 119954 1312
rect 121178 1300 121184 1312
rect 121236 1300 121242 1352
rect 125870 1300 125876 1352
rect 125928 1340 125934 1352
rect 126974 1340 126980 1352
rect 125928 1312 126980 1340
rect 125928 1300 125934 1312
rect 126974 1300 126980 1312
rect 127032 1300 127038 1352
rect 129366 1300 129372 1352
rect 129424 1340 129430 1352
rect 130470 1340 130476 1352
rect 129424 1312 130476 1340
rect 129424 1300 129430 1312
rect 130470 1300 130476 1312
rect 130528 1300 130534 1352
rect 130562 1300 130568 1352
rect 130620 1340 130626 1352
rect 131574 1340 131580 1352
rect 130620 1312 131580 1340
rect 130620 1300 130626 1312
rect 131574 1300 131580 1312
rect 131632 1300 131638 1352
rect 131758 1300 131764 1352
rect 131816 1340 131822 1352
rect 132770 1340 132776 1352
rect 131816 1312 132776 1340
rect 131816 1300 131822 1312
rect 132770 1300 132776 1312
rect 132828 1300 132834 1352
rect 132954 1300 132960 1352
rect 133012 1340 133018 1352
rect 133966 1340 133972 1352
rect 133012 1312 133972 1340
rect 133012 1300 133018 1312
rect 133966 1300 133972 1312
rect 134024 1300 134030 1352
rect 137646 1300 137652 1352
rect 137704 1340 137710 1352
rect 138566 1340 138572 1352
rect 137704 1312 138572 1340
rect 137704 1300 137710 1312
rect 138566 1300 138572 1312
rect 138624 1300 138630 1352
rect 144730 1300 144736 1352
rect 144788 1340 144794 1352
rect 145558 1340 145564 1352
rect 144788 1312 145564 1340
rect 144788 1300 144794 1312
rect 145558 1300 145564 1312
rect 145616 1300 145622 1352
rect 145926 1300 145932 1352
rect 145984 1340 145990 1352
rect 146662 1340 146668 1352
rect 145984 1312 146668 1340
rect 145984 1300 145990 1312
rect 146662 1300 146668 1312
rect 146720 1300 146726 1352
rect 148318 1300 148324 1352
rect 148376 1340 148382 1352
rect 149054 1340 149060 1352
rect 148376 1312 149060 1340
rect 148376 1300 148382 1312
rect 149054 1300 149060 1312
rect 149112 1300 149118 1352
rect 154206 1300 154212 1352
rect 154264 1340 154270 1352
rect 154850 1340 154856 1352
rect 154264 1312 154856 1340
rect 154264 1300 154270 1312
rect 154850 1300 154856 1312
rect 154908 1300 154914 1352
rect 162486 1300 162492 1352
rect 162544 1340 162550 1352
rect 162946 1340 162952 1352
rect 162544 1312 162952 1340
rect 162544 1300 162550 1312
rect 162946 1300 162952 1312
rect 163004 1300 163010 1352
rect 266262 1300 266268 1352
rect 266320 1340 266326 1352
rect 267734 1340 267740 1352
rect 266320 1312 267740 1340
rect 266320 1300 266326 1312
rect 267734 1300 267740 1312
rect 267792 1300 267798 1352
rect 273162 1300 273168 1352
rect 273220 1340 273226 1352
rect 274818 1340 274824 1352
rect 273220 1312 274824 1340
rect 273220 1300 273226 1312
rect 274818 1300 274824 1312
rect 274876 1300 274882 1352
rect 280062 1300 280068 1352
rect 280120 1340 280126 1352
rect 281902 1340 281908 1352
rect 280120 1312 281908 1340
rect 280120 1300 280126 1312
rect 281902 1300 281908 1312
rect 281960 1300 281966 1352
rect 282546 1300 282552 1352
rect 282604 1340 282610 1352
rect 284294 1340 284300 1352
rect 282604 1312 284300 1340
rect 282604 1300 282610 1312
rect 284294 1300 284300 1312
rect 284352 1300 284358 1352
rect 288342 1300 288348 1352
rect 288400 1340 288406 1352
rect 290182 1340 290188 1352
rect 288400 1312 290188 1340
rect 288400 1300 288406 1312
rect 290182 1300 290188 1312
rect 290240 1300 290246 1352
rect 295242 1300 295248 1352
rect 295300 1340 295306 1352
rect 297266 1340 297272 1352
rect 295300 1312 297272 1340
rect 295300 1300 295306 1312
rect 297266 1300 297272 1312
rect 297324 1300 297330 1352
rect 297542 1300 297548 1352
rect 297600 1340 297606 1352
rect 299658 1340 299664 1352
rect 297600 1312 299664 1340
rect 297600 1300 297606 1312
rect 299658 1300 299664 1312
rect 299716 1300 299722 1352
rect 302142 1300 302148 1352
rect 302200 1340 302206 1352
rect 304350 1340 304356 1352
rect 302200 1312 304356 1340
rect 302200 1300 302206 1312
rect 304350 1300 304356 1312
rect 304408 1300 304414 1352
rect 305730 1300 305736 1352
rect 305788 1340 305794 1352
rect 307938 1340 307944 1352
rect 305788 1312 307944 1340
rect 305788 1300 305794 1312
rect 307938 1300 307944 1312
rect 307996 1300 308002 1352
rect 310330 1300 310336 1352
rect 310388 1340 310394 1352
rect 312630 1340 312636 1352
rect 310388 1312 312636 1340
rect 310388 1300 310394 1312
rect 312630 1300 312636 1312
rect 312688 1300 312694 1352
rect 313826 1300 313832 1352
rect 313884 1340 313890 1352
rect 316218 1340 316224 1352
rect 313884 1312 316224 1340
rect 313884 1300 313890 1312
rect 316218 1300 316224 1312
rect 316276 1300 316282 1352
rect 317230 1300 317236 1352
rect 317288 1340 317294 1352
rect 319714 1340 319720 1352
rect 317288 1312 319720 1340
rect 317288 1300 317294 1312
rect 319714 1300 319720 1312
rect 319772 1300 319778 1352
rect 321922 1300 321928 1352
rect 321980 1340 321986 1352
rect 324406 1340 324412 1352
rect 321980 1312 324412 1340
rect 321980 1300 321986 1312
rect 324406 1300 324412 1312
rect 324464 1300 324470 1352
rect 325418 1300 325424 1352
rect 325476 1340 325482 1352
rect 327994 1340 328000 1352
rect 325476 1312 328000 1340
rect 325476 1300 325482 1312
rect 327994 1300 328000 1312
rect 328052 1300 328058 1352
rect 328914 1300 328920 1352
rect 328972 1340 328978 1352
rect 331582 1340 331588 1352
rect 328972 1312 331588 1340
rect 328972 1300 328978 1312
rect 331582 1300 331588 1312
rect 331640 1300 331646 1352
rect 332410 1300 332416 1352
rect 332468 1340 332474 1352
rect 335078 1340 335084 1352
rect 332468 1312 335084 1340
rect 332468 1300 332474 1312
rect 335078 1300 335084 1312
rect 335136 1300 335142 1352
rect 335906 1300 335912 1352
rect 335964 1340 335970 1352
rect 338666 1340 338672 1352
rect 335964 1312 338672 1340
rect 335964 1300 335970 1312
rect 338666 1300 338672 1312
rect 338724 1300 338730 1352
rect 339310 1300 339316 1352
rect 339368 1340 339374 1352
rect 342162 1340 342168 1352
rect 339368 1312 342168 1340
rect 339368 1300 339374 1312
rect 342162 1300 342168 1312
rect 342220 1300 342226 1352
rect 345106 1300 345112 1352
rect 345164 1340 345170 1352
rect 348050 1340 348056 1352
rect 345164 1312 348056 1340
rect 345164 1300 345170 1312
rect 348050 1300 348056 1312
rect 348108 1300 348114 1352
rect 349798 1300 349804 1352
rect 349856 1340 349862 1352
rect 352834 1340 352840 1352
rect 349856 1312 352840 1340
rect 349856 1300 349862 1312
rect 352834 1300 352840 1312
rect 352892 1300 352898 1352
rect 353202 1300 353208 1352
rect 353260 1340 353266 1352
rect 356330 1340 356336 1352
rect 353260 1312 356336 1340
rect 353260 1300 353266 1312
rect 356330 1300 356336 1312
rect 356388 1300 356394 1352
rect 356698 1300 356704 1352
rect 356756 1340 356762 1352
rect 359918 1340 359924 1352
rect 356756 1312 359924 1340
rect 356756 1300 356762 1312
rect 359918 1300 359924 1312
rect 359976 1300 359982 1352
rect 362586 1300 362592 1352
rect 362644 1340 362650 1352
rect 365806 1340 365812 1352
rect 362644 1312 365812 1340
rect 362644 1300 362650 1312
rect 365806 1300 365812 1312
rect 365864 1300 365870 1352
rect 367186 1300 367192 1352
rect 367244 1340 367250 1352
rect 370590 1340 370596 1352
rect 367244 1312 370596 1340
rect 367244 1300 367250 1312
rect 370590 1300 370596 1312
rect 370648 1300 370654 1352
rect 370682 1300 370688 1352
rect 370740 1340 370746 1352
rect 374086 1340 374092 1352
rect 370740 1312 374092 1340
rect 370740 1300 370746 1312
rect 374086 1300 374092 1312
rect 374144 1300 374150 1352
rect 376386 1300 376392 1352
rect 376444 1340 376450 1352
rect 379974 1340 379980 1352
rect 376444 1312 379980 1340
rect 376444 1300 376450 1312
rect 379974 1300 379980 1312
rect 380032 1300 380038 1352
rect 385770 1300 385776 1352
rect 385828 1340 385834 1352
rect 389450 1340 389456 1352
rect 385828 1312 389456 1340
rect 385828 1300 385834 1312
rect 389450 1300 389456 1312
rect 389508 1300 389514 1352
rect 395062 1300 395068 1352
rect 395120 1340 395126 1352
rect 398926 1340 398932 1352
rect 395120 1312 398932 1340
rect 395120 1300 395126 1312
rect 398926 1300 398932 1312
rect 398984 1300 398990 1352
rect 399662 1300 399668 1352
rect 399720 1340 399726 1352
rect 403618 1340 403624 1352
rect 399720 1312 403624 1340
rect 399720 1300 399726 1312
rect 403618 1300 403624 1312
rect 403676 1300 403682 1352
rect 405458 1300 405464 1352
rect 405516 1340 405522 1352
rect 409598 1340 409604 1352
rect 405516 1312 409604 1340
rect 405516 1300 405522 1312
rect 409598 1300 409604 1312
rect 409656 1300 409662 1352
rect 415946 1300 415952 1352
rect 416004 1340 416010 1352
rect 420178 1340 420184 1352
rect 416004 1312 420184 1340
rect 416004 1300 416010 1312
rect 420178 1300 420184 1312
rect 420236 1300 420242 1352
rect 427538 1300 427544 1352
rect 427596 1340 427602 1352
rect 431862 1340 431868 1352
rect 427596 1312 431868 1340
rect 427596 1300 427602 1312
rect 431862 1300 431868 1312
rect 431920 1300 431926 1352
rect 433242 1300 433248 1352
rect 433300 1340 433306 1352
rect 437842 1340 437848 1352
rect 433300 1312 437848 1340
rect 433300 1300 433306 1312
rect 437842 1300 437848 1312
rect 437900 1300 437906 1352
rect 442626 1300 442632 1352
rect 442684 1340 442690 1352
rect 447410 1340 447416 1352
rect 442684 1312 447416 1340
rect 442684 1300 442690 1312
rect 447410 1300 447416 1312
rect 447468 1300 447474 1352
rect 448422 1300 448428 1352
rect 448480 1340 448486 1352
rect 453298 1340 453304 1352
rect 448480 1312 453304 1340
rect 448480 1300 448486 1312
rect 453298 1300 453304 1312
rect 453356 1300 453362 1352
rect 458818 1300 458824 1352
rect 458876 1340 458882 1352
rect 463970 1340 463976 1352
rect 458876 1312 463976 1340
rect 458876 1300 458882 1312
rect 463970 1300 463976 1312
rect 464028 1300 464034 1352
rect 468110 1300 468116 1352
rect 468168 1340 468174 1352
rect 473078 1340 473084 1352
rect 468168 1312 473084 1340
rect 468168 1300 468174 1312
rect 473078 1300 473084 1312
rect 473136 1300 473142 1352
rect 480898 1300 480904 1352
rect 480956 1340 480962 1352
rect 486418 1340 486424 1352
rect 480956 1312 486424 1340
rect 480956 1300 480962 1312
rect 486418 1300 486424 1312
rect 486476 1300 486482 1352
rect 487798 1300 487804 1352
rect 487856 1340 487862 1352
rect 493134 1340 493140 1352
rect 487856 1312 493140 1340
rect 487856 1300 487862 1312
rect 493134 1300 493140 1312
rect 493192 1300 493198 1352
rect 497090 1300 497096 1352
rect 497148 1340 497154 1352
rect 502978 1340 502984 1352
rect 497148 1312 502984 1340
rect 497148 1300 497154 1312
rect 502978 1300 502984 1312
rect 503036 1300 503042 1352
rect 504082 1300 504088 1352
rect 504140 1340 504146 1352
rect 509694 1340 509700 1352
rect 504140 1312 509700 1340
rect 504140 1300 504146 1312
rect 509694 1300 509700 1312
rect 509752 1300 509758 1352
rect 509878 1300 509884 1352
rect 509936 1340 509942 1352
rect 515766 1340 515772 1352
rect 509936 1312 515772 1340
rect 509936 1300 509942 1312
rect 515766 1300 515772 1312
rect 515824 1300 515830 1352
rect 519170 1300 519176 1352
rect 519228 1340 519234 1352
rect 525426 1340 525432 1352
rect 519228 1312 525432 1340
rect 519228 1300 519234 1312
rect 525426 1300 525432 1312
rect 525484 1300 525490 1352
rect 526070 1300 526076 1352
rect 526128 1340 526134 1352
rect 532142 1340 532148 1352
rect 526128 1312 532148 1340
rect 526128 1300 526134 1312
rect 532142 1300 532148 1312
rect 532200 1300 532206 1352
rect 534258 1300 534264 1352
rect 534316 1340 534322 1352
rect 540422 1340 540428 1352
rect 534316 1312 540428 1340
rect 534316 1300 534322 1312
rect 540422 1300 540428 1312
rect 540480 1300 540486 1352
rect 542262 1300 542268 1352
rect 542320 1340 542326 1352
rect 549070 1340 549076 1352
rect 542320 1312 549076 1340
rect 542320 1300 542326 1312
rect 549070 1300 549076 1312
rect 549128 1300 549134 1352
rect 551646 1300 551652 1352
rect 551704 1340 551710 1352
rect 558546 1340 558552 1352
rect 551704 1312 558552 1340
rect 551704 1300 551710 1312
rect 558546 1300 558552 1312
rect 558604 1300 558610 1352
rect 560938 1300 560944 1352
rect 560996 1340 561002 1352
rect 568022 1340 568028 1352
rect 560996 1312 568028 1340
rect 560996 1300 561002 1312
rect 568022 1300 568028 1312
rect 568080 1300 568086 1352
rect 571242 1300 571248 1352
rect 571300 1340 571306 1352
rect 578602 1340 578608 1352
rect 571300 1312 578608 1340
rect 571300 1300 571306 1312
rect 578602 1300 578608 1312
rect 578660 1300 578666 1352
rect 74994 1232 75000 1284
rect 75052 1272 75058 1284
rect 77110 1272 77116 1284
rect 75052 1244 77116 1272
rect 75052 1232 75058 1244
rect 77110 1232 77116 1244
rect 77168 1232 77174 1284
rect 77386 1232 77392 1284
rect 77444 1272 77450 1284
rect 79410 1272 79416 1284
rect 77444 1244 79416 1272
rect 77444 1232 77450 1244
rect 79410 1232 79416 1244
rect 79468 1232 79474 1284
rect 82078 1232 82084 1284
rect 82136 1272 82142 1284
rect 84010 1272 84016 1284
rect 82136 1244 84016 1272
rect 82136 1232 82142 1244
rect 84010 1232 84016 1244
rect 84068 1232 84074 1284
rect 84470 1232 84476 1284
rect 84528 1272 84534 1284
rect 86402 1272 86408 1284
rect 84528 1244 86408 1272
rect 84528 1232 84534 1244
rect 86402 1232 86408 1244
rect 86460 1232 86466 1284
rect 90358 1232 90364 1284
rect 90416 1272 90422 1284
rect 92198 1272 92204 1284
rect 90416 1244 92204 1272
rect 90416 1232 90422 1244
rect 92198 1232 92204 1244
rect 92256 1232 92262 1284
rect 92750 1232 92756 1284
rect 92808 1272 92814 1284
rect 94498 1272 94504 1284
rect 92808 1244 94504 1272
rect 92808 1232 92814 1244
rect 94498 1232 94504 1244
rect 94556 1232 94562 1284
rect 98638 1232 98644 1284
rect 98696 1272 98702 1284
rect 100294 1272 100300 1284
rect 98696 1244 100300 1272
rect 98696 1232 98702 1244
rect 100294 1232 100300 1244
rect 100352 1232 100358 1284
rect 102226 1232 102232 1284
rect 102284 1272 102290 1284
rect 103790 1272 103796 1284
rect 102284 1244 103796 1272
rect 102284 1232 102290 1244
rect 103790 1232 103796 1244
rect 103848 1232 103854 1284
rect 108114 1232 108120 1284
rect 108172 1272 108178 1284
rect 109586 1272 109592 1284
rect 108172 1244 109592 1272
rect 108172 1232 108178 1244
rect 109586 1232 109592 1244
rect 109644 1232 109650 1284
rect 110506 1232 110512 1284
rect 110564 1272 110570 1284
rect 111886 1272 111892 1284
rect 110564 1244 111892 1272
rect 110564 1232 110570 1244
rect 111886 1232 111892 1244
rect 111944 1232 111950 1284
rect 115198 1232 115204 1284
rect 115256 1272 115262 1284
rect 116578 1272 116584 1284
rect 115256 1244 116584 1272
rect 115256 1232 115262 1244
rect 116578 1232 116584 1244
rect 116636 1232 116642 1284
rect 117590 1232 117596 1284
rect 117648 1272 117654 1284
rect 118878 1272 118884 1284
rect 117648 1244 118884 1272
rect 117648 1232 117654 1244
rect 118878 1232 118884 1244
rect 118936 1232 118942 1284
rect 122282 1232 122288 1284
rect 122340 1272 122346 1284
rect 123478 1272 123484 1284
rect 122340 1244 123484 1272
rect 122340 1232 122346 1244
rect 123478 1232 123484 1244
rect 123536 1232 123542 1284
rect 124674 1232 124680 1284
rect 124732 1272 124738 1284
rect 125778 1272 125784 1284
rect 124732 1244 125784 1272
rect 124732 1232 124738 1244
rect 125778 1232 125784 1244
rect 125836 1232 125842 1284
rect 128170 1232 128176 1284
rect 128228 1272 128234 1284
rect 129274 1272 129280 1284
rect 128228 1244 129280 1272
rect 128228 1232 128234 1244
rect 129274 1232 129280 1244
rect 129332 1232 129338 1284
rect 136450 1232 136456 1284
rect 136508 1272 136514 1284
rect 137370 1272 137376 1284
rect 136508 1244 137376 1272
rect 136508 1232 136514 1244
rect 137370 1232 137376 1244
rect 137428 1232 137434 1284
rect 138842 1232 138848 1284
rect 138900 1272 138906 1284
rect 139762 1272 139768 1284
rect 138900 1244 139768 1272
rect 138900 1232 138906 1244
rect 139762 1232 139768 1244
rect 139820 1232 139826 1284
rect 140038 1232 140044 1284
rect 140096 1272 140102 1284
rect 140866 1272 140872 1284
rect 140096 1244 140872 1272
rect 140096 1232 140102 1244
rect 140866 1232 140872 1244
rect 140924 1232 140930 1284
rect 281350 1232 281356 1284
rect 281408 1272 281414 1284
rect 283098 1272 283104 1284
rect 281408 1244 283104 1272
rect 281408 1232 281414 1244
rect 283098 1232 283104 1244
rect 283156 1232 283162 1284
rect 289446 1232 289452 1284
rect 289504 1272 289510 1284
rect 291378 1272 291384 1284
rect 289504 1244 291384 1272
rect 289504 1232 289510 1244
rect 291378 1232 291384 1244
rect 291436 1232 291442 1284
rect 296438 1232 296444 1284
rect 296496 1272 296502 1284
rect 298462 1272 298468 1284
rect 296496 1244 298468 1272
rect 296496 1232 296502 1244
rect 298462 1232 298468 1244
rect 298520 1232 298526 1284
rect 303338 1232 303344 1284
rect 303396 1272 303402 1284
rect 305546 1272 305552 1284
rect 303396 1244 305552 1272
rect 303396 1232 303402 1244
rect 305546 1232 305552 1244
rect 305604 1232 305610 1284
rect 312538 1232 312544 1284
rect 312596 1272 312602 1284
rect 315022 1272 315028 1284
rect 312596 1244 315028 1272
rect 312596 1232 312602 1244
rect 315022 1232 315028 1244
rect 315080 1232 315086 1284
rect 318426 1232 318432 1284
rect 318484 1272 318490 1284
rect 320910 1272 320916 1284
rect 318484 1244 320916 1272
rect 318484 1232 318490 1244
rect 320910 1232 320916 1244
rect 320968 1232 320974 1284
rect 324222 1232 324228 1284
rect 324280 1272 324286 1284
rect 326798 1272 326804 1284
rect 324280 1244 326804 1272
rect 324280 1232 324286 1244
rect 326798 1232 326804 1244
rect 326856 1232 326862 1284
rect 330018 1232 330024 1284
rect 330076 1272 330082 1284
rect 332686 1272 332692 1284
rect 330076 1244 332692 1272
rect 330076 1232 330082 1244
rect 332686 1232 332692 1244
rect 332744 1232 332750 1284
rect 334710 1232 334716 1284
rect 334768 1272 334774 1284
rect 337470 1272 337476 1284
rect 334768 1244 337476 1272
rect 334768 1232 334774 1244
rect 337470 1232 337476 1244
rect 337528 1232 337534 1284
rect 340506 1232 340512 1284
rect 340564 1272 340570 1284
rect 343358 1272 343364 1284
rect 340564 1244 343364 1272
rect 340564 1232 340570 1244
rect 343358 1232 343364 1244
rect 343416 1232 343422 1284
rect 344002 1232 344008 1284
rect 344060 1272 344066 1284
rect 346946 1272 346952 1284
rect 344060 1244 346952 1272
rect 344060 1232 344066 1244
rect 346946 1232 346952 1244
rect 347004 1232 347010 1284
rect 348602 1232 348608 1284
rect 348660 1272 348666 1284
rect 351638 1272 351644 1284
rect 348660 1244 351644 1272
rect 348660 1232 348666 1244
rect 351638 1232 351644 1244
rect 351696 1232 351702 1284
rect 352098 1232 352104 1284
rect 352156 1272 352162 1284
rect 355226 1272 355232 1284
rect 352156 1244 355232 1272
rect 352156 1232 352162 1244
rect 355226 1232 355232 1244
rect 355284 1232 355290 1284
rect 355594 1232 355600 1284
rect 355652 1272 355658 1284
rect 358722 1272 358728 1284
rect 355652 1244 358728 1272
rect 355652 1232 355658 1244
rect 358722 1232 358728 1244
rect 358780 1232 358786 1284
rect 359090 1232 359096 1284
rect 359148 1272 359154 1284
rect 362310 1272 362316 1284
rect 359148 1244 362316 1272
rect 359148 1232 359154 1244
rect 362310 1232 362316 1244
rect 362368 1232 362374 1284
rect 363690 1232 363696 1284
rect 363748 1272 363754 1284
rect 367002 1272 367008 1284
rect 363748 1244 367008 1272
rect 363748 1232 363754 1244
rect 367002 1232 367008 1244
rect 367060 1232 367066 1284
rect 372982 1232 372988 1284
rect 373040 1272 373046 1284
rect 376478 1272 376484 1284
rect 373040 1244 376484 1272
rect 373040 1232 373046 1244
rect 376478 1232 376484 1244
rect 376536 1232 376542 1284
rect 377582 1232 377588 1284
rect 377640 1272 377646 1284
rect 381170 1272 381176 1284
rect 377640 1244 381176 1272
rect 377640 1232 377646 1244
rect 381170 1232 381176 1244
rect 381228 1232 381234 1284
rect 388070 1232 388076 1284
rect 388128 1272 388134 1284
rect 391842 1272 391848 1284
rect 388128 1244 391848 1272
rect 388128 1232 388134 1244
rect 391842 1232 391848 1244
rect 391900 1232 391906 1284
rect 393866 1232 393872 1284
rect 393924 1272 393930 1284
rect 397730 1272 397736 1284
rect 393924 1244 397736 1272
rect 393924 1232 393930 1244
rect 397730 1232 397736 1244
rect 397788 1232 397794 1284
rect 398466 1232 398472 1284
rect 398524 1272 398530 1284
rect 402514 1272 402520 1284
rect 398524 1244 402520 1272
rect 398524 1232 398530 1244
rect 402514 1232 402520 1244
rect 402572 1232 402578 1284
rect 403158 1232 403164 1284
rect 403216 1272 403222 1284
rect 407206 1272 407212 1284
rect 403216 1244 407212 1272
rect 403216 1232 403222 1244
rect 407206 1232 407212 1244
rect 407264 1232 407270 1284
rect 410058 1232 410064 1284
rect 410116 1272 410122 1284
rect 414290 1272 414296 1284
rect 410116 1244 414296 1272
rect 410116 1232 410122 1244
rect 414290 1232 414296 1244
rect 414348 1232 414354 1284
rect 418246 1232 418252 1284
rect 418304 1272 418310 1284
rect 422570 1272 422576 1284
rect 418304 1244 422576 1272
rect 418304 1232 418310 1244
rect 422570 1232 422576 1244
rect 422628 1232 422634 1284
rect 424042 1232 424048 1284
rect 424100 1272 424106 1284
rect 428458 1272 428464 1284
rect 424100 1244 428464 1272
rect 424100 1232 424106 1244
rect 428458 1232 428464 1244
rect 428516 1232 428522 1284
rect 435634 1232 435640 1284
rect 435692 1272 435698 1284
rect 439958 1272 439964 1284
rect 435692 1244 439964 1272
rect 435692 1232 435698 1244
rect 439958 1232 439964 1244
rect 440016 1232 440022 1284
rect 444926 1232 444932 1284
rect 444984 1272 444990 1284
rect 449802 1272 449808 1284
rect 444984 1244 449808 1272
rect 444984 1232 444990 1244
rect 449802 1232 449808 1244
rect 449860 1232 449866 1284
rect 450722 1232 450728 1284
rect 450780 1272 450786 1284
rect 455690 1272 455696 1284
rect 450780 1244 455696 1272
rect 450780 1232 450786 1244
rect 455690 1232 455696 1244
rect 455748 1232 455754 1284
rect 456518 1232 456524 1284
rect 456576 1272 456582 1284
rect 461578 1272 461584 1284
rect 456576 1244 461584 1272
rect 456576 1232 456582 1244
rect 461578 1232 461584 1244
rect 461636 1232 461642 1284
rect 462222 1232 462228 1284
rect 462280 1272 462286 1284
rect 467466 1272 467472 1284
rect 462280 1244 467472 1272
rect 462280 1232 462286 1244
rect 467466 1232 467472 1244
rect 467524 1232 467530 1284
rect 471606 1232 471612 1284
rect 471664 1272 471670 1284
rect 476574 1272 476580 1284
rect 471664 1244 476580 1272
rect 471664 1232 471670 1244
rect 476574 1232 476580 1244
rect 476632 1232 476638 1284
rect 479702 1232 479708 1284
rect 479760 1272 479766 1284
rect 484854 1272 484860 1284
rect 479760 1244 484860 1272
rect 479760 1232 479766 1244
rect 484854 1232 484860 1244
rect 484912 1232 484918 1284
rect 488994 1232 489000 1284
rect 489052 1272 489058 1284
rect 494698 1272 494704 1284
rect 489052 1244 494704 1272
rect 489052 1232 489058 1244
rect 494698 1232 494704 1244
rect 494756 1232 494762 1284
rect 498286 1232 498292 1284
rect 498344 1272 498350 1284
rect 503806 1272 503812 1284
rect 498344 1244 503812 1272
rect 498344 1232 498350 1244
rect 503806 1232 503812 1244
rect 503864 1232 503870 1284
rect 510982 1232 510988 1284
rect 511040 1272 511046 1284
rect 517146 1272 517152 1284
rect 511040 1244 517152 1272
rect 511040 1232 511046 1244
rect 517146 1232 517152 1244
rect 517204 1232 517210 1284
rect 517974 1232 517980 1284
rect 518032 1272 518038 1284
rect 523862 1272 523868 1284
rect 518032 1244 523868 1272
rect 518032 1232 518038 1244
rect 523862 1232 523868 1244
rect 523920 1232 523926 1284
rect 527266 1232 527272 1284
rect 527324 1272 527330 1284
rect 533706 1272 533712 1284
rect 527324 1244 533712 1272
rect 527324 1232 527330 1244
rect 533706 1232 533712 1244
rect 533764 1232 533770 1284
rect 543458 1232 543464 1284
rect 543516 1272 543522 1284
rect 550266 1272 550272 1284
rect 543516 1244 550272 1272
rect 543516 1232 543522 1244
rect 550266 1232 550272 1244
rect 550324 1232 550330 1284
rect 550450 1232 550456 1284
rect 550508 1272 550514 1284
rect 557350 1272 557356 1284
rect 550508 1244 557356 1272
rect 550508 1232 550514 1244
rect 557350 1232 557356 1244
rect 557408 1232 557414 1284
rect 562042 1232 562048 1284
rect 562100 1272 562106 1284
rect 569126 1272 569132 1284
rect 562100 1244 569132 1272
rect 562100 1232 562106 1244
rect 569126 1232 569132 1244
rect 569184 1232 569190 1284
rect 570138 1232 570144 1284
rect 570196 1272 570202 1284
rect 577406 1272 577412 1284
rect 570196 1244 577412 1272
rect 570196 1232 570202 1244
rect 577406 1232 577412 1244
rect 577464 1232 577470 1284
rect 99834 1164 99840 1216
rect 99892 1204 99898 1216
rect 101490 1204 101496 1216
rect 99892 1176 101496 1204
rect 99892 1164 99898 1176
rect 101490 1164 101496 1176
rect 101548 1164 101554 1216
rect 114002 1164 114008 1216
rect 114060 1204 114066 1216
rect 115382 1204 115388 1216
rect 114060 1176 115388 1204
rect 114060 1164 114066 1176
rect 115382 1164 115388 1176
rect 115440 1164 115446 1216
rect 311526 1164 311532 1216
rect 311584 1204 311590 1216
rect 313826 1204 313832 1216
rect 311584 1176 313832 1204
rect 311584 1164 311590 1176
rect 313826 1164 313832 1176
rect 313884 1164 313890 1216
rect 319622 1164 319628 1216
rect 319680 1204 319686 1216
rect 322106 1204 322112 1216
rect 319680 1176 322112 1204
rect 319680 1164 319686 1176
rect 322106 1164 322112 1176
rect 322164 1164 322170 1216
rect 326614 1164 326620 1216
rect 326672 1204 326678 1216
rect 329190 1204 329196 1216
rect 326672 1176 329196 1204
rect 326672 1164 326678 1176
rect 329190 1164 329196 1176
rect 329248 1164 329254 1216
rect 331122 1164 331128 1216
rect 331180 1204 331186 1216
rect 333882 1204 333888 1216
rect 331180 1176 333888 1204
rect 331180 1164 331186 1176
rect 333882 1164 333888 1176
rect 333940 1164 333946 1216
rect 337010 1164 337016 1216
rect 337068 1204 337074 1216
rect 339862 1204 339868 1216
rect 337068 1176 339868 1204
rect 337068 1164 337074 1176
rect 339862 1164 339868 1176
rect 339920 1164 339926 1216
rect 341702 1164 341708 1216
rect 341760 1204 341766 1216
rect 344554 1204 344560 1216
rect 341760 1176 344560 1204
rect 341760 1164 341766 1176
rect 344554 1164 344560 1176
rect 344612 1164 344618 1216
rect 357894 1164 357900 1216
rect 357952 1204 357958 1216
rect 361114 1204 361120 1216
rect 357952 1176 361120 1204
rect 357952 1164 357958 1176
rect 361114 1164 361120 1176
rect 361172 1164 361178 1216
rect 364886 1164 364892 1216
rect 364944 1204 364950 1216
rect 368198 1204 368204 1216
rect 364944 1176 368204 1204
rect 364944 1164 364950 1176
rect 368198 1164 368204 1176
rect 368256 1164 368262 1216
rect 375282 1164 375288 1216
rect 375340 1204 375346 1216
rect 378870 1204 378876 1216
rect 375340 1176 378876 1204
rect 375340 1164 375346 1176
rect 378870 1164 378876 1176
rect 378928 1164 378934 1216
rect 381078 1164 381084 1216
rect 381136 1204 381142 1216
rect 384758 1204 384764 1216
rect 381136 1176 384764 1204
rect 381136 1164 381142 1176
rect 384758 1164 384764 1176
rect 384816 1164 384822 1216
rect 390370 1164 390376 1216
rect 390428 1204 390434 1216
rect 394234 1204 394240 1216
rect 390428 1176 394240 1204
rect 390428 1164 390434 1176
rect 394234 1164 394240 1176
rect 394292 1164 394298 1216
rect 400858 1164 400864 1216
rect 400916 1204 400922 1216
rect 404814 1204 404820 1216
rect 400916 1176 404820 1204
rect 400916 1164 400922 1176
rect 404814 1164 404820 1176
rect 404872 1164 404878 1216
rect 407758 1164 407764 1216
rect 407816 1204 407822 1216
rect 411898 1204 411904 1216
rect 407816 1176 411904 1204
rect 407816 1164 407822 1176
rect 411898 1164 411904 1176
rect 411956 1164 411962 1216
rect 413554 1164 413560 1216
rect 413612 1204 413618 1216
rect 417878 1204 417884 1216
rect 413612 1176 417884 1204
rect 413612 1164 413618 1176
rect 417878 1164 417884 1176
rect 417936 1164 417942 1216
rect 419350 1164 419356 1216
rect 419408 1204 419414 1216
rect 423398 1204 423404 1216
rect 419408 1176 423404 1204
rect 419408 1164 419414 1176
rect 423398 1164 423404 1176
rect 423456 1164 423462 1216
rect 426342 1164 426348 1216
rect 426400 1204 426406 1216
rect 430850 1204 430856 1216
rect 426400 1176 430856 1204
rect 426400 1164 426406 1176
rect 430850 1164 430856 1176
rect 430908 1164 430914 1216
rect 441430 1164 441436 1216
rect 441488 1204 441494 1216
rect 445846 1204 445852 1216
rect 441488 1176 445852 1204
rect 441488 1164 441494 1176
rect 445846 1164 445852 1176
rect 445904 1164 445910 1216
rect 446030 1164 446036 1216
rect 446088 1204 446094 1216
rect 450906 1204 450912 1216
rect 446088 1176 450912 1204
rect 446088 1164 446094 1176
rect 450906 1164 450912 1176
rect 450964 1164 450970 1216
rect 457622 1164 457628 1216
rect 457680 1204 457686 1216
rect 462406 1204 462412 1216
rect 457680 1176 462412 1204
rect 457680 1164 457686 1176
rect 462406 1164 462412 1176
rect 462464 1164 462470 1216
rect 465810 1164 465816 1216
rect 465868 1204 465874 1216
rect 470686 1204 470692 1216
rect 465868 1176 470692 1204
rect 465868 1164 465874 1176
rect 470686 1164 470692 1176
rect 470744 1164 470750 1216
rect 475102 1164 475108 1216
rect 475160 1204 475166 1216
rect 480530 1204 480536 1216
rect 475160 1176 480536 1204
rect 475160 1164 475166 1176
rect 480530 1164 480536 1176
rect 480588 1164 480594 1216
rect 482002 1164 482008 1216
rect 482060 1204 482066 1216
rect 487246 1204 487252 1216
rect 482060 1176 487252 1204
rect 482060 1164 482066 1176
rect 487246 1164 487252 1176
rect 487304 1164 487310 1216
rect 492490 1164 492496 1216
rect 492548 1204 492554 1216
rect 498194 1204 498200 1216
rect 492548 1176 498200 1204
rect 492548 1164 492554 1176
rect 498194 1164 498200 1176
rect 498252 1164 498258 1216
rect 505186 1164 505192 1216
rect 505244 1204 505250 1216
rect 511258 1204 511264 1216
rect 505244 1176 511264 1204
rect 505244 1164 505250 1176
rect 511258 1164 511264 1176
rect 511316 1164 511322 1216
rect 513282 1164 513288 1216
rect 513340 1204 513346 1216
rect 519538 1204 519544 1216
rect 513340 1176 519544 1204
rect 513340 1164 513346 1176
rect 519538 1164 519544 1176
rect 519596 1164 519602 1216
rect 522666 1164 522672 1216
rect 522724 1204 522730 1216
rect 529014 1204 529020 1216
rect 522724 1176 529020 1204
rect 522724 1164 522730 1176
rect 529014 1164 529020 1176
rect 529072 1164 529078 1216
rect 531866 1164 531872 1216
rect 531924 1204 531930 1216
rect 538398 1204 538404 1216
rect 531924 1176 538404 1204
rect 531924 1164 531930 1176
rect 538398 1164 538404 1176
rect 538456 1164 538462 1216
rect 540054 1164 540060 1216
rect 540112 1204 540118 1216
rect 546678 1204 546684 1216
rect 540112 1176 546684 1204
rect 540112 1164 540118 1176
rect 546678 1164 546684 1176
rect 546736 1164 546742 1216
rect 548150 1164 548156 1216
rect 548208 1204 548214 1216
rect 554958 1204 554964 1216
rect 548208 1176 554964 1204
rect 548208 1164 548214 1176
rect 554958 1164 554964 1176
rect 555016 1164 555022 1216
rect 558454 1164 558460 1216
rect 558512 1204 558518 1216
rect 565630 1204 565636 1216
rect 558512 1176 565636 1204
rect 558512 1164 558518 1176
rect 565630 1164 565636 1176
rect 565688 1164 565694 1216
rect 569034 1164 569040 1216
rect 569092 1204 569098 1216
rect 576302 1204 576308 1216
rect 569092 1176 576308 1204
rect 569092 1164 569098 1176
rect 576302 1164 576308 1176
rect 576360 1164 576366 1216
rect 5626 1096 5632 1148
rect 5684 1136 5690 1148
rect 8662 1136 8668 1148
rect 5684 1108 8668 1136
rect 5684 1096 5690 1108
rect 8662 1096 8668 1108
rect 8720 1096 8726 1148
rect 111610 1096 111616 1148
rect 111668 1136 111674 1148
rect 113082 1136 113088 1148
rect 111668 1108 113088 1136
rect 111668 1096 111674 1108
rect 113082 1096 113088 1108
rect 113140 1096 113146 1148
rect 123478 1096 123484 1148
rect 123536 1136 123542 1148
rect 124766 1136 124772 1148
rect 123536 1108 124772 1136
rect 123536 1096 123542 1108
rect 124766 1096 124772 1108
rect 124824 1096 124830 1148
rect 320818 1096 320824 1148
rect 320876 1136 320882 1148
rect 323302 1136 323308 1148
rect 320876 1108 323308 1136
rect 320876 1096 320882 1108
rect 323302 1096 323308 1108
rect 323360 1096 323366 1148
rect 327718 1096 327724 1148
rect 327776 1136 327782 1148
rect 330386 1136 330392 1148
rect 327776 1108 330392 1136
rect 327776 1096 327782 1108
rect 330386 1096 330392 1108
rect 330444 1096 330450 1148
rect 360102 1096 360108 1148
rect 360160 1136 360166 1148
rect 363506 1136 363512 1148
rect 360160 1108 363512 1136
rect 360160 1096 360166 1108
rect 363506 1096 363512 1108
rect 363564 1096 363570 1148
rect 382182 1096 382188 1148
rect 382240 1136 382246 1148
rect 385954 1136 385960 1148
rect 382240 1108 385960 1136
rect 382240 1096 382246 1108
rect 385954 1096 385960 1108
rect 386012 1096 386018 1148
rect 389266 1096 389272 1148
rect 389324 1136 389330 1148
rect 393038 1136 393044 1148
rect 389324 1108 393044 1136
rect 389324 1096 389330 1108
rect 393038 1096 393044 1108
rect 393096 1096 393102 1148
rect 397362 1096 397368 1148
rect 397420 1136 397426 1148
rect 401318 1136 401324 1148
rect 397420 1108 401324 1136
rect 397420 1096 397426 1108
rect 401318 1096 401324 1108
rect 401376 1096 401382 1148
rect 404262 1096 404268 1148
rect 404320 1136 404326 1148
rect 408402 1136 408408 1148
rect 404320 1108 408408 1136
rect 404320 1096 404326 1108
rect 408402 1096 408408 1108
rect 408460 1096 408466 1148
rect 408954 1096 408960 1148
rect 409012 1136 409018 1148
rect 413094 1136 413100 1148
rect 409012 1108 413100 1136
rect 409012 1096 409018 1108
rect 413094 1096 413100 1108
rect 413152 1096 413158 1148
rect 420546 1096 420552 1148
rect 420604 1136 420610 1148
rect 424962 1136 424968 1148
rect 420604 1108 424968 1136
rect 420604 1096 420610 1108
rect 424962 1096 424968 1108
rect 425020 1096 425026 1148
rect 428642 1096 428648 1148
rect 428700 1136 428706 1148
rect 433242 1136 433248 1148
rect 428700 1108 433248 1136
rect 428700 1096 428706 1108
rect 433242 1096 433248 1108
rect 433300 1096 433306 1148
rect 436738 1096 436744 1148
rect 436796 1136 436802 1148
rect 441522 1136 441528 1148
rect 436796 1108 441528 1136
rect 436796 1096 436802 1108
rect 441522 1096 441528 1108
rect 441580 1096 441586 1148
rect 454218 1096 454224 1148
rect 454276 1136 454282 1148
rect 459186 1136 459192 1148
rect 454276 1108 459192 1136
rect 454276 1096 454282 1108
rect 459186 1096 459192 1108
rect 459244 1096 459250 1148
rect 461118 1096 461124 1148
rect 461176 1136 461182 1148
rect 466270 1136 466276 1148
rect 461176 1108 466276 1136
rect 461176 1096 461182 1108
rect 466270 1096 466276 1108
rect 466328 1096 466334 1148
rect 472710 1096 472716 1148
rect 472768 1136 472774 1148
rect 478138 1136 478144 1148
rect 472768 1108 478144 1136
rect 472768 1096 472774 1108
rect 478138 1096 478144 1108
rect 478196 1096 478202 1148
rect 486694 1096 486700 1148
rect 486752 1136 486758 1148
rect 492306 1136 492312 1148
rect 486752 1108 492312 1136
rect 486752 1096 486758 1108
rect 492306 1096 492312 1108
rect 492364 1096 492370 1148
rect 493594 1096 493600 1148
rect 493652 1136 493658 1148
rect 499390 1136 499396 1148
rect 493652 1108 499396 1136
rect 493652 1096 493658 1108
rect 499390 1096 499396 1108
rect 499448 1096 499454 1148
rect 500494 1096 500500 1148
rect 500552 1136 500558 1148
rect 506474 1136 506480 1148
rect 500552 1108 506480 1136
rect 500552 1096 500558 1108
rect 506474 1096 506480 1108
rect 506532 1096 506538 1148
rect 512178 1096 512184 1148
rect 512236 1136 512242 1148
rect 517974 1136 517980 1148
rect 512236 1108 517980 1136
rect 512236 1096 512242 1108
rect 517974 1096 517980 1108
rect 518032 1096 518038 1148
rect 523770 1096 523776 1148
rect 523828 1136 523834 1148
rect 530118 1136 530124 1148
rect 523828 1108 530124 1136
rect 523828 1096 523834 1108
rect 530118 1096 530124 1108
rect 530176 1096 530182 1148
rect 530762 1096 530768 1148
rect 530820 1136 530826 1148
rect 537202 1136 537208 1148
rect 530820 1108 537208 1136
rect 530820 1096 530826 1108
rect 537202 1096 537208 1108
rect 537260 1096 537266 1148
rect 538858 1096 538864 1148
rect 538916 1136 538922 1148
rect 545482 1136 545488 1148
rect 538916 1108 545488 1136
rect 538916 1096 538922 1108
rect 545482 1096 545488 1108
rect 545540 1096 545546 1148
rect 552750 1096 552756 1148
rect 552808 1136 552814 1148
rect 559742 1136 559748 1148
rect 552808 1108 559748 1136
rect 552808 1096 552814 1108
rect 559742 1096 559748 1108
rect 559800 1096 559806 1148
rect 567838 1096 567844 1148
rect 567896 1136 567902 1148
rect 575106 1136 575112 1148
rect 567896 1108 575112 1136
rect 567896 1096 567902 1108
rect 575106 1096 575112 1108
rect 575164 1096 575170 1148
rect 378778 1028 378784 1080
rect 378836 1068 378842 1080
rect 382366 1068 382372 1080
rect 378836 1040 382372 1068
rect 378836 1028 378842 1040
rect 382366 1028 382372 1040
rect 382424 1028 382430 1080
rect 386874 1028 386880 1080
rect 386932 1068 386938 1080
rect 390646 1068 390652 1080
rect 386932 1040 390652 1068
rect 386932 1028 386938 1040
rect 390646 1028 390652 1040
rect 390704 1028 390710 1080
rect 425146 1028 425152 1080
rect 425204 1068 425210 1080
rect 429654 1068 429660 1080
rect 425204 1040 429660 1068
rect 425204 1028 425210 1040
rect 429654 1028 429660 1040
rect 429712 1028 429718 1080
rect 439130 1028 439136 1080
rect 439188 1068 439194 1080
rect 443822 1068 443828 1080
rect 439188 1040 443828 1068
rect 439188 1028 439194 1040
rect 443822 1028 443828 1040
rect 443880 1028 443886 1080
rect 447226 1028 447232 1080
rect 447284 1068 447290 1080
rect 452102 1068 452108 1080
rect 447284 1040 452108 1068
rect 447284 1028 447290 1040
rect 452102 1028 452108 1040
rect 452160 1028 452166 1080
rect 455322 1028 455328 1080
rect 455380 1068 455386 1080
rect 460106 1068 460112 1080
rect 455380 1040 460112 1068
rect 455380 1028 455386 1040
rect 460106 1028 460112 1040
rect 460164 1028 460170 1080
rect 466914 1028 466920 1080
rect 466972 1068 466978 1080
rect 472250 1068 472256 1080
rect 466972 1040 472256 1068
rect 466972 1028 466978 1040
rect 472250 1028 472256 1040
rect 472308 1028 472314 1080
rect 477402 1028 477408 1080
rect 477460 1068 477466 1080
rect 482462 1068 482468 1080
rect 477460 1040 482468 1068
rect 477460 1028 477466 1040
rect 482462 1028 482468 1040
rect 482520 1028 482526 1080
rect 485498 1028 485504 1080
rect 485556 1068 485562 1080
rect 490742 1068 490748 1080
rect 485556 1040 490748 1068
rect 485556 1028 485562 1040
rect 490742 1028 490748 1040
rect 490800 1028 490806 1080
rect 494790 1028 494796 1080
rect 494848 1068 494854 1080
rect 500586 1068 500592 1080
rect 494848 1040 500592 1068
rect 494848 1028 494854 1040
rect 500586 1028 500592 1040
rect 500644 1028 500650 1080
rect 501690 1028 501696 1080
rect 501748 1068 501754 1080
rect 507302 1068 507308 1080
rect 501748 1040 507308 1068
rect 501748 1028 501754 1040
rect 507302 1028 507308 1040
rect 507360 1028 507366 1080
rect 514478 1028 514484 1080
rect 514536 1068 514542 1080
rect 520734 1068 520740 1080
rect 514536 1040 520740 1068
rect 514536 1028 514542 1040
rect 520734 1028 520740 1040
rect 520792 1028 520798 1080
rect 521470 1028 521476 1080
rect 521528 1068 521534 1080
rect 527818 1068 527824 1080
rect 521528 1040 527824 1068
rect 521528 1028 521534 1040
rect 527818 1028 527824 1040
rect 527876 1028 527882 1080
rect 529566 1028 529572 1080
rect 529624 1068 529630 1080
rect 536098 1068 536104 1080
rect 529624 1040 536104 1068
rect 529624 1028 529630 1040
rect 536098 1028 536104 1040
rect 536156 1028 536162 1080
rect 549346 1028 549352 1080
rect 549404 1068 549410 1080
rect 556154 1068 556160 1080
rect 549404 1040 556160 1068
rect 549404 1028 549410 1040
rect 556154 1028 556160 1040
rect 556212 1028 556218 1080
rect 559650 1028 559656 1080
rect 559708 1068 559714 1080
rect 566826 1068 566832 1080
rect 559708 1040 566832 1068
rect 559708 1028 559714 1040
rect 566826 1028 566832 1040
rect 566884 1028 566890 1080
rect 374178 960 374184 1012
rect 374236 1000 374242 1012
rect 377674 1000 377680 1012
rect 374236 972 377680 1000
rect 374236 960 374242 972
rect 377674 960 377680 972
rect 377732 960 377738 1012
rect 379882 960 379888 1012
rect 379940 1000 379946 1012
rect 383562 1000 383568 1012
rect 379940 972 383568 1000
rect 379940 960 379946 972
rect 383562 960 383568 972
rect 383620 960 383626 1012
rect 414750 960 414756 1012
rect 414808 1000 414814 1012
rect 418982 1000 418988 1012
rect 414808 972 418988 1000
rect 414808 960 414814 972
rect 418982 960 418988 972
rect 419040 960 419046 1012
rect 422846 960 422852 1012
rect 422904 1000 422910 1012
rect 427262 1000 427268 1012
rect 422904 972 427268 1000
rect 422904 960 422910 972
rect 427262 960 427268 972
rect 427320 960 427326 1012
rect 432138 960 432144 1012
rect 432196 1000 432202 1012
rect 436738 1000 436744 1012
rect 432196 972 436744 1000
rect 432196 960 432202 972
rect 436738 960 436744 972
rect 436796 960 436802 1012
rect 453022 960 453028 1012
rect 453080 1000 453086 1012
rect 458082 1000 458088 1012
rect 453080 972 458088 1000
rect 453080 960 453086 972
rect 458082 960 458088 972
rect 458140 960 458146 1012
rect 464614 960 464620 1012
rect 464672 1000 464678 1012
rect 469858 1000 469864 1012
rect 464672 972 469864 1000
rect 464672 960 464678 972
rect 469858 960 469864 972
rect 469916 960 469922 1012
rect 473906 960 473912 1012
rect 473964 1000 473970 1012
rect 479334 1000 479340 1012
rect 473964 972 479340 1000
rect 473964 960 473970 972
rect 479334 960 479340 972
rect 479392 960 479398 1012
rect 484302 960 484308 1012
rect 484360 1000 484366 1012
rect 489914 1000 489920 1012
rect 484360 972 489920 1000
rect 484360 960 484366 972
rect 489914 960 489920 972
rect 489972 960 489978 1012
rect 490098 960 490104 1012
rect 490156 1000 490162 1012
rect 495526 1000 495532 1012
rect 490156 972 495532 1000
rect 490156 960 490162 972
rect 495526 960 495532 972
rect 495584 960 495590 1012
rect 495986 960 495992 1012
rect 496044 1000 496050 1012
rect 501782 1000 501788 1012
rect 496044 972 501788 1000
rect 496044 960 496050 972
rect 501782 960 501788 972
rect 501840 960 501846 1012
rect 502886 960 502892 1012
rect 502944 1000 502950 1012
rect 508866 1000 508872 1012
rect 502944 972 508872 1000
rect 502944 960 502950 972
rect 508866 960 508872 972
rect 508924 960 508930 1012
rect 520182 960 520188 1012
rect 520240 1000 520246 1012
rect 526622 1000 526628 1012
rect 520240 972 526628 1000
rect 520240 960 520246 972
rect 526622 960 526628 972
rect 526680 960 526686 1012
rect 533062 960 533068 1012
rect 533120 1000 533126 1012
rect 539594 1000 539600 1012
rect 533120 972 539600 1000
rect 533120 960 533126 972
rect 539594 960 539600 972
rect 539652 960 539658 1012
rect 8754 892 8760 944
rect 8812 932 8818 944
rect 12158 932 12164 944
rect 8812 904 12164 932
rect 8812 892 8818 904
rect 12158 892 12164 904
rect 12216 892 12222 944
rect 121086 892 121092 944
rect 121144 932 121150 944
rect 122374 932 122380 944
rect 121144 904 122380 932
rect 121144 892 121150 904
rect 122374 892 122380 904
rect 122432 892 122438 944
rect 437934 892 437940 944
rect 437992 932 437998 944
rect 442626 932 442632 944
rect 437992 904 442632 932
rect 437992 892 437998 904
rect 442626 892 442632 904
rect 442684 892 442690 944
rect 483198 892 483204 944
rect 483256 932 483262 944
rect 488810 932 488816 944
rect 483256 904 488816 932
rect 483256 892 483262 904
rect 488810 892 488816 904
rect 488868 892 488874 944
rect 491202 892 491208 944
rect 491260 932 491266 944
rect 497090 932 497096 944
rect 491260 904 497096 932
rect 491260 892 491266 904
rect 497090 892 497096 904
rect 497148 892 497154 944
rect 347498 824 347504 876
rect 347556 864 347562 876
rect 350442 864 350448 876
rect 347556 836 350448 864
rect 347556 824 347562 836
rect 350442 824 350448 836
rect 350500 824 350506 876
rect 361390 824 361396 876
rect 361448 864 361454 876
rect 364610 864 364616 876
rect 361448 836 364616 864
rect 361448 824 361454 836
rect 364610 824 364616 836
rect 364668 824 364674 876
rect 368382 824 368388 876
rect 368440 864 368446 876
rect 371694 864 371700 876
rect 368440 836 371700 864
rect 368440 824 368446 836
rect 371694 824 371700 836
rect 371752 824 371758 876
rect 371786 824 371792 876
rect 371844 864 371850 876
rect 375282 864 375288 876
rect 371844 836 375288 864
rect 371844 824 371850 836
rect 375282 824 375288 836
rect 375340 824 375346 876
rect 384574 824 384580 876
rect 384632 864 384638 876
rect 388254 864 388260 876
rect 384632 836 388260 864
rect 384632 824 384638 836
rect 388254 824 388260 836
rect 388312 824 388318 876
rect 391566 824 391572 876
rect 391624 864 391630 876
rect 395338 864 395344 876
rect 391624 836 395344 864
rect 391624 824 391630 836
rect 395338 824 395344 836
rect 395396 824 395402 876
rect 396166 824 396172 876
rect 396224 864 396230 876
rect 400122 864 400128 876
rect 396224 836 400128 864
rect 396224 824 396230 836
rect 400122 824 400128 836
rect 400180 824 400186 876
rect 406654 824 406660 876
rect 406712 864 406718 876
rect 410794 864 410800 876
rect 406712 836 410800 864
rect 406712 824 406718 836
rect 410794 824 410800 836
rect 410852 824 410858 876
rect 417050 824 417056 876
rect 417108 864 417114 876
rect 421374 864 421380 876
rect 417108 836 421380 864
rect 417108 824 417114 836
rect 421374 824 421380 836
rect 421432 824 421438 876
rect 429838 824 429844 876
rect 429896 864 429902 876
rect 434438 864 434444 876
rect 429896 836 434444 864
rect 429896 824 429902 836
rect 434438 824 434444 836
rect 434496 824 434502 876
rect 443730 824 443736 876
rect 443788 864 443794 876
rect 448238 864 448244 876
rect 443788 836 448244 864
rect 443788 824 443794 836
rect 448238 824 448244 836
rect 448296 824 448302 876
rect 451826 824 451832 876
rect 451884 864 451890 876
rect 456518 864 456524 876
rect 451884 836 456524 864
rect 451884 824 451890 836
rect 456518 824 456524 836
rect 456576 824 456582 876
rect 463418 824 463424 876
rect 463476 864 463482 876
rect 468662 864 468668 876
rect 463476 836 468668 864
rect 463476 824 463482 836
rect 468662 824 468668 836
rect 468720 824 468726 876
rect 476206 824 476212 876
rect 476264 864 476270 876
rect 481358 864 481364 876
rect 476264 836 481364 864
rect 476264 824 476270 836
rect 481358 824 481364 836
rect 481416 824 481422 876
rect 434346 756 434352 808
rect 434404 796 434410 808
rect 439130 796 439136 808
rect 434404 768 439136 796
rect 434404 756 434410 768
rect 439130 756 439136 768
rect 439188 756 439194 808
rect 52546 688 52552 740
rect 52604 728 52610 740
rect 55030 728 55036 740
rect 52604 700 55036 728
rect 52604 688 52610 700
rect 55030 688 55036 700
rect 55088 688 55094 740
rect 59630 688 59636 740
rect 59688 728 59694 740
rect 61930 728 61936 740
rect 59688 700 61936 728
rect 59688 688 59694 700
rect 61930 688 61936 700
rect 61988 688 61994 740
rect 105722 688 105728 740
rect 105780 728 105786 740
rect 107286 728 107292 740
rect 105780 700 107292 728
rect 105780 688 105786 700
rect 107286 688 107292 700
rect 107344 688 107350 740
rect 274358 688 274364 740
rect 274416 728 274422 740
rect 276014 728 276020 740
rect 274416 700 276020 728
rect 274416 688 274422 700
rect 276014 688 276020 700
rect 276072 688 276078 740
rect 333514 688 333520 740
rect 333572 728 333578 740
rect 336274 728 336280 740
rect 333572 700 336280 728
rect 333572 688 333578 700
rect 336274 688 336280 700
rect 336332 688 336338 740
rect 338206 688 338212 740
rect 338264 728 338270 740
rect 340966 728 340972 740
rect 338264 700 340972 728
rect 338264 688 338270 700
rect 340966 688 340972 700
rect 341024 688 341030 740
rect 342806 688 342812 740
rect 342864 728 342870 740
rect 345750 728 345756 740
rect 342864 700 345756 728
rect 342864 688 342870 700
rect 345750 688 345756 700
rect 345808 688 345814 740
rect 346302 688 346308 740
rect 346360 728 346366 740
rect 349246 728 349252 740
rect 346360 700 349252 728
rect 346360 688 346366 700
rect 349246 688 349252 700
rect 349304 688 349310 740
rect 350902 688 350908 740
rect 350960 728 350966 740
rect 354030 728 354036 740
rect 350960 700 354036 728
rect 350960 688 350966 700
rect 354030 688 354036 700
rect 354088 688 354094 740
rect 365990 688 365996 740
rect 366048 728 366054 740
rect 369394 728 369400 740
rect 366048 700 369400 728
rect 366048 688 366054 700
rect 369394 688 369400 700
rect 369452 688 369458 740
rect 369486 688 369492 740
rect 369544 728 369550 740
rect 372890 728 372896 740
rect 369544 700 372896 728
rect 369544 688 369550 700
rect 372890 688 372896 700
rect 372948 688 372954 740
rect 541158 688 541164 740
rect 541216 728 541222 740
rect 547874 728 547880 740
rect 541216 700 547880 728
rect 541216 688 541222 700
rect 547874 688 547880 700
rect 547932 688 547938 740
rect 557534 688 557540 740
rect 557592 728 557598 740
rect 564434 728 564440 740
rect 557592 700 564440 728
rect 557592 688 557598 700
rect 564434 688 564440 700
rect 564492 688 564498 740
rect 553946 620 553952 672
rect 554004 660 554010 672
rect 554004 632 557534 660
rect 554004 620 554010 632
rect 69106 552 69112 604
rect 69164 592 69170 604
rect 71314 592 71320 604
rect 69164 564 71320 592
rect 69164 552 69170 564
rect 71314 552 71320 564
rect 71372 552 71378 604
rect 290642 552 290648 604
rect 290700 592 290706 604
rect 292574 592 292580 604
rect 290700 564 292580 592
rect 290700 552 290706 564
rect 292574 552 292580 564
rect 292632 552 292638 604
rect 304534 552 304540 604
rect 304592 592 304598 604
rect 306742 592 306748 604
rect 304592 564 306748 592
rect 304592 552 304598 564
rect 306742 552 306748 564
rect 306800 552 306806 604
rect 556246 552 556252 604
rect 556304 552 556310 604
rect 557506 592 557534 632
rect 563146 620 563152 672
rect 563204 660 563210 672
rect 570322 660 570328 672
rect 563204 632 570328 660
rect 563204 620 563210 632
rect 570322 620 570328 632
rect 570380 620 570386 672
rect 560846 592 560852 604
rect 557506 564 560852 592
rect 560846 552 560852 564
rect 560904 552 560910 604
rect 563238 552 563244 604
rect 563296 552 563302 604
rect 556264 524 556292 552
rect 563256 524 563284 552
rect 556264 496 563284 524
rect 507486 416 507492 468
rect 507544 456 507550 468
rect 513374 456 513380 468
rect 507544 428 513380 456
rect 507544 416 507550 428
rect 513374 416 513380 428
rect 513432 416 513438 468
rect 536558 416 536564 468
rect 536616 456 536622 468
rect 542814 456 542820 468
rect 536616 428 542820 456
rect 536616 416 536622 428
rect 542814 416 542820 428
rect 542872 416 542878 468
rect 544654 416 544660 468
rect 544712 456 544718 468
rect 551094 456 551100 468
rect 544712 428 551100 456
rect 544712 416 544718 428
rect 551094 416 551100 428
rect 551152 416 551158 468
rect 566642 416 566648 468
rect 566700 456 566706 468
rect 573726 456 573732 468
rect 566700 428 573732 456
rect 566700 416 566706 428
rect 573726 416 573732 428
rect 573784 416 573790 468
rect 383378 348 383384 400
rect 383436 388 383442 400
rect 386782 388 386788 400
rect 383436 360 386788 388
rect 383436 348 383442 360
rect 386782 348 386788 360
rect 386840 348 386846 400
rect 535362 348 535368 400
rect 535420 388 535426 400
rect 542170 388 542176 400
rect 535420 360 542176 388
rect 535420 348 535426 360
rect 542170 348 542176 360
rect 542228 348 542234 400
rect 546954 348 546960 400
rect 547012 388 547018 400
rect 553946 388 553952 400
rect 547012 360 553952 388
rect 547012 348 547018 360
rect 553946 348 553952 360
rect 554004 348 554010 400
rect 537662 280 537668 332
rect 537720 320 537726 332
rect 544562 320 544568 332
rect 537720 292 544568 320
rect 537720 280 537726 292
rect 544562 280 544568 292
rect 544620 280 544626 332
rect 545850 280 545856 332
rect 545908 320 545914 332
rect 552382 320 552388 332
rect 545908 292 552388 320
rect 545908 280 545914 292
rect 552382 280 552388 292
rect 552440 280 552446 332
rect 573634 280 573640 332
rect 573692 320 573698 332
rect 581178 320 581184 332
rect 573692 292 581184 320
rect 573692 280 573698 292
rect 581178 280 581184 292
rect 581236 280 581242 332
rect 392670 212 392676 264
rect 392728 252 392734 264
rect 396166 252 396172 264
rect 392728 224 396172 252
rect 392728 212 392734 224
rect 396166 212 396172 224
rect 396224 212 396230 264
rect 412450 212 412456 264
rect 412508 252 412514 264
rect 416866 252 416872 264
rect 412508 224 416872 252
rect 412508 212 412514 224
rect 416866 212 416872 224
rect 416924 212 416930 264
rect 421742 212 421748 264
rect 421800 252 421806 264
rect 425790 252 425796 264
rect 421800 224 425796 252
rect 421800 212 421806 224
rect 425790 212 425796 224
rect 425848 212 425854 264
rect 469306 212 469312 264
rect 469364 252 469370 264
rect 474182 252 474188 264
rect 469364 224 474188 252
rect 469364 212 469370 224
rect 474182 212 474188 224
rect 474240 212 474246 264
rect 508682 212 508688 264
rect 508740 252 508746 264
rect 514938 252 514944 264
rect 508740 224 514944 252
rect 508740 212 508746 224
rect 514938 212 514944 224
rect 514996 212 515002 264
rect 528462 212 528468 264
rect 528520 252 528526 264
rect 534534 252 534540 264
rect 528520 224 534540 252
rect 528520 212 528526 224
rect 534534 212 534540 224
rect 534592 212 534598 264
rect 564250 144 564256 196
rect 564308 184 564314 196
rect 571334 184 571340 196
rect 564308 156 571340 184
rect 564308 144 564314 156
rect 571334 144 571340 156
rect 571392 144 571398 196
rect 574830 144 574836 196
rect 574888 184 574894 196
rect 581822 184 581828 196
rect 574888 156 581828 184
rect 574888 144 574894 156
rect 581822 144 581828 156
rect 581880 144 581886 196
rect 431034 76 431040 128
rect 431092 116 431098 128
rect 435174 116 435180 128
rect 431092 88 435180 116
rect 431092 76 431098 88
rect 435174 76 435180 88
rect 435232 76 435238 128
rect 460014 76 460020 128
rect 460072 116 460078 128
rect 464982 116 464988 128
rect 460072 88 464988 116
rect 460072 76 460078 88
rect 464982 76 464988 88
rect 465040 76 465046 128
rect 470410 76 470416 128
rect 470468 116 470474 128
rect 475930 116 475936 128
rect 470468 88 475936 116
rect 470468 76 470474 88
rect 475930 76 475936 88
rect 475988 76 475994 128
rect 515674 76 515680 128
rect 515732 116 515738 128
rect 521654 116 521660 128
rect 515732 88 521660 116
rect 515732 76 515738 88
rect 521654 76 521660 88
rect 521712 76 521718 128
rect 524966 76 524972 128
rect 525024 116 525030 128
rect 531498 116 531504 128
rect 525024 88 531504 116
rect 525024 76 525030 88
rect 531498 76 531504 88
rect 531556 76 531562 128
rect 555142 76 555148 128
rect 555200 116 555206 128
rect 562226 116 562232 128
rect 555200 88 562232 116
rect 555200 76 555206 88
rect 562226 76 562232 88
rect 562284 76 562290 128
rect 565446 76 565452 128
rect 565504 116 565510 128
rect 572898 116 572904 128
rect 565504 88 572904 116
rect 565504 76 565510 88
rect 572898 76 572904 88
rect 572956 76 572962 128
rect 576118 76 576124 128
rect 576176 116 576182 128
rect 583570 116 583576 128
rect 576176 88 583576 116
rect 576176 76 576182 88
rect 583570 76 583576 88
rect 583628 76 583634 128
rect 354398 8 354404 60
rect 354456 48 354462 60
rect 357342 48 357348 60
rect 354456 20 357348 48
rect 354456 8 354462 20
rect 357342 8 357348 20
rect 357400 8 357406 60
rect 401962 8 401968 60
rect 402020 48 402026 60
rect 406194 48 406200 60
rect 402020 20 406200 48
rect 402020 8 402026 20
rect 406194 8 406200 20
rect 406252 8 406258 60
rect 499206 8 499212 60
rect 499264 48 499270 60
rect 505554 48 505560 60
rect 499264 20 505560 48
rect 499264 8 499270 20
rect 505554 8 505560 20
rect 505612 8 505618 60
rect 506290 8 506296 60
rect 506348 48 506354 60
rect 512086 48 512092 60
rect 506348 20 512092 48
rect 506348 8 506354 20
rect 512086 8 512092 20
rect 512144 8 512150 60
rect 516778 8 516784 60
rect 516836 48 516842 60
rect 523218 48 523224 60
rect 516836 20 523224 48
rect 516836 8 516842 20
rect 523218 8 523224 20
rect 523276 8 523282 60
rect 572530 8 572536 60
rect 572588 48 572594 60
rect 579614 48 579620 60
rect 572588 20 579620 48
rect 572588 8 572594 20
rect 579614 8 579620 20
rect 579672 8 579678 60
<< via1 >>
rect 102048 700748 102100 700800
rect 105452 700748 105504 700800
rect 200028 700748 200080 700800
rect 202788 700748 202840 700800
rect 314476 700748 314528 700800
rect 316316 700748 316368 700800
rect 53012 700544 53064 700596
rect 56784 700544 56836 700596
rect 151084 700544 151136 700596
rect 154120 700544 154172 700596
rect 412456 700408 412508 700460
rect 413652 700408 413704 700460
rect 363512 700340 363564 700392
rect 364984 700340 365036 700392
rect 20352 700204 20404 700256
rect 24308 700204 24360 700256
rect 36728 700204 36780 700256
rect 40500 700204 40552 700256
rect 69388 700204 69440 700256
rect 72976 700204 73028 700256
rect 85764 700204 85816 700256
rect 89168 700204 89220 700256
rect 134708 700204 134760 700256
rect 137836 700204 137888 700256
rect 167368 700204 167420 700256
rect 170312 700204 170364 700256
rect 183744 700204 183796 700256
rect 186504 700204 186556 700256
rect 232780 700204 232832 700256
rect 235172 700204 235224 700256
rect 249064 700204 249116 700256
rect 251456 700204 251508 700256
rect 265440 700204 265492 700256
rect 267648 700204 267700 700256
rect 281816 700204 281868 700256
rect 283840 700204 283892 700256
rect 330760 700204 330812 700256
rect 332508 700204 332560 700256
rect 347136 700204 347188 700256
rect 348792 700204 348844 700256
rect 396172 700204 396224 700256
rect 397460 700204 397512 700256
rect 428832 700204 428884 700256
rect 429844 700204 429896 700256
rect 445208 700204 445260 700256
rect 446128 700204 446180 700256
rect 461492 700204 461544 700256
rect 462320 700204 462372 700256
rect 118424 700136 118476 700188
rect 121644 700136 121696 700188
rect 216404 700136 216456 700188
rect 218980 700136 219032 700188
rect 298008 700136 298060 700188
rect 300124 700136 300176 700188
rect 477868 700136 477920 700188
rect 478512 700136 478564 700188
rect 494244 700136 494296 700188
rect 494796 700136 494848 700188
rect 379796 699864 379848 699916
rect 381176 699864 381228 699916
rect 576768 698232 576820 698284
rect 580172 698232 580224 698284
rect 4020 698164 4072 698216
rect 8116 698164 8168 698216
rect 578332 644512 578384 644564
rect 580908 644512 580960 644564
rect 578884 257796 578936 257848
rect 580908 257796 580960 257848
rect 578516 151444 578568 151496
rect 580908 151444 580960 151496
rect 578332 44956 578384 45008
rect 579988 44956 580040 45008
rect 576860 5516 576912 5568
rect 579620 5516 579672 5568
rect 11152 3884 11204 3936
rect 14508 3884 14560 3936
rect 14740 3884 14792 3936
rect 18004 3884 18056 3936
rect 20628 3884 20680 3936
rect 23800 3884 23852 3936
rect 24216 3884 24268 3936
rect 27296 3884 27348 3936
rect 27712 3884 27764 3936
rect 30700 3884 30752 3936
rect 32404 3884 32456 3936
rect 35392 3884 35444 3936
rect 38384 3884 38436 3936
rect 41188 3884 41240 3936
rect 43076 3884 43128 3936
rect 45788 3884 45840 3936
rect 46664 3884 46716 3936
rect 49284 3884 49336 3936
rect 50160 3884 50212 3936
rect 52780 3884 52832 3936
rect 56048 3884 56100 3936
rect 58576 3884 58628 3936
rect 72608 3884 72660 3936
rect 74860 3884 74912 3936
rect 247636 3884 247688 3936
rect 248604 3884 248656 3936
rect 285908 3884 285960 3936
rect 287796 3884 287848 3936
rect 1676 3816 1728 3868
rect 5216 3816 5268 3868
rect 13544 3816 13596 3868
rect 16808 3816 16860 3868
rect 19432 3816 19484 3868
rect 22604 3816 22656 3868
rect 23020 3816 23072 3868
rect 26100 3816 26152 3868
rect 26516 3816 26568 3868
rect 29596 3816 29648 3868
rect 30104 3816 30156 3868
rect 33092 3816 33144 3868
rect 33600 3816 33652 3868
rect 36588 3816 36640 3868
rect 37188 3816 37240 3868
rect 39992 3816 40044 3868
rect 41880 3816 41932 3868
rect 44684 3816 44736 3868
rect 45468 3816 45520 3868
rect 48180 3816 48232 3868
rect 48964 3816 49016 3868
rect 51584 3816 51636 3868
rect 53748 3816 53800 3868
rect 56276 3816 56328 3868
rect 57244 3816 57296 3868
rect 59772 3816 59824 3868
rect 71504 3816 71556 3868
rect 73664 3816 73716 3868
rect 78588 3816 78640 3868
rect 80656 3816 80708 3868
rect 80888 3816 80940 3868
rect 82956 3816 83008 3868
rect 87972 3816 88024 3868
rect 89948 3816 90000 3868
rect 96252 3816 96304 3868
rect 98044 3816 98096 3868
rect 244140 3816 244192 3868
rect 245200 3816 245252 3868
rect 256928 3816 256980 3868
rect 258264 3816 258316 3868
rect 259228 3816 259280 3868
rect 260656 3816 260708 3868
rect 261620 3816 261672 3868
rect 262956 3816 263008 3868
rect 263920 3816 263972 3868
rect 265348 3816 265400 3868
rect 268520 3816 268572 3868
rect 270040 3816 270092 3868
rect 270820 3816 270872 3868
rect 272432 3816 272484 3868
rect 275512 3816 275564 3868
rect 277124 3816 277176 3868
rect 277812 3816 277864 3868
rect 279516 3816 279568 3868
rect 284804 3816 284856 3868
rect 286600 3816 286652 3868
rect 292900 3816 292952 3868
rect 294880 3816 294932 3868
rect 299892 3816 299944 3868
rect 301964 3816 302016 3868
rect 306792 3816 306844 3868
rect 309048 3816 309100 3868
rect 572 3748 624 3800
rect 4112 3748 4164 3800
rect 7656 3748 7708 3800
rect 11012 3748 11064 3800
rect 12348 3748 12400 3800
rect 15704 3748 15756 3800
rect 15936 3748 15988 3800
rect 19108 3748 19160 3800
rect 21824 3748 21876 3800
rect 24904 3748 24956 3800
rect 25320 3748 25372 3800
rect 28400 3748 28452 3800
rect 31300 3748 31352 3800
rect 34196 3748 34248 3800
rect 34796 3748 34848 3800
rect 37692 3748 37744 3800
rect 40684 3748 40736 3800
rect 43488 3748 43540 3800
rect 44272 3748 44324 3800
rect 46984 3748 47036 3800
rect 47860 3748 47912 3800
rect 50480 3748 50532 3800
rect 51356 3748 51408 3800
rect 53976 3748 54028 3800
rect 54944 3748 54996 3800
rect 57380 3748 57432 3800
rect 58440 3748 58492 3800
rect 60876 3748 60928 3800
rect 64328 3748 64380 3800
rect 66672 3748 66724 3800
rect 67088 3748 67140 3800
rect 69064 3748 69116 3800
rect 70308 3748 70360 3800
rect 72468 3748 72520 3800
rect 73804 3748 73856 3800
rect 75964 3748 76016 3800
rect 79692 3748 79744 3800
rect 81760 3748 81812 3800
rect 86868 3748 86920 3800
rect 88752 3748 88804 3800
rect 95148 3748 95200 3800
rect 96848 3748 96900 3800
rect 103336 3748 103388 3800
rect 104944 3748 104996 3800
rect 216356 3748 216408 3800
rect 216864 3748 216916 3800
rect 222152 3748 222204 3800
rect 222752 3748 222804 3800
rect 224452 3748 224504 3800
rect 225144 3748 225196 3800
rect 230248 3748 230300 3800
rect 231032 3748 231084 3800
rect 231444 3748 231496 3800
rect 232228 3748 232280 3800
rect 232548 3748 232600 3800
rect 233424 3748 233476 3800
rect 233744 3748 233796 3800
rect 234620 3748 234672 3800
rect 237240 3748 237292 3800
rect 238116 3748 238168 3800
rect 238344 3748 238396 3800
rect 239312 3748 239364 3800
rect 239540 3748 239592 3800
rect 240508 3748 240560 3800
rect 240736 3748 240788 3800
rect 241704 3748 241756 3800
rect 241840 3748 241892 3800
rect 242900 3748 242952 3800
rect 245336 3748 245388 3800
rect 246396 3748 246448 3800
rect 246532 3748 246584 3800
rect 247592 3748 247644 3800
rect 250028 3748 250080 3800
rect 251180 3748 251232 3800
rect 252328 3748 252380 3800
rect 253480 3748 253532 3800
rect 255824 3748 255876 3800
rect 257068 3748 257120 3800
rect 258124 3748 258176 3800
rect 259460 3748 259512 3800
rect 260424 3748 260476 3800
rect 261760 3748 261812 3800
rect 262724 3748 262776 3800
rect 264152 3748 264204 3800
rect 265024 3748 265076 3800
rect 266544 3748 266596 3800
rect 267416 3748 267468 3800
rect 268844 3748 268896 3800
rect 269716 3748 269768 3800
rect 271236 3748 271288 3800
rect 272016 3748 272068 3800
rect 273628 3748 273680 3800
rect 276708 3748 276760 3800
rect 278320 3748 278372 3800
rect 279008 3748 279060 3800
rect 280712 3748 280764 3800
rect 283608 3748 283660 3800
rect 285404 3748 285456 3800
rect 287104 3748 287156 3800
rect 288992 3748 289044 3800
rect 291704 3748 291756 3800
rect 293684 3748 293736 3800
rect 294096 3748 294148 3800
rect 296076 3748 296128 3800
rect 298696 3748 298748 3800
rect 300768 3748 300820 3800
rect 300996 3748 301048 3800
rect 303160 3748 303212 3800
rect 307988 3748 308040 3800
rect 310244 3748 310296 3800
rect 316084 3748 316136 3800
rect 318524 3748 318576 3800
rect 323076 3748 323128 3800
rect 325608 3748 325660 3800
rect 6460 3000 6512 3052
rect 9864 3000 9916 3052
rect 63224 3000 63276 3052
rect 65524 3000 65576 3052
rect 18236 2864 18288 2916
rect 21456 2864 21508 2916
rect 253388 2864 253440 2916
rect 254676 2864 254728 2916
rect 4068 2796 4120 2848
rect 7472 2796 7524 2848
rect 9956 2796 10008 2848
rect 13268 2796 13320 2848
rect 17040 2796 17092 2848
rect 20260 2796 20312 2848
rect 28908 2796 28960 2848
rect 31852 2796 31904 2848
rect 35992 2796 36044 2848
rect 38844 2796 38896 2848
rect 39580 2796 39632 2848
rect 42340 2796 42392 2848
rect 62028 2796 62080 2848
rect 64420 2796 64472 2848
rect 65524 2796 65576 2848
rect 67824 2796 67876 2848
rect 248880 2796 248932 2848
rect 249984 2796 250036 2848
rect 251088 2796 251140 2848
rect 252376 2796 252428 2848
rect 254584 2796 254636 2848
rect 255872 2796 255924 2848
rect 309232 2796 309284 2848
rect 311440 2796 311492 2848
rect 315028 2796 315080 2848
rect 317328 2796 317380 2848
rect 411168 2796 411220 2848
rect 415492 2796 415544 2848
rect 440148 2796 440200 2848
rect 445024 2796 445076 2848
rect 449532 2796 449584 2848
rect 454500 2796 454552 2848
rect 478512 2796 478564 2848
rect 484032 2796 484084 2848
rect 3240 1300 3292 1352
rect 6368 1300 6420 1352
rect 60832 1300 60884 1352
rect 63316 1300 63368 1352
rect 67916 1300 67968 1352
rect 70124 1300 70176 1352
rect 76196 1300 76248 1352
rect 78220 1300 78272 1352
rect 83280 1300 83332 1352
rect 85212 1300 85264 1352
rect 85672 1300 85724 1352
rect 87512 1300 87564 1352
rect 89168 1300 89220 1352
rect 91008 1300 91060 1352
rect 91560 1300 91612 1352
rect 93308 1300 93360 1352
rect 93952 1300 94004 1352
rect 95700 1300 95752 1352
rect 97448 1300 97500 1352
rect 99104 1300 99156 1352
rect 101036 1300 101088 1352
rect 102600 1300 102652 1352
rect 104532 1300 104584 1352
rect 106096 1300 106148 1352
rect 106924 1300 106976 1352
rect 108396 1300 108448 1352
rect 109316 1300 109368 1352
rect 110696 1300 110748 1352
rect 112812 1300 112864 1352
rect 114192 1300 114244 1352
rect 116400 1300 116452 1352
rect 117688 1300 117740 1352
rect 119896 1300 119948 1352
rect 121184 1300 121236 1352
rect 125876 1300 125928 1352
rect 126980 1300 127032 1352
rect 129372 1300 129424 1352
rect 130476 1300 130528 1352
rect 130568 1300 130620 1352
rect 131580 1300 131632 1352
rect 131764 1300 131816 1352
rect 132776 1300 132828 1352
rect 132960 1300 133012 1352
rect 133972 1300 134024 1352
rect 137652 1300 137704 1352
rect 138572 1300 138624 1352
rect 144736 1300 144788 1352
rect 145564 1300 145616 1352
rect 145932 1300 145984 1352
rect 146668 1300 146720 1352
rect 148324 1300 148376 1352
rect 149060 1300 149112 1352
rect 154212 1300 154264 1352
rect 154856 1300 154908 1352
rect 162492 1300 162544 1352
rect 162952 1300 163004 1352
rect 266268 1300 266320 1352
rect 267740 1300 267792 1352
rect 273168 1300 273220 1352
rect 274824 1300 274876 1352
rect 280068 1300 280120 1352
rect 281908 1300 281960 1352
rect 282552 1300 282604 1352
rect 284300 1300 284352 1352
rect 288348 1300 288400 1352
rect 290188 1300 290240 1352
rect 295248 1300 295300 1352
rect 297272 1300 297324 1352
rect 297548 1300 297600 1352
rect 299664 1300 299716 1352
rect 302148 1300 302200 1352
rect 304356 1300 304408 1352
rect 305736 1300 305788 1352
rect 307944 1300 307996 1352
rect 310336 1300 310388 1352
rect 312636 1300 312688 1352
rect 313832 1300 313884 1352
rect 316224 1300 316276 1352
rect 317236 1300 317288 1352
rect 319720 1300 319772 1352
rect 321928 1300 321980 1352
rect 324412 1300 324464 1352
rect 325424 1300 325476 1352
rect 328000 1300 328052 1352
rect 328920 1300 328972 1352
rect 331588 1300 331640 1352
rect 332416 1300 332468 1352
rect 335084 1300 335136 1352
rect 335912 1300 335964 1352
rect 338672 1300 338724 1352
rect 339316 1300 339368 1352
rect 342168 1300 342220 1352
rect 345112 1300 345164 1352
rect 348056 1300 348108 1352
rect 349804 1300 349856 1352
rect 352840 1300 352892 1352
rect 353208 1300 353260 1352
rect 356336 1300 356388 1352
rect 356704 1300 356756 1352
rect 359924 1300 359976 1352
rect 362592 1300 362644 1352
rect 365812 1300 365864 1352
rect 367192 1300 367244 1352
rect 370596 1300 370648 1352
rect 370688 1300 370740 1352
rect 374092 1300 374144 1352
rect 376392 1300 376444 1352
rect 379980 1300 380032 1352
rect 385776 1300 385828 1352
rect 389456 1300 389508 1352
rect 395068 1300 395120 1352
rect 398932 1300 398984 1352
rect 399668 1300 399720 1352
rect 403624 1300 403676 1352
rect 405464 1300 405516 1352
rect 409604 1300 409656 1352
rect 415952 1300 416004 1352
rect 420184 1300 420236 1352
rect 427544 1300 427596 1352
rect 431868 1300 431920 1352
rect 433248 1300 433300 1352
rect 437848 1300 437900 1352
rect 442632 1300 442684 1352
rect 447416 1300 447468 1352
rect 448428 1300 448480 1352
rect 453304 1300 453356 1352
rect 458824 1300 458876 1352
rect 463976 1300 464028 1352
rect 468116 1300 468168 1352
rect 473084 1300 473136 1352
rect 480904 1300 480956 1352
rect 486424 1300 486476 1352
rect 487804 1300 487856 1352
rect 493140 1300 493192 1352
rect 497096 1300 497148 1352
rect 502984 1300 503036 1352
rect 504088 1300 504140 1352
rect 509700 1300 509752 1352
rect 509884 1300 509936 1352
rect 515772 1300 515824 1352
rect 519176 1300 519228 1352
rect 525432 1300 525484 1352
rect 526076 1300 526128 1352
rect 532148 1300 532200 1352
rect 534264 1300 534316 1352
rect 540428 1300 540480 1352
rect 542268 1300 542320 1352
rect 549076 1300 549128 1352
rect 551652 1300 551704 1352
rect 558552 1300 558604 1352
rect 560944 1300 560996 1352
rect 568028 1300 568080 1352
rect 571248 1300 571300 1352
rect 578608 1300 578660 1352
rect 75000 1232 75052 1284
rect 77116 1232 77168 1284
rect 77392 1232 77444 1284
rect 79416 1232 79468 1284
rect 82084 1232 82136 1284
rect 84016 1232 84068 1284
rect 84476 1232 84528 1284
rect 86408 1232 86460 1284
rect 90364 1232 90416 1284
rect 92204 1232 92256 1284
rect 92756 1232 92808 1284
rect 94504 1232 94556 1284
rect 98644 1232 98696 1284
rect 100300 1232 100352 1284
rect 102232 1232 102284 1284
rect 103796 1232 103848 1284
rect 108120 1232 108172 1284
rect 109592 1232 109644 1284
rect 110512 1232 110564 1284
rect 111892 1232 111944 1284
rect 115204 1232 115256 1284
rect 116584 1232 116636 1284
rect 117596 1232 117648 1284
rect 118884 1232 118936 1284
rect 122288 1232 122340 1284
rect 123484 1232 123536 1284
rect 124680 1232 124732 1284
rect 125784 1232 125836 1284
rect 128176 1232 128228 1284
rect 129280 1232 129332 1284
rect 136456 1232 136508 1284
rect 137376 1232 137428 1284
rect 138848 1232 138900 1284
rect 139768 1232 139820 1284
rect 140044 1232 140096 1284
rect 140872 1232 140924 1284
rect 281356 1232 281408 1284
rect 283104 1232 283156 1284
rect 289452 1232 289504 1284
rect 291384 1232 291436 1284
rect 296444 1232 296496 1284
rect 298468 1232 298520 1284
rect 303344 1232 303396 1284
rect 305552 1232 305604 1284
rect 312544 1232 312596 1284
rect 315028 1232 315080 1284
rect 318432 1232 318484 1284
rect 320916 1232 320968 1284
rect 324228 1232 324280 1284
rect 326804 1232 326856 1284
rect 330024 1232 330076 1284
rect 332692 1232 332744 1284
rect 334716 1232 334768 1284
rect 337476 1232 337528 1284
rect 340512 1232 340564 1284
rect 343364 1232 343416 1284
rect 344008 1232 344060 1284
rect 346952 1232 347004 1284
rect 348608 1232 348660 1284
rect 351644 1232 351696 1284
rect 352104 1232 352156 1284
rect 355232 1232 355284 1284
rect 355600 1232 355652 1284
rect 358728 1232 358780 1284
rect 359096 1232 359148 1284
rect 362316 1232 362368 1284
rect 363696 1232 363748 1284
rect 367008 1232 367060 1284
rect 372988 1232 373040 1284
rect 376484 1232 376536 1284
rect 377588 1232 377640 1284
rect 381176 1232 381228 1284
rect 388076 1232 388128 1284
rect 391848 1232 391900 1284
rect 393872 1232 393924 1284
rect 397736 1232 397788 1284
rect 398472 1232 398524 1284
rect 402520 1232 402572 1284
rect 403164 1232 403216 1284
rect 407212 1232 407264 1284
rect 410064 1232 410116 1284
rect 414296 1232 414348 1284
rect 418252 1232 418304 1284
rect 422576 1232 422628 1284
rect 424048 1232 424100 1284
rect 428464 1232 428516 1284
rect 435640 1232 435692 1284
rect 439964 1232 440016 1284
rect 444932 1232 444984 1284
rect 449808 1232 449860 1284
rect 450728 1232 450780 1284
rect 455696 1232 455748 1284
rect 456524 1232 456576 1284
rect 461584 1232 461636 1284
rect 462228 1232 462280 1284
rect 467472 1232 467524 1284
rect 471612 1232 471664 1284
rect 476580 1232 476632 1284
rect 479708 1232 479760 1284
rect 484860 1232 484912 1284
rect 489000 1232 489052 1284
rect 494704 1232 494756 1284
rect 498292 1232 498344 1284
rect 503812 1232 503864 1284
rect 510988 1232 511040 1284
rect 517152 1232 517204 1284
rect 517980 1232 518032 1284
rect 523868 1232 523920 1284
rect 527272 1232 527324 1284
rect 533712 1232 533764 1284
rect 543464 1232 543516 1284
rect 550272 1232 550324 1284
rect 550456 1232 550508 1284
rect 557356 1232 557408 1284
rect 562048 1232 562100 1284
rect 569132 1232 569184 1284
rect 570144 1232 570196 1284
rect 577412 1232 577464 1284
rect 99840 1164 99892 1216
rect 101496 1164 101548 1216
rect 114008 1164 114060 1216
rect 115388 1164 115440 1216
rect 311532 1164 311584 1216
rect 313832 1164 313884 1216
rect 319628 1164 319680 1216
rect 322112 1164 322164 1216
rect 326620 1164 326672 1216
rect 329196 1164 329248 1216
rect 331128 1164 331180 1216
rect 333888 1164 333940 1216
rect 337016 1164 337068 1216
rect 339868 1164 339920 1216
rect 341708 1164 341760 1216
rect 344560 1164 344612 1216
rect 357900 1164 357952 1216
rect 361120 1164 361172 1216
rect 364892 1164 364944 1216
rect 368204 1164 368256 1216
rect 375288 1164 375340 1216
rect 378876 1164 378928 1216
rect 381084 1164 381136 1216
rect 384764 1164 384816 1216
rect 390376 1164 390428 1216
rect 394240 1164 394292 1216
rect 400864 1164 400916 1216
rect 404820 1164 404872 1216
rect 407764 1164 407816 1216
rect 411904 1164 411956 1216
rect 413560 1164 413612 1216
rect 417884 1164 417936 1216
rect 419356 1164 419408 1216
rect 423404 1164 423456 1216
rect 426348 1164 426400 1216
rect 430856 1164 430908 1216
rect 441436 1164 441488 1216
rect 445852 1164 445904 1216
rect 446036 1164 446088 1216
rect 450912 1164 450964 1216
rect 457628 1164 457680 1216
rect 462412 1164 462464 1216
rect 465816 1164 465868 1216
rect 470692 1164 470744 1216
rect 475108 1164 475160 1216
rect 480536 1164 480588 1216
rect 482008 1164 482060 1216
rect 487252 1164 487304 1216
rect 492496 1164 492548 1216
rect 498200 1164 498252 1216
rect 505192 1164 505244 1216
rect 511264 1164 511316 1216
rect 513288 1164 513340 1216
rect 519544 1164 519596 1216
rect 522672 1164 522724 1216
rect 529020 1164 529072 1216
rect 531872 1164 531924 1216
rect 538404 1164 538456 1216
rect 540060 1164 540112 1216
rect 546684 1164 546736 1216
rect 548156 1164 548208 1216
rect 554964 1164 555016 1216
rect 558460 1164 558512 1216
rect 565636 1164 565688 1216
rect 569040 1164 569092 1216
rect 576308 1164 576360 1216
rect 5632 1096 5684 1148
rect 8668 1096 8720 1148
rect 111616 1096 111668 1148
rect 113088 1096 113140 1148
rect 123484 1096 123536 1148
rect 124772 1096 124824 1148
rect 320824 1096 320876 1148
rect 323308 1096 323360 1148
rect 327724 1096 327776 1148
rect 330392 1096 330444 1148
rect 360108 1096 360160 1148
rect 363512 1096 363564 1148
rect 382188 1096 382240 1148
rect 385960 1096 386012 1148
rect 389272 1096 389324 1148
rect 393044 1096 393096 1148
rect 397368 1096 397420 1148
rect 401324 1096 401376 1148
rect 404268 1096 404320 1148
rect 408408 1096 408460 1148
rect 408960 1096 409012 1148
rect 413100 1096 413152 1148
rect 420552 1096 420604 1148
rect 424968 1096 425020 1148
rect 428648 1096 428700 1148
rect 433248 1096 433300 1148
rect 436744 1096 436796 1148
rect 441528 1096 441580 1148
rect 454224 1096 454276 1148
rect 459192 1096 459244 1148
rect 461124 1096 461176 1148
rect 466276 1096 466328 1148
rect 472716 1096 472768 1148
rect 478144 1096 478196 1148
rect 486700 1096 486752 1148
rect 492312 1096 492364 1148
rect 493600 1096 493652 1148
rect 499396 1096 499448 1148
rect 500500 1096 500552 1148
rect 506480 1096 506532 1148
rect 512184 1096 512236 1148
rect 517980 1096 518032 1148
rect 523776 1096 523828 1148
rect 530124 1096 530176 1148
rect 530768 1096 530820 1148
rect 537208 1096 537260 1148
rect 538864 1096 538916 1148
rect 545488 1096 545540 1148
rect 552756 1096 552808 1148
rect 559748 1096 559800 1148
rect 567844 1096 567896 1148
rect 575112 1096 575164 1148
rect 378784 1028 378836 1080
rect 382372 1028 382424 1080
rect 386880 1028 386932 1080
rect 390652 1028 390704 1080
rect 425152 1028 425204 1080
rect 429660 1028 429712 1080
rect 439136 1028 439188 1080
rect 443828 1028 443880 1080
rect 447232 1028 447284 1080
rect 452108 1028 452160 1080
rect 455328 1028 455380 1080
rect 460112 1028 460164 1080
rect 466920 1028 466972 1080
rect 472256 1028 472308 1080
rect 477408 1028 477460 1080
rect 482468 1028 482520 1080
rect 485504 1028 485556 1080
rect 490748 1028 490800 1080
rect 494796 1028 494848 1080
rect 500592 1028 500644 1080
rect 501696 1028 501748 1080
rect 507308 1028 507360 1080
rect 514484 1028 514536 1080
rect 520740 1028 520792 1080
rect 521476 1028 521528 1080
rect 527824 1028 527876 1080
rect 529572 1028 529624 1080
rect 536104 1028 536156 1080
rect 549352 1028 549404 1080
rect 556160 1028 556212 1080
rect 559656 1028 559708 1080
rect 566832 1028 566884 1080
rect 374184 960 374236 1012
rect 377680 960 377732 1012
rect 379888 960 379940 1012
rect 383568 960 383620 1012
rect 414756 960 414808 1012
rect 418988 960 419040 1012
rect 422852 960 422904 1012
rect 427268 960 427320 1012
rect 432144 960 432196 1012
rect 436744 960 436796 1012
rect 453028 960 453080 1012
rect 458088 960 458140 1012
rect 464620 960 464672 1012
rect 469864 960 469916 1012
rect 473912 960 473964 1012
rect 479340 960 479392 1012
rect 484308 960 484360 1012
rect 489920 960 489972 1012
rect 490104 960 490156 1012
rect 495532 960 495584 1012
rect 495992 960 496044 1012
rect 501788 960 501840 1012
rect 502892 960 502944 1012
rect 508872 960 508924 1012
rect 520188 960 520240 1012
rect 526628 960 526680 1012
rect 533068 960 533120 1012
rect 539600 960 539652 1012
rect 8760 892 8812 944
rect 12164 892 12216 944
rect 121092 892 121144 944
rect 122380 892 122432 944
rect 437940 892 437992 944
rect 442632 892 442684 944
rect 483204 892 483256 944
rect 488816 892 488868 944
rect 491208 892 491260 944
rect 497096 892 497148 944
rect 347504 824 347556 876
rect 350448 824 350500 876
rect 361396 824 361448 876
rect 364616 824 364668 876
rect 368388 824 368440 876
rect 371700 824 371752 876
rect 371792 824 371844 876
rect 375288 824 375340 876
rect 384580 824 384632 876
rect 388260 824 388312 876
rect 391572 824 391624 876
rect 395344 824 395396 876
rect 396172 824 396224 876
rect 400128 824 400180 876
rect 406660 824 406712 876
rect 410800 824 410852 876
rect 417056 824 417108 876
rect 421380 824 421432 876
rect 429844 824 429896 876
rect 434444 824 434496 876
rect 443736 824 443788 876
rect 448244 824 448296 876
rect 451832 824 451884 876
rect 456524 824 456576 876
rect 463424 824 463476 876
rect 468668 824 468720 876
rect 476212 824 476264 876
rect 481364 824 481416 876
rect 434352 756 434404 808
rect 439136 756 439188 808
rect 52552 688 52604 740
rect 55036 688 55088 740
rect 59636 688 59688 740
rect 61936 688 61988 740
rect 105728 688 105780 740
rect 107292 688 107344 740
rect 274364 688 274416 740
rect 276020 688 276072 740
rect 333520 688 333572 740
rect 336280 688 336332 740
rect 338212 688 338264 740
rect 340972 688 341024 740
rect 342812 688 342864 740
rect 345756 688 345808 740
rect 346308 688 346360 740
rect 349252 688 349304 740
rect 350908 688 350960 740
rect 354036 688 354088 740
rect 365996 688 366048 740
rect 369400 688 369452 740
rect 369492 688 369544 740
rect 372896 688 372948 740
rect 541164 688 541216 740
rect 547880 688 547932 740
rect 557540 688 557592 740
rect 564440 688 564492 740
rect 553952 620 554004 672
rect 69112 552 69164 604
rect 71320 552 71372 604
rect 290648 552 290700 604
rect 292580 552 292632 604
rect 304540 552 304592 604
rect 306748 552 306800 604
rect 556252 552 556304 604
rect 563152 620 563204 672
rect 570328 620 570380 672
rect 560852 552 560904 604
rect 563244 552 563296 604
rect 507492 416 507544 468
rect 513380 416 513432 468
rect 536564 416 536616 468
rect 542820 416 542872 468
rect 544660 416 544712 468
rect 551100 416 551152 468
rect 566648 416 566700 468
rect 573732 416 573784 468
rect 383384 348 383436 400
rect 386788 348 386840 400
rect 535368 348 535420 400
rect 542176 348 542228 400
rect 546960 348 547012 400
rect 553952 348 554004 400
rect 537668 280 537720 332
rect 544568 280 544620 332
rect 545856 280 545908 332
rect 552388 280 552440 332
rect 573640 280 573692 332
rect 581184 280 581236 332
rect 392676 212 392728 264
rect 396172 212 396224 264
rect 412456 212 412508 264
rect 416872 212 416924 264
rect 421748 212 421800 264
rect 425796 212 425848 264
rect 469312 212 469364 264
rect 474188 212 474240 264
rect 508688 212 508740 264
rect 514944 212 514996 264
rect 528468 212 528520 264
rect 534540 212 534592 264
rect 564256 144 564308 196
rect 571340 144 571392 196
rect 574836 144 574888 196
rect 581828 144 581880 196
rect 431040 76 431092 128
rect 435180 76 435232 128
rect 460020 76 460072 128
rect 464988 76 465040 128
rect 470416 76 470468 128
rect 475936 76 475988 128
rect 515680 76 515732 128
rect 521660 76 521712 128
rect 524972 76 525024 128
rect 531504 76 531556 128
rect 555148 76 555200 128
rect 562232 76 562284 128
rect 565452 76 565504 128
rect 572904 76 572956 128
rect 576124 76 576176 128
rect 583576 76 583628 128
rect 354404 8 354456 60
rect 357348 8 357400 60
rect 401968 8 402020 60
rect 406200 8 406252 60
rect 499212 8 499264 60
rect 505560 8 505612 60
rect 506296 8 506348 60
rect 512092 8 512144 60
rect 516784 8 516836 60
rect 523224 8 523276 60
rect 572536 8 572588 60
rect 579620 8 579672 60
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510632 703582 510844 703610
rect 8128 698222 8156 703520
rect 24320 700262 24348 703520
rect 40512 700262 40540 703520
rect 56796 700602 56824 703520
rect 53012 700596 53064 700602
rect 53012 700538 53064 700544
rect 56784 700596 56836 700602
rect 56784 700538 56836 700544
rect 20352 700256 20404 700262
rect 20352 700198 20404 700204
rect 24308 700256 24360 700262
rect 24308 700198 24360 700204
rect 36728 700256 36780 700262
rect 36728 700198 36780 700204
rect 40500 700256 40552 700262
rect 40500 700198 40552 700204
rect 4020 698216 4072 698222
rect 4020 698158 4072 698164
rect 8116 698216 8168 698222
rect 20364 698170 20392 700198
rect 36740 698170 36768 700198
rect 53024 698170 53052 700538
rect 72988 700262 73016 703520
rect 89180 700262 89208 703520
rect 105464 700806 105492 703520
rect 102048 700800 102100 700806
rect 102048 700742 102100 700748
rect 105452 700800 105504 700806
rect 105452 700742 105504 700748
rect 69388 700256 69440 700262
rect 69388 700198 69440 700204
rect 72976 700256 73028 700262
rect 72976 700198 73028 700204
rect 85764 700256 85816 700262
rect 85764 700198 85816 700204
rect 89168 700256 89220 700262
rect 89168 700198 89220 700204
rect 69400 698170 69428 700198
rect 85776 698170 85804 700198
rect 102060 698170 102088 700742
rect 121656 700194 121684 703520
rect 137848 700262 137876 703520
rect 154132 700602 154160 703520
rect 151084 700596 151136 700602
rect 151084 700538 151136 700544
rect 154120 700596 154172 700602
rect 154120 700538 154172 700544
rect 134708 700256 134760 700262
rect 134708 700198 134760 700204
rect 137836 700256 137888 700262
rect 137836 700198 137888 700204
rect 118424 700188 118476 700194
rect 118424 700130 118476 700136
rect 121644 700188 121696 700194
rect 121644 700130 121696 700136
rect 118436 698170 118464 700130
rect 134720 698170 134748 700198
rect 151096 698170 151124 700538
rect 170324 700262 170352 703520
rect 186516 700262 186544 703520
rect 202800 700806 202828 703520
rect 200028 700800 200080 700806
rect 200028 700742 200080 700748
rect 202788 700800 202840 700806
rect 202788 700742 202840 700748
rect 167368 700256 167420 700262
rect 167368 700198 167420 700204
rect 170312 700256 170364 700262
rect 170312 700198 170364 700204
rect 183744 700256 183796 700262
rect 183744 700198 183796 700204
rect 186504 700256 186556 700262
rect 186504 700198 186556 700204
rect 167380 698170 167408 700198
rect 183756 698170 183784 700198
rect 8116 698158 8168 698164
rect 3514 697976 3570 697985
rect 4032 697959 4060 698158
rect 20316 698142 20392 698170
rect 36692 698142 36768 698170
rect 52976 698142 53052 698170
rect 69352 698142 69428 698170
rect 85728 698142 85804 698170
rect 102012 698142 102088 698170
rect 118388 698142 118464 698170
rect 134672 698142 134748 698170
rect 151048 698142 151124 698170
rect 167332 698142 167408 698170
rect 183708 698142 183784 698170
rect 200040 698170 200068 700742
rect 218992 700194 219020 703520
rect 235184 700262 235212 703520
rect 251468 700262 251496 703520
rect 267660 700262 267688 703520
rect 283852 700262 283880 703520
rect 232780 700256 232832 700262
rect 232780 700198 232832 700204
rect 235172 700256 235224 700262
rect 235172 700198 235224 700204
rect 249064 700256 249116 700262
rect 249064 700198 249116 700204
rect 251456 700256 251508 700262
rect 251456 700198 251508 700204
rect 265440 700256 265492 700262
rect 265440 700198 265492 700204
rect 267648 700256 267700 700262
rect 267648 700198 267700 700204
rect 281816 700256 281868 700262
rect 281816 700198 281868 700204
rect 283840 700256 283892 700262
rect 283840 700198 283892 700204
rect 216404 700188 216456 700194
rect 216404 700130 216456 700136
rect 218980 700188 219032 700194
rect 218980 700130 219032 700136
rect 216416 698170 216444 700130
rect 232792 698170 232820 700198
rect 249076 698170 249104 700198
rect 265452 698170 265480 700198
rect 281828 698170 281856 700198
rect 300136 700194 300164 703520
rect 316328 700806 316356 703520
rect 314476 700800 314528 700806
rect 314476 700742 314528 700748
rect 316316 700800 316368 700806
rect 316316 700742 316368 700748
rect 298008 700188 298060 700194
rect 298008 700130 298060 700136
rect 300124 700188 300176 700194
rect 300124 700130 300176 700136
rect 200040 698142 200112 698170
rect 20316 697959 20344 698142
rect 36692 697959 36720 698142
rect 52976 697959 53004 698142
rect 69352 697959 69380 698142
rect 85728 697959 85756 698142
rect 102012 697959 102040 698142
rect 118388 697959 118416 698142
rect 134672 697959 134700 698142
rect 151048 697959 151076 698142
rect 167332 697959 167360 698142
rect 183708 697959 183736 698142
rect 200084 697959 200112 698142
rect 216368 698142 216444 698170
rect 232744 698142 232820 698170
rect 249028 698142 249104 698170
rect 265404 698142 265480 698170
rect 281780 698142 281856 698170
rect 298020 698170 298048 700130
rect 314488 698170 314516 700742
rect 332520 700262 332548 703520
rect 348804 700262 348832 703520
rect 364996 700398 365024 703520
rect 363512 700392 363564 700398
rect 363512 700334 363564 700340
rect 364984 700392 365036 700398
rect 364984 700334 365036 700340
rect 330760 700256 330812 700262
rect 330760 700198 330812 700204
rect 332508 700256 332560 700262
rect 332508 700198 332560 700204
rect 347136 700256 347188 700262
rect 347136 700198 347188 700204
rect 348792 700256 348844 700262
rect 348792 700198 348844 700204
rect 330772 698170 330800 700198
rect 347148 698170 347176 700198
rect 363524 698170 363552 700334
rect 381188 699922 381216 703520
rect 397472 700262 397500 703520
rect 413664 700466 413692 703520
rect 412456 700460 412508 700466
rect 412456 700402 412508 700408
rect 413652 700460 413704 700466
rect 413652 700402 413704 700408
rect 396172 700256 396224 700262
rect 396172 700198 396224 700204
rect 397460 700256 397512 700262
rect 397460 700198 397512 700204
rect 379796 699916 379848 699922
rect 379796 699858 379848 699864
rect 381176 699916 381228 699922
rect 381176 699858 381228 699864
rect 379808 698170 379836 699858
rect 396184 698170 396212 700198
rect 412468 698170 412496 700402
rect 429856 700262 429884 703520
rect 446140 700262 446168 703520
rect 462332 700262 462360 703520
rect 428832 700256 428884 700262
rect 428832 700198 428884 700204
rect 429844 700256 429896 700262
rect 429844 700198 429896 700204
rect 445208 700256 445260 700262
rect 445208 700198 445260 700204
rect 446128 700256 446180 700262
rect 446128 700198 446180 700204
rect 461492 700256 461544 700262
rect 461492 700198 461544 700204
rect 462320 700256 462372 700262
rect 462320 700198 462372 700204
rect 428844 698170 428872 700198
rect 445220 698170 445248 700198
rect 461504 698170 461532 700198
rect 478524 700194 478552 703520
rect 494808 700194 494836 703520
rect 477868 700188 477920 700194
rect 477868 700130 477920 700136
rect 478512 700188 478564 700194
rect 478512 700130 478564 700136
rect 494244 700188 494296 700194
rect 494244 700130 494296 700136
rect 494796 700188 494848 700194
rect 494796 700130 494848 700136
rect 477880 698170 477908 700130
rect 494256 698170 494284 700130
rect 510632 699802 510660 703582
rect 510816 703474 510844 703582
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 511000 703474 511028 703520
rect 510816 703446 511028 703474
rect 527192 699802 527220 703520
rect 543476 702434 543504 703520
rect 559668 702434 559696 703520
rect 510540 699774 510660 699802
rect 526916 699774 527220 699802
rect 543200 702406 543504 702434
rect 559576 702406 559696 702434
rect 510540 698170 510568 699774
rect 526916 698170 526944 699774
rect 543200 698170 543228 702406
rect 559576 698170 559604 702406
rect 298020 698142 298092 698170
rect 216368 697959 216396 698142
rect 232744 697959 232772 698142
rect 249028 697959 249056 698142
rect 265404 697959 265432 698142
rect 281780 697959 281808 698142
rect 298064 697959 298092 698142
rect 314440 698142 314516 698170
rect 330724 698142 330800 698170
rect 347100 698142 347176 698170
rect 363476 698142 363552 698170
rect 379760 698142 379836 698170
rect 396136 698142 396212 698170
rect 412420 698142 412496 698170
rect 428796 698142 428872 698170
rect 445172 698142 445248 698170
rect 461456 698142 461532 698170
rect 477832 698142 477908 698170
rect 494208 698142 494284 698170
rect 510492 698142 510568 698170
rect 526868 698142 526944 698170
rect 543152 698142 543228 698170
rect 559528 698142 559604 698170
rect 575860 698170 575888 703520
rect 576768 698284 576820 698290
rect 576768 698226 576820 698232
rect 580172 698284 580224 698290
rect 580172 698226 580224 698232
rect 576780 698193 576808 698226
rect 576766 698184 576822 698193
rect 575860 698142 575932 698170
rect 314440 697959 314468 698142
rect 330724 697959 330752 698142
rect 347100 697959 347128 698142
rect 363476 697959 363504 698142
rect 379760 697959 379788 698142
rect 396136 697959 396164 698142
rect 412420 697959 412448 698142
rect 428796 697959 428824 698142
rect 445172 697959 445200 698142
rect 461456 697959 461484 698142
rect 477832 697959 477860 698142
rect 494208 697959 494236 698142
rect 510492 697959 510520 698142
rect 526868 697959 526896 698142
rect 543152 697959 543180 698142
rect 559528 697959 559556 698142
rect 575904 697959 575932 698142
rect 576766 698119 576822 698128
rect 3514 697911 3570 697920
rect 3528 697377 3556 697911
rect 3514 697368 3570 697377
rect 3514 697303 3570 697312
rect 580184 697241 580212 698226
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 579526 684720 579582 684729
rect 579582 684678 579660 684706
rect 579526 684655 579582 684664
rect 579632 683913 579660 684678
rect 579618 683904 579674 683913
rect 579618 683839 579674 683848
rect 578330 644600 578386 644609
rect 578330 644535 578332 644544
rect 578384 644535 578386 644544
rect 580908 644564 580960 644570
rect 578332 644506 578384 644512
rect 580908 644506 580960 644512
rect 580920 644065 580948 644506
rect 580906 644056 580962 644065
rect 580906 643991 580962 644000
rect 3422 436656 3478 436665
rect 3422 436591 3478 436600
rect 3436 436051 3464 436591
rect 3422 436042 3478 436051
rect 3422 435977 3478 435986
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3436 422997 3464 423535
rect 3422 422988 3478 422997
rect 3422 422923 3478 422932
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 3436 409943 3464 410479
rect 3422 409934 3478 409943
rect 3422 409869 3478 409878
rect 3422 397488 3478 397497
rect 3422 397423 3478 397432
rect 3436 396889 3464 397423
rect 3422 396880 3478 396889
rect 3422 396815 3478 396824
rect 3422 384432 3478 384441
rect 3422 384367 3478 384376
rect 3436 383713 3464 384367
rect 3422 383704 3478 383713
rect 3422 383639 3478 383648
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 3436 370659 3464 371311
rect 3422 370650 3478 370659
rect 3422 370585 3478 370594
rect 3422 358456 3478 358465
rect 3422 358391 3478 358400
rect 3436 357605 3464 358391
rect 3422 357596 3478 357605
rect 3422 357531 3478 357540
rect 579526 351928 579582 351937
rect 579526 351863 579582 351872
rect 579540 351121 579568 351863
rect 579526 351112 579582 351121
rect 579526 351047 579582 351056
rect 3422 345400 3478 345409
rect 3422 345335 3478 345344
rect 3436 344429 3464 345335
rect 3422 344420 3478 344429
rect 3422 344355 3478 344364
rect 579618 338600 579674 338609
rect 579618 338535 579674 338544
rect 579526 337920 579582 337929
rect 579632 337906 579660 338535
rect 579582 337878 579660 337906
rect 579526 337855 579582 337864
rect 3422 332344 3478 332353
rect 3422 332279 3478 332288
rect 3436 331375 3464 332279
rect 3422 331366 3478 331375
rect 3422 331301 3478 331310
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324465 580212 325207
rect 580170 324456 580226 324465
rect 580170 324391 580226 324400
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 318321 3464 319223
rect 3422 318312 3478 318321
rect 3422 318247 3478 318256
rect 579618 312080 579674 312089
rect 579618 312015 579674 312024
rect 579526 311128 579582 311137
rect 579632 311114 579660 312015
rect 579582 311086 579660 311114
rect 579526 311063 579582 311072
rect 3422 306232 3478 306241
rect 3422 306167 3478 306176
rect 3436 305145 3464 306167
rect 3422 305136 3478 305145
rect 3422 305071 3478 305080
rect 579618 298752 579674 298761
rect 579618 298687 579674 298696
rect 579526 297800 579582 297809
rect 579632 297786 579660 298687
rect 579582 297758 579660 297786
rect 579526 297735 579582 297744
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 3436 292091 3464 293111
rect 3422 292082 3478 292091
rect 3422 292017 3478 292026
rect 580170 285424 580226 285433
rect 580170 285359 580226 285368
rect 580184 284481 580212 285359
rect 580170 284472 580226 284481
rect 580170 284407 580226 284416
rect 3422 280120 3478 280129
rect 3422 280055 3478 280064
rect 3436 279037 3464 280055
rect 3422 279028 3478 279037
rect 3422 278963 3478 278972
rect 579618 272232 579674 272241
rect 579618 272167 579674 272176
rect 579526 271144 579582 271153
rect 579632 271130 579660 272167
rect 579582 271102 579660 271130
rect 579526 271079 579582 271088
rect 3422 267200 3478 267209
rect 3422 267135 3478 267144
rect 3436 265983 3464 267135
rect 3422 265974 3478 265983
rect 3422 265909 3478 265918
rect 580906 258904 580962 258913
rect 580906 258839 580962 258848
rect 580920 257854 580948 258839
rect 578884 257848 578936 257854
rect 578884 257790 578936 257796
rect 580908 257848 580960 257854
rect 580908 257790 580960 257796
rect 578896 257689 578924 257790
rect 578882 257680 578938 257689
rect 578882 257615 578938 257624
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3436 252807 3464 254079
rect 3422 252798 3478 252807
rect 3422 252733 3478 252742
rect 580170 245576 580226 245585
rect 580170 245511 580226 245520
rect 580184 244497 580212 245511
rect 580170 244488 580226 244497
rect 580170 244423 580226 244432
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 3436 239753 3464 241023
rect 3422 239744 3478 239753
rect 3422 239679 3478 239688
rect 579618 232384 579674 232393
rect 579618 232319 579674 232328
rect 579526 231160 579582 231169
rect 579632 231146 579660 232319
rect 579582 231118 579660 231146
rect 579526 231095 579582 231104
rect 3422 228032 3478 228041
rect 3422 227967 3478 227976
rect 3436 226699 3464 227967
rect 3422 226690 3478 226699
rect 3422 226625 3478 226634
rect 579618 219056 579674 219065
rect 579618 218991 579674 219000
rect 579526 217696 579582 217705
rect 579632 217682 579660 218991
rect 579582 217654 579660 217682
rect 579526 217631 579582 217640
rect 3422 214976 3478 214985
rect 3422 214911 3478 214920
rect 3436 213523 3464 214911
rect 3422 213514 3478 213523
rect 3422 213449 3478 213458
rect 579618 205728 579674 205737
rect 579618 205663 579674 205672
rect 579526 204368 579582 204377
rect 579632 204354 579660 205663
rect 579582 204326 579660 204354
rect 579526 204303 579582 204312
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 3436 200469 3464 201855
rect 3422 200460 3478 200469
rect 3422 200395 3478 200404
rect 579618 192536 579674 192545
rect 579618 192471 579674 192480
rect 579526 191040 579582 191049
rect 579632 191026 579660 192471
rect 579582 190998 579660 191026
rect 579526 190975 579582 190984
rect 3606 188864 3662 188873
rect 3606 188799 3662 188808
rect 3620 187415 3648 188799
rect 3606 187406 3662 187415
rect 3606 187341 3662 187350
rect 579618 179208 579674 179217
rect 579618 179143 579674 179152
rect 579526 177712 579582 177721
rect 579632 177698 579660 179143
rect 579582 177670 579660 177698
rect 579526 177647 579582 177656
rect 3422 175944 3478 175953
rect 3422 175879 3478 175888
rect 3436 174239 3464 175879
rect 3422 174230 3478 174239
rect 3422 174165 3478 174174
rect 579618 165880 579674 165889
rect 579618 165815 579674 165824
rect 579526 164384 579582 164393
rect 579632 164370 579660 165815
rect 579582 164342 579660 164370
rect 579526 164319 579582 164328
rect 2134 162888 2190 162897
rect 2134 162823 2190 162832
rect 2148 161129 2176 162823
rect 2134 161120 2190 161129
rect 2134 161055 2190 161064
rect 580906 152688 580962 152697
rect 580906 152623 580962 152632
rect 580920 151502 580948 152623
rect 578516 151496 578568 151502
rect 578516 151438 578568 151444
rect 580908 151496 580960 151502
rect 580908 151438 580960 151444
rect 578528 151065 578556 151438
rect 578514 151056 578570 151065
rect 578514 150991 578570 151000
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3436 148131 3464 149767
rect 3422 148122 3478 148131
rect 3422 148057 3478 148066
rect 579618 139360 579674 139369
rect 579618 139295 579674 139304
rect 579526 137592 579582 137601
rect 579632 137578 579660 139295
rect 579582 137550 579660 137578
rect 579526 137527 579582 137536
rect 2134 136776 2190 136785
rect 2134 136711 2190 136720
rect 2148 135017 2176 136711
rect 2134 135008 2190 135017
rect 2134 134943 2190 134952
rect 579618 126032 579674 126041
rect 579618 125967 579674 125976
rect 579526 124400 579582 124409
rect 579632 124386 579660 125967
rect 579582 124358 579660 124386
rect 579526 124335 579582 124344
rect 3422 123720 3478 123729
rect 3422 123655 3478 123664
rect 3436 121901 3464 123655
rect 3422 121892 3478 121901
rect 3422 121827 3478 121836
rect 579618 112840 579674 112849
rect 579618 112775 579674 112784
rect 579526 110936 579582 110945
rect 579632 110922 579660 112775
rect 579582 110894 579660 110922
rect 579526 110871 579582 110880
rect 2134 110664 2190 110673
rect 2134 110599 2190 110608
rect 2148 108905 2176 110599
rect 2134 108896 2190 108905
rect 2134 108831 2190 108840
rect 579618 99512 579674 99521
rect 579618 99447 579674 99456
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 579526 97608 579582 97617
rect 579632 97594 579660 99447
rect 579582 97566 579660 97594
rect 579526 97543 579582 97552
rect 3436 95793 3464 97543
rect 3422 95784 3478 95793
rect 3422 95719 3478 95728
rect 579618 86184 579674 86193
rect 579618 86119 579674 86128
rect 2134 84688 2190 84697
rect 2134 84623 2190 84632
rect 2148 82657 2176 84623
rect 579526 84280 579582 84289
rect 579632 84266 579660 86119
rect 579582 84238 579660 84266
rect 579526 84215 579582 84224
rect 2134 82648 2190 82657
rect 2134 82583 2190 82592
rect 579618 72992 579674 73001
rect 579618 72927 579674 72936
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3436 69563 3464 71567
rect 579526 70952 579582 70961
rect 579632 70938 579660 72927
rect 579582 70910 579660 70938
rect 579526 70887 579582 70896
rect 3422 69554 3478 69563
rect 3422 69489 3478 69498
rect 579618 59664 579674 59673
rect 579618 59599 579674 59608
rect 2134 58576 2190 58585
rect 2134 58511 2190 58520
rect 2148 56545 2176 58511
rect 579526 57624 579582 57633
rect 579632 57610 579660 59599
rect 579582 57582 579660 57610
rect 579526 57559 579582 57568
rect 2134 56536 2190 56545
rect 2134 56471 2190 56480
rect 579986 46336 580042 46345
rect 579986 46271 580042 46280
rect 3422 45520 3478 45529
rect 3422 45455 3478 45464
rect 3436 43333 3464 45455
rect 580000 45014 580028 46271
rect 578332 45008 578384 45014
rect 578332 44950 578384 44956
rect 579988 45008 580040 45014
rect 579988 44950 580040 44956
rect 578344 44305 578372 44950
rect 578330 44296 578386 44305
rect 578330 44231 578386 44240
rect 3422 43324 3478 43333
rect 3422 43259 3478 43268
rect 579618 33144 579674 33153
rect 579618 33079 579674 33088
rect 2134 32464 2190 32473
rect 2134 32399 2190 32408
rect 2148 30297 2176 32399
rect 579526 30968 579582 30977
rect 579632 30954 579660 33079
rect 579582 30926 579660 30954
rect 579526 30903 579582 30912
rect 2134 30288 2190 30297
rect 2134 30223 2190 30232
rect 579618 19816 579674 19825
rect 579618 19751 579674 19760
rect 2042 19408 2098 19417
rect 2042 19343 2098 19352
rect 2056 17241 2084 19343
rect 579526 17640 579582 17649
rect 579632 17626 579660 19751
rect 579582 17598 579660 17626
rect 579526 17575 579582 17584
rect 2042 17232 2098 17241
rect 2042 17167 2098 17176
rect 579618 6624 579674 6633
rect 579618 6559 579674 6568
rect 2778 6488 2834 6497
rect 2778 6423 2834 6432
rect 2792 4185 2820 6423
rect 579632 5574 579660 6559
rect 576860 5568 576912 5574
rect 576860 5510 576912 5516
rect 579620 5568 579672 5574
rect 579620 5510 579672 5516
rect 2778 4176 2834 4185
rect 2778 4111 2834 4120
rect 576766 4176 576822 4185
rect 576872 4162 576900 5510
rect 576822 4134 576900 4162
rect 576766 4111 576822 4120
rect 1676 3868 1728 3874
rect 1676 3810 1728 3816
rect 572 3800 624 3806
rect 572 3742 624 3748
rect 584 480 612 3742
rect 1688 480 1716 3810
rect 4124 3806 4152 4012
rect 5228 3874 5256 4012
rect 5216 3868 5268 3874
rect 5216 3810 5268 3816
rect 4112 3800 4164 3806
rect 6424 3754 6452 4012
rect 7528 3754 7556 4012
rect 4112 3742 4164 3748
rect 6380 3726 6452 3754
rect 7484 3726 7556 3754
rect 7656 3800 7708 3806
rect 8724 3754 8752 4012
rect 9920 3754 9948 4012
rect 11024 3806 11052 4012
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 7656 3742 7708 3748
rect 4068 2848 4120 2854
rect 4068 2790 4120 2796
rect 3240 1352 3292 1358
rect 3240 1294 3292 1300
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 354 2954 480
rect 3252 354 3280 1294
rect 4080 480 4108 2790
rect 6380 1358 6408 3726
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6368 1352 6420 1358
rect 6368 1294 6420 1300
rect 5632 1148 5684 1154
rect 5632 1090 5684 1096
rect 2842 326 3280 354
rect 2842 -960 2954 326
rect 4038 -960 4150 480
rect 5234 354 5346 480
rect 5644 354 5672 1090
rect 6472 480 6500 2994
rect 7484 2854 7512 3726
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 7668 480 7696 3742
rect 8680 3726 8752 3754
rect 9876 3726 9948 3754
rect 11012 3800 11064 3806
rect 11012 3742 11064 3748
rect 8680 1154 8708 3726
rect 9876 3058 9904 3726
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 8668 1148 8720 1154
rect 8668 1090 8720 1096
rect 8760 944 8812 950
rect 8760 886 8812 892
rect 8772 480 8800 886
rect 9968 480 9996 2790
rect 11164 480 11192 3878
rect 12220 3754 12248 4012
rect 12176 3726 12248 3754
rect 12348 3800 12400 3806
rect 13324 3754 13352 4012
rect 14520 3942 14548 4012
rect 14508 3936 14560 3942
rect 14508 3878 14560 3884
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 13544 3868 13596 3874
rect 13544 3810 13596 3816
rect 12348 3742 12400 3748
rect 12176 950 12204 3726
rect 12164 944 12216 950
rect 12164 886 12216 892
rect 12360 480 12388 3742
rect 13280 3726 13352 3754
rect 13280 2854 13308 3726
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 13556 480 13584 3810
rect 14752 480 14780 3878
rect 15716 3806 15744 4012
rect 16820 3874 16848 4012
rect 18016 3942 18044 4012
rect 18004 3936 18056 3942
rect 18004 3878 18056 3884
rect 16808 3868 16860 3874
rect 16808 3810 16860 3816
rect 19120 3806 19148 4012
rect 19432 3868 19484 3874
rect 19432 3810 19484 3816
rect 15704 3800 15756 3806
rect 15704 3742 15756 3748
rect 15936 3800 15988 3806
rect 15936 3742 15988 3748
rect 19108 3800 19160 3806
rect 19108 3742 19160 3748
rect 15948 480 15976 3742
rect 18236 2916 18288 2922
rect 18236 2858 18288 2864
rect 17040 2848 17092 2854
rect 17040 2790 17092 2796
rect 17052 480 17080 2790
rect 18248 480 18276 2858
rect 19444 480 19472 3810
rect 20316 3754 20344 4012
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 20272 3726 20344 3754
rect 20272 2854 20300 3726
rect 20260 2848 20312 2854
rect 20260 2790 20312 2796
rect 20640 480 20668 3878
rect 21512 3754 21540 4012
rect 22616 3874 22644 4012
rect 23812 3942 23840 4012
rect 23800 3936 23852 3942
rect 23800 3878 23852 3884
rect 24216 3936 24268 3942
rect 24216 3878 24268 3884
rect 22604 3868 22656 3874
rect 22604 3810 22656 3816
rect 23020 3868 23072 3874
rect 23020 3810 23072 3816
rect 21468 3726 21540 3754
rect 21824 3800 21876 3806
rect 21824 3742 21876 3748
rect 21468 2922 21496 3726
rect 21456 2916 21508 2922
rect 21456 2858 21508 2864
rect 21836 480 21864 3742
rect 23032 480 23060 3810
rect 24228 480 24256 3878
rect 24916 3806 24944 4012
rect 26112 3874 26140 4012
rect 27308 3942 27336 4012
rect 27296 3936 27348 3942
rect 27296 3878 27348 3884
rect 27712 3936 27764 3942
rect 27712 3878 27764 3884
rect 26100 3868 26152 3874
rect 26100 3810 26152 3816
rect 26516 3868 26568 3874
rect 26516 3810 26568 3816
rect 24904 3800 24956 3806
rect 24904 3742 24956 3748
rect 25320 3800 25372 3806
rect 25320 3742 25372 3748
rect 25332 480 25360 3742
rect 26528 480 26556 3810
rect 27724 480 27752 3878
rect 28412 3806 28440 4012
rect 29608 3874 29636 4012
rect 30712 3942 30740 4012
rect 30700 3936 30752 3942
rect 30700 3878 30752 3884
rect 29596 3868 29648 3874
rect 29596 3810 29648 3816
rect 30104 3868 30156 3874
rect 30104 3810 30156 3816
rect 28400 3800 28452 3806
rect 28400 3742 28452 3748
rect 28908 2848 28960 2854
rect 28908 2790 28960 2796
rect 28920 480 28948 2790
rect 30116 480 30144 3810
rect 31300 3800 31352 3806
rect 31908 3754 31936 4012
rect 32404 3936 32456 3942
rect 32404 3878 32456 3884
rect 31300 3742 31352 3748
rect 31312 480 31340 3742
rect 31864 3726 31936 3754
rect 31864 2854 31892 3726
rect 31852 2848 31904 2854
rect 31852 2790 31904 2796
rect 32416 480 32444 3878
rect 33104 3874 33132 4012
rect 33092 3868 33144 3874
rect 33092 3810 33144 3816
rect 33600 3868 33652 3874
rect 33600 3810 33652 3816
rect 33612 480 33640 3810
rect 34208 3806 34236 4012
rect 35404 3942 35432 4012
rect 35392 3936 35444 3942
rect 35392 3878 35444 3884
rect 36600 3874 36628 4012
rect 36588 3868 36640 3874
rect 36588 3810 36640 3816
rect 37188 3868 37240 3874
rect 37188 3810 37240 3816
rect 34196 3800 34248 3806
rect 34196 3742 34248 3748
rect 34796 3800 34848 3806
rect 34796 3742 34848 3748
rect 34808 480 34836 3742
rect 35992 2848 36044 2854
rect 35992 2790 36044 2796
rect 36004 480 36032 2790
rect 37200 480 37228 3810
rect 37704 3806 37732 4012
rect 38384 3936 38436 3942
rect 38384 3878 38436 3884
rect 37692 3800 37744 3806
rect 37692 3742 37744 3748
rect 38396 480 38424 3878
rect 38900 3754 38928 4012
rect 40004 3874 40032 4012
rect 41200 3942 41228 4012
rect 41188 3936 41240 3942
rect 41188 3878 41240 3884
rect 39992 3868 40044 3874
rect 39992 3810 40044 3816
rect 41880 3868 41932 3874
rect 41880 3810 41932 3816
rect 38856 3726 38928 3754
rect 40684 3800 40736 3806
rect 40684 3742 40736 3748
rect 38856 2854 38884 3726
rect 38844 2848 38896 2854
rect 38844 2790 38896 2796
rect 39580 2848 39632 2854
rect 39580 2790 39632 2796
rect 39592 480 39620 2790
rect 40696 480 40724 3742
rect 41892 480 41920 3810
rect 42396 3754 42424 4012
rect 43076 3936 43128 3942
rect 43076 3878 43128 3884
rect 42352 3726 42424 3754
rect 42352 2854 42380 3726
rect 42340 2848 42392 2854
rect 42340 2790 42392 2796
rect 43088 480 43116 3878
rect 43500 3806 43528 4012
rect 44696 3874 44724 4012
rect 45800 3942 45828 4012
rect 45788 3936 45840 3942
rect 45788 3878 45840 3884
rect 46664 3936 46716 3942
rect 46664 3878 46716 3884
rect 44684 3868 44736 3874
rect 44684 3810 44736 3816
rect 45468 3868 45520 3874
rect 45468 3810 45520 3816
rect 43488 3800 43540 3806
rect 43488 3742 43540 3748
rect 44272 3800 44324 3806
rect 44272 3742 44324 3748
rect 44284 480 44312 3742
rect 45480 480 45508 3810
rect 46676 480 46704 3878
rect 46996 3806 47024 4012
rect 48192 3874 48220 4012
rect 49296 3942 49324 4012
rect 49284 3936 49336 3942
rect 49284 3878 49336 3884
rect 50160 3936 50212 3942
rect 50160 3878 50212 3884
rect 48180 3868 48232 3874
rect 48180 3810 48232 3816
rect 48964 3868 49016 3874
rect 48964 3810 49016 3816
rect 46984 3800 47036 3806
rect 46984 3742 47036 3748
rect 47860 3800 47912 3806
rect 47860 3742 47912 3748
rect 47872 480 47900 3742
rect 48976 480 49004 3810
rect 50172 480 50200 3878
rect 50492 3806 50520 4012
rect 51596 3874 51624 4012
rect 52792 3942 52820 4012
rect 52780 3936 52832 3942
rect 52780 3878 52832 3884
rect 51584 3868 51636 3874
rect 51584 3810 51636 3816
rect 53748 3868 53800 3874
rect 53748 3810 53800 3816
rect 50480 3800 50532 3806
rect 50480 3742 50532 3748
rect 51356 3800 51408 3806
rect 51356 3742 51408 3748
rect 51368 480 51396 3742
rect 52552 740 52604 746
rect 52552 682 52604 688
rect 52564 480 52592 682
rect 53760 480 53788 3810
rect 53988 3806 54016 4012
rect 53976 3800 54028 3806
rect 53976 3742 54028 3748
rect 54944 3800 54996 3806
rect 55092 3754 55120 4012
rect 56048 3936 56100 3942
rect 56048 3878 56100 3884
rect 54944 3742 54996 3748
rect 54956 480 54984 3742
rect 55048 3726 55120 3754
rect 55048 746 55076 3726
rect 55036 740 55088 746
rect 55036 682 55088 688
rect 56060 480 56088 3878
rect 56288 3874 56316 4012
rect 56276 3868 56328 3874
rect 56276 3810 56328 3816
rect 57244 3868 57296 3874
rect 57244 3810 57296 3816
rect 57256 480 57284 3810
rect 57392 3806 57420 4012
rect 58588 3942 58616 4012
rect 58576 3936 58628 3942
rect 58576 3878 58628 3884
rect 59784 3874 59812 4012
rect 59772 3868 59824 3874
rect 59772 3810 59824 3816
rect 60888 3806 60916 4012
rect 62084 3890 62112 4012
rect 61948 3862 62112 3890
rect 57380 3800 57432 3806
rect 57380 3742 57432 3748
rect 58440 3800 58492 3806
rect 58440 3742 58492 3748
rect 60876 3800 60928 3806
rect 60876 3742 60928 3748
rect 58452 480 58480 3742
rect 60832 1352 60884 1358
rect 60832 1294 60884 1300
rect 59636 740 59688 746
rect 59636 682 59688 688
rect 59648 480 59676 682
rect 60844 480 60872 1294
rect 61948 746 61976 3862
rect 63280 3754 63308 4012
rect 64384 3890 64412 4012
rect 64384 3862 64460 3890
rect 64328 3800 64380 3806
rect 63280 3726 63356 3754
rect 64328 3742 64380 3748
rect 63224 3052 63276 3058
rect 63224 2994 63276 3000
rect 62028 2848 62080 2854
rect 62028 2790 62080 2796
rect 61936 740 61988 746
rect 61936 682 61988 688
rect 62040 480 62068 2790
rect 63236 480 63264 2994
rect 63328 1358 63356 3726
rect 63316 1352 63368 1358
rect 63316 1294 63368 1300
rect 64340 480 64368 3742
rect 64432 2854 64460 3862
rect 65580 3754 65608 4012
rect 66684 3806 66712 4012
rect 65536 3726 65608 3754
rect 66672 3800 66724 3806
rect 66672 3742 66724 3748
rect 67088 3800 67140 3806
rect 67880 3754 67908 4012
rect 69076 3806 69104 4012
rect 67088 3742 67140 3748
rect 65536 3058 65564 3726
rect 65524 3052 65576 3058
rect 65524 2994 65576 3000
rect 64420 2848 64472 2854
rect 64420 2790 64472 2796
rect 65524 2848 65576 2854
rect 65524 2790 65576 2796
rect 65536 480 65564 2790
rect 5234 326 5672 354
rect 5234 -960 5346 326
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 354 66802 480
rect 67100 354 67128 3742
rect 67836 3726 67908 3754
rect 69064 3800 69116 3806
rect 70180 3754 70208 4012
rect 69064 3742 69116 3748
rect 70136 3726 70208 3754
rect 70308 3800 70360 3806
rect 71376 3754 71404 4012
rect 71504 3868 71556 3874
rect 71504 3810 71556 3816
rect 70308 3742 70360 3748
rect 67836 2854 67864 3726
rect 67824 2848 67876 2854
rect 67824 2790 67876 2796
rect 70136 1358 70164 3726
rect 67916 1352 67968 1358
rect 67916 1294 67968 1300
rect 70124 1352 70176 1358
rect 70124 1294 70176 1300
rect 67928 480 67956 1294
rect 69112 604 69164 610
rect 69112 546 69164 552
rect 69124 480 69152 546
rect 70320 480 70348 3742
rect 71332 3726 71404 3754
rect 71332 610 71360 3726
rect 71320 604 71372 610
rect 71320 546 71372 552
rect 71516 480 71544 3810
rect 72480 3806 72508 4012
rect 72608 3936 72660 3942
rect 72608 3878 72660 3884
rect 72468 3800 72520 3806
rect 72468 3742 72520 3748
rect 72620 480 72648 3878
rect 73676 3874 73704 4012
rect 74872 3942 74900 4012
rect 74860 3936 74912 3942
rect 74860 3878 74912 3884
rect 73664 3868 73716 3874
rect 73664 3810 73716 3816
rect 75976 3806 76004 4012
rect 73804 3800 73856 3806
rect 73804 3742 73856 3748
rect 75964 3800 76016 3806
rect 77172 3754 77200 4012
rect 78276 3754 78304 4012
rect 78588 3868 78640 3874
rect 78588 3810 78640 3816
rect 75964 3742 76016 3748
rect 73816 480 73844 3742
rect 77128 3726 77200 3754
rect 78232 3726 78304 3754
rect 76196 1352 76248 1358
rect 76196 1294 76248 1300
rect 75000 1284 75052 1290
rect 75000 1226 75052 1232
rect 75012 480 75040 1226
rect 76208 480 76236 1294
rect 77128 1290 77156 3726
rect 78232 1358 78260 3726
rect 78220 1352 78272 1358
rect 78220 1294 78272 1300
rect 77116 1284 77168 1290
rect 77116 1226 77168 1232
rect 77392 1284 77444 1290
rect 77392 1226 77444 1232
rect 77404 480 77432 1226
rect 78600 480 78628 3810
rect 79472 3754 79500 4012
rect 80668 3874 80696 4012
rect 80656 3868 80708 3874
rect 80656 3810 80708 3816
rect 80888 3868 80940 3874
rect 80888 3810 80940 3816
rect 79428 3726 79500 3754
rect 79692 3800 79744 3806
rect 79692 3742 79744 3748
rect 79428 1290 79456 3726
rect 79416 1284 79468 1290
rect 79416 1226 79468 1232
rect 79704 480 79732 3742
rect 80900 480 80928 3810
rect 81772 3806 81800 4012
rect 82968 3874 82996 4012
rect 82956 3868 83008 3874
rect 82956 3810 83008 3816
rect 81760 3800 81812 3806
rect 84072 3754 84100 4012
rect 85268 3754 85296 4012
rect 86464 3754 86492 4012
rect 81760 3742 81812 3748
rect 84028 3726 84100 3754
rect 85224 3726 85296 3754
rect 86420 3726 86492 3754
rect 86868 3800 86920 3806
rect 87568 3754 87596 4012
rect 87972 3868 88024 3874
rect 87972 3810 88024 3816
rect 86868 3742 86920 3748
rect 83280 1352 83332 1358
rect 83280 1294 83332 1300
rect 82084 1284 82136 1290
rect 82084 1226 82136 1232
rect 82096 480 82124 1226
rect 83292 480 83320 1294
rect 84028 1290 84056 3726
rect 85224 1358 85252 3726
rect 85212 1352 85264 1358
rect 85212 1294 85264 1300
rect 85672 1352 85724 1358
rect 85672 1294 85724 1300
rect 84016 1284 84068 1290
rect 84016 1226 84068 1232
rect 84476 1284 84528 1290
rect 84476 1226 84528 1232
rect 84488 480 84516 1226
rect 85684 480 85712 1294
rect 86420 1290 86448 3726
rect 86408 1284 86460 1290
rect 86408 1226 86460 1232
rect 86880 480 86908 3742
rect 87524 3726 87596 3754
rect 87524 1358 87552 3726
rect 87512 1352 87564 1358
rect 87512 1294 87564 1300
rect 87984 480 88012 3810
rect 88764 3806 88792 4012
rect 89960 3874 89988 4012
rect 89948 3868 90000 3874
rect 89948 3810 90000 3816
rect 88752 3800 88804 3806
rect 91064 3754 91092 4012
rect 92260 3754 92288 4012
rect 93364 3754 93392 4012
rect 94560 3754 94588 4012
rect 88752 3742 88804 3748
rect 91020 3726 91092 3754
rect 92216 3726 92288 3754
rect 93320 3726 93392 3754
rect 94516 3726 94588 3754
rect 95148 3800 95200 3806
rect 95756 3754 95784 4012
rect 96252 3868 96304 3874
rect 96252 3810 96304 3816
rect 95148 3742 95200 3748
rect 91020 1358 91048 3726
rect 89168 1352 89220 1358
rect 89168 1294 89220 1300
rect 91008 1352 91060 1358
rect 91008 1294 91060 1300
rect 91560 1352 91612 1358
rect 91560 1294 91612 1300
rect 89180 480 89208 1294
rect 90364 1284 90416 1290
rect 90364 1226 90416 1232
rect 90376 480 90404 1226
rect 91572 480 91600 1294
rect 92216 1290 92244 3726
rect 93320 1358 93348 3726
rect 93308 1352 93360 1358
rect 93308 1294 93360 1300
rect 93952 1352 94004 1358
rect 93952 1294 94004 1300
rect 92204 1284 92256 1290
rect 92204 1226 92256 1232
rect 92756 1284 92808 1290
rect 92756 1226 92808 1232
rect 92768 480 92796 1226
rect 93964 480 93992 1294
rect 94516 1290 94544 3726
rect 94504 1284 94556 1290
rect 94504 1226 94556 1232
rect 95160 480 95188 3742
rect 95712 3726 95784 3754
rect 95712 1358 95740 3726
rect 95700 1352 95752 1358
rect 95700 1294 95752 1300
rect 96264 480 96292 3810
rect 96860 3806 96888 4012
rect 98056 3874 98084 4012
rect 98044 3868 98096 3874
rect 98044 3810 98096 3816
rect 96848 3800 96900 3806
rect 99160 3754 99188 4012
rect 100356 3754 100384 4012
rect 101552 3754 101580 4012
rect 102656 3754 102684 4012
rect 96848 3742 96900 3748
rect 99116 3726 99188 3754
rect 100312 3726 100384 3754
rect 101508 3726 101580 3754
rect 102612 3726 102684 3754
rect 103336 3800 103388 3806
rect 103852 3754 103880 4012
rect 104956 3806 104984 4012
rect 103336 3742 103388 3748
rect 99116 1358 99144 3726
rect 97448 1352 97500 1358
rect 97448 1294 97500 1300
rect 99104 1352 99156 1358
rect 99104 1294 99156 1300
rect 97460 480 97488 1294
rect 100312 1290 100340 3726
rect 101036 1352 101088 1358
rect 101036 1294 101088 1300
rect 98644 1284 98696 1290
rect 98644 1226 98696 1232
rect 100300 1284 100352 1290
rect 100300 1226 100352 1232
rect 98656 480 98684 1226
rect 99840 1216 99892 1222
rect 99840 1158 99892 1164
rect 99852 480 99880 1158
rect 101048 480 101076 1294
rect 101508 1222 101536 3726
rect 102612 1358 102640 3726
rect 102600 1352 102652 1358
rect 102600 1294 102652 1300
rect 102232 1284 102284 1290
rect 102232 1226 102284 1232
rect 101496 1216 101548 1222
rect 101496 1158 101548 1164
rect 102244 480 102272 1226
rect 103348 480 103376 3742
rect 103808 3726 103880 3754
rect 104944 3800 104996 3806
rect 106152 3754 106180 4012
rect 107348 3754 107376 4012
rect 108452 3754 108480 4012
rect 109648 3754 109676 4012
rect 110752 3754 110780 4012
rect 111948 3754 111976 4012
rect 113144 3754 113172 4012
rect 114248 3754 114276 4012
rect 115444 3754 115472 4012
rect 116640 3754 116668 4012
rect 117744 3754 117772 4012
rect 118940 3754 118968 4012
rect 120044 3754 120072 4012
rect 121240 3754 121268 4012
rect 122436 3754 122464 4012
rect 123540 3754 123568 4012
rect 104944 3742 104996 3748
rect 106108 3726 106180 3754
rect 107304 3726 107376 3754
rect 108408 3726 108480 3754
rect 109604 3726 109676 3754
rect 110708 3726 110780 3754
rect 111904 3726 111976 3754
rect 113100 3726 113172 3754
rect 114204 3726 114276 3754
rect 115400 3726 115472 3754
rect 116596 3726 116668 3754
rect 117700 3726 117772 3754
rect 118896 3726 118968 3754
rect 119264 3726 120072 3754
rect 121196 3726 121268 3754
rect 122392 3726 122464 3754
rect 123496 3726 123568 3754
rect 124736 3754 124764 4012
rect 125840 3754 125868 4012
rect 127036 3754 127064 4012
rect 128232 3754 128260 4012
rect 129336 3754 129364 4012
rect 130532 3754 130560 4012
rect 131636 3754 131664 4012
rect 132832 3754 132860 4012
rect 134028 3754 134056 4012
rect 135132 3754 135160 4012
rect 136328 3754 136356 4012
rect 137432 3754 137460 4012
rect 138628 3754 138656 4012
rect 139824 3754 139852 4012
rect 140928 3754 140956 4012
rect 142124 3754 142152 4012
rect 143320 3754 143348 4012
rect 144424 3754 144452 4012
rect 145620 3754 145648 4012
rect 146724 3754 146752 4012
rect 147920 3754 147948 4012
rect 149116 3754 149144 4012
rect 150220 3754 150248 4012
rect 151416 3754 151444 4012
rect 152520 3754 152548 4012
rect 153716 3754 153744 4012
rect 154912 3754 154940 4012
rect 156016 3754 156044 4012
rect 157212 3754 157240 4012
rect 158316 3754 158344 4012
rect 159512 3754 159540 4012
rect 160708 3754 160736 4012
rect 161812 3754 161840 4012
rect 163008 3754 163036 4012
rect 164112 3754 164140 4012
rect 165308 3754 165336 4012
rect 166504 3754 166532 4012
rect 167608 3754 167636 4012
rect 168804 3754 168832 4012
rect 170000 3754 170028 4012
rect 171104 3754 171132 4012
rect 172300 3754 172328 4012
rect 173404 3754 173432 4012
rect 174600 3754 174628 4012
rect 175796 3754 175824 4012
rect 176900 3754 176928 4012
rect 178096 3754 178124 4012
rect 179200 3754 179228 4012
rect 124736 3726 124812 3754
rect 103808 1290 103836 3726
rect 106108 1358 106136 3726
rect 104532 1352 104584 1358
rect 104532 1294 104584 1300
rect 106096 1352 106148 1358
rect 106096 1294 106148 1300
rect 106924 1352 106976 1358
rect 106924 1294 106976 1300
rect 103796 1284 103848 1290
rect 103796 1226 103848 1232
rect 104544 480 104572 1294
rect 105728 740 105780 746
rect 105728 682 105780 688
rect 105740 480 105768 682
rect 106936 480 106964 1294
rect 107304 746 107332 3726
rect 108408 1358 108436 3726
rect 108396 1352 108448 1358
rect 108396 1294 108448 1300
rect 109316 1352 109368 1358
rect 109316 1294 109368 1300
rect 108120 1284 108172 1290
rect 108120 1226 108172 1232
rect 107292 740 107344 746
rect 107292 682 107344 688
rect 108132 480 108160 1226
rect 109328 480 109356 1294
rect 109604 1290 109632 3726
rect 110708 1358 110736 3726
rect 110696 1352 110748 1358
rect 110696 1294 110748 1300
rect 111904 1290 111932 3726
rect 112812 1352 112864 1358
rect 112812 1294 112864 1300
rect 109592 1284 109644 1290
rect 109592 1226 109644 1232
rect 110512 1284 110564 1290
rect 110512 1226 110564 1232
rect 111892 1284 111944 1290
rect 111892 1226 111944 1232
rect 110524 480 110552 1226
rect 111616 1148 111668 1154
rect 111616 1090 111668 1096
rect 111628 480 111656 1090
rect 112824 480 112852 1294
rect 113100 1154 113128 3726
rect 114204 1358 114232 3726
rect 114192 1352 114244 1358
rect 114192 1294 114244 1300
rect 115204 1284 115256 1290
rect 115204 1226 115256 1232
rect 114008 1216 114060 1222
rect 114008 1158 114060 1164
rect 113088 1148 113140 1154
rect 113088 1090 113140 1096
rect 114020 480 114048 1158
rect 115216 480 115244 1226
rect 115400 1222 115428 3726
rect 116400 1352 116452 1358
rect 116400 1294 116452 1300
rect 115388 1216 115440 1222
rect 115388 1158 115440 1164
rect 116412 480 116440 1294
rect 116596 1290 116624 3726
rect 117700 1358 117728 3726
rect 117688 1352 117740 1358
rect 117688 1294 117740 1300
rect 118896 1290 118924 3726
rect 116584 1284 116636 1290
rect 116584 1226 116636 1232
rect 117596 1284 117648 1290
rect 117596 1226 117648 1232
rect 118884 1284 118936 1290
rect 118884 1226 118936 1232
rect 117608 480 117636 1226
rect 66690 326 67128 354
rect 66690 -960 66802 326
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 354 118874 480
rect 119264 354 119292 3726
rect 121196 1358 121224 3726
rect 119896 1352 119948 1358
rect 119896 1294 119948 1300
rect 121184 1352 121236 1358
rect 121184 1294 121236 1300
rect 119908 480 119936 1294
rect 122288 1284 122340 1290
rect 122288 1226 122340 1232
rect 121092 944 121144 950
rect 121092 886 121144 892
rect 121104 480 121132 886
rect 122300 480 122328 1226
rect 122392 950 122420 3726
rect 123496 1290 123524 3726
rect 123484 1284 123536 1290
rect 123484 1226 123536 1232
rect 124680 1284 124732 1290
rect 124680 1226 124732 1232
rect 123484 1148 123536 1154
rect 123484 1090 123536 1096
rect 122380 944 122432 950
rect 122380 886 122432 892
rect 123496 480 123524 1090
rect 124692 480 124720 1226
rect 124784 1154 124812 3726
rect 125796 3726 125868 3754
rect 126992 3726 127064 3754
rect 127176 3726 128260 3754
rect 129292 3726 129364 3754
rect 130488 3726 130560 3754
rect 131592 3726 131664 3754
rect 132788 3726 132860 3754
rect 133984 3726 134056 3754
rect 134168 3726 135160 3754
rect 135272 3726 136356 3754
rect 137388 3726 137460 3754
rect 138584 3726 138656 3754
rect 139780 3726 139852 3754
rect 140884 3726 140956 3754
rect 141712 3726 142152 3754
rect 142448 3726 143348 3754
rect 143552 3726 144452 3754
rect 145576 3726 145648 3754
rect 146680 3726 146752 3754
rect 147600 3726 147948 3754
rect 149072 3726 149144 3754
rect 149992 3726 150248 3754
rect 151096 3726 151444 3754
rect 151832 3726 152548 3754
rect 153488 3726 153744 3754
rect 154868 3726 154940 3754
rect 155880 3726 156044 3754
rect 156616 3726 157240 3754
rect 158272 3726 158344 3754
rect 159376 3726 159540 3754
rect 160112 3726 160736 3754
rect 161584 3726 161840 3754
rect 162964 3726 163036 3754
rect 164068 3726 164140 3754
rect 164896 3726 165336 3754
rect 166460 3726 166532 3754
rect 167564 3726 167636 3754
rect 168392 3726 168832 3754
rect 169956 3726 170028 3754
rect 170784 3726 171132 3754
rect 172256 3726 172328 3754
rect 173176 3726 173432 3754
rect 174280 3726 174628 3754
rect 175752 3726 175824 3754
rect 176672 3726 176928 3754
rect 178052 3726 178124 3754
rect 179064 3726 179228 3754
rect 180396 3754 180424 4012
rect 181592 3754 181620 4012
rect 182696 3754 182724 4012
rect 180396 3726 180472 3754
rect 125796 1290 125824 3726
rect 126992 1358 127020 3726
rect 125876 1352 125928 1358
rect 125876 1294 125928 1300
rect 126980 1352 127032 1358
rect 126980 1294 127032 1300
rect 125784 1284 125836 1290
rect 125784 1226 125836 1232
rect 124772 1148 124824 1154
rect 124772 1090 124824 1096
rect 125888 480 125916 1294
rect 127176 1170 127204 3726
rect 129292 1290 129320 3726
rect 130488 1358 130516 3726
rect 131592 1358 131620 3726
rect 132788 1358 132816 3726
rect 133984 1358 134012 3726
rect 129372 1352 129424 1358
rect 129372 1294 129424 1300
rect 130476 1352 130528 1358
rect 130476 1294 130528 1300
rect 130568 1352 130620 1358
rect 130568 1294 130620 1300
rect 131580 1352 131632 1358
rect 131580 1294 131632 1300
rect 131764 1352 131816 1358
rect 131764 1294 131816 1300
rect 132776 1352 132828 1358
rect 132776 1294 132828 1300
rect 132960 1352 133012 1358
rect 132960 1294 133012 1300
rect 133972 1352 134024 1358
rect 133972 1294 134024 1300
rect 128176 1284 128228 1290
rect 128176 1226 128228 1232
rect 129280 1284 129332 1290
rect 129280 1226 129332 1232
rect 126992 1142 127204 1170
rect 126992 480 127020 1142
rect 128188 480 128216 1226
rect 129384 480 129412 1294
rect 130580 480 130608 1294
rect 131776 480 131804 1294
rect 132972 480 133000 1294
rect 134168 480 134196 3726
rect 135272 480 135300 3726
rect 137388 1290 137416 3726
rect 138584 1358 138612 3726
rect 137652 1352 137704 1358
rect 137652 1294 137704 1300
rect 138572 1352 138624 1358
rect 138572 1294 138624 1300
rect 136456 1284 136508 1290
rect 136456 1226 136508 1232
rect 137376 1284 137428 1290
rect 137376 1226 137428 1232
rect 136468 480 136496 1226
rect 137664 480 137692 1294
rect 139780 1290 139808 3726
rect 140884 1290 140912 3726
rect 138848 1284 138900 1290
rect 138848 1226 138900 1232
rect 139768 1284 139820 1290
rect 139768 1226 139820 1232
rect 140044 1284 140096 1290
rect 140044 1226 140096 1232
rect 140872 1284 140924 1290
rect 140872 1226 140924 1232
rect 138860 480 138888 1226
rect 140056 480 140084 1226
rect 118762 326 119292 354
rect 118762 -960 118874 326
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 354 141322 480
rect 141712 354 141740 3726
rect 142448 480 142476 3726
rect 143552 480 143580 3726
rect 145576 1358 145604 3726
rect 146680 1358 146708 3726
rect 144736 1352 144788 1358
rect 144736 1294 144788 1300
rect 145564 1352 145616 1358
rect 145564 1294 145616 1300
rect 145932 1352 145984 1358
rect 145932 1294 145984 1300
rect 146668 1352 146720 1358
rect 146668 1294 146720 1300
rect 144748 480 144776 1294
rect 145944 480 145972 1294
rect 141210 326 141740 354
rect 141210 -960 141322 326
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 354 147210 480
rect 147600 354 147628 3726
rect 149072 1358 149100 3726
rect 148324 1352 148376 1358
rect 148324 1294 148376 1300
rect 149060 1352 149112 1358
rect 149060 1294 149112 1300
rect 148336 480 148364 1294
rect 147098 326 147628 354
rect 147098 -960 147210 326
rect 148294 -960 148406 480
rect 149490 354 149602 480
rect 149992 354 150020 3726
rect 149490 326 150020 354
rect 150594 354 150706 480
rect 151096 354 151124 3726
rect 151832 480 151860 3726
rect 150594 326 151124 354
rect 149490 -960 149602 326
rect 150594 -960 150706 326
rect 151790 -960 151902 480
rect 152986 354 153098 480
rect 153488 354 153516 3726
rect 154868 1358 154896 3726
rect 154212 1352 154264 1358
rect 154212 1294 154264 1300
rect 154856 1352 154908 1358
rect 154856 1294 154908 1300
rect 154224 480 154252 1294
rect 152986 326 153516 354
rect 152986 -960 153098 326
rect 154182 -960 154294 480
rect 155378 354 155490 480
rect 155880 354 155908 3726
rect 156616 480 156644 3726
rect 155378 326 155908 354
rect 155378 -960 155490 326
rect 156574 -960 156686 480
rect 157770 354 157882 480
rect 158272 354 158300 3726
rect 157770 326 158300 354
rect 158874 354 158986 480
rect 159376 354 159404 3726
rect 160112 480 160140 3726
rect 158874 326 159404 354
rect 157770 -960 157882 326
rect 158874 -960 158986 326
rect 160070 -960 160182 480
rect 161266 354 161378 480
rect 161584 354 161612 3726
rect 162964 1358 162992 3726
rect 162492 1352 162544 1358
rect 162492 1294 162544 1300
rect 162952 1352 163004 1358
rect 162952 1294 163004 1300
rect 162504 480 162532 1294
rect 161266 326 161612 354
rect 161266 -960 161378 326
rect 162462 -960 162574 480
rect 163658 354 163770 480
rect 164068 354 164096 3726
rect 164896 480 164924 3726
rect 163658 326 164096 354
rect 163658 -960 163770 326
rect 164854 -960 164966 480
rect 166050 354 166162 480
rect 166460 354 166488 3726
rect 166050 326 166488 354
rect 167154 354 167266 480
rect 167564 354 167592 3726
rect 168392 480 168420 3726
rect 167154 326 167592 354
rect 166050 -960 166162 326
rect 167154 -960 167266 326
rect 168350 -960 168462 480
rect 169546 354 169658 480
rect 169956 354 169984 3726
rect 170784 480 170812 3726
rect 169546 326 169984 354
rect 169546 -960 169658 326
rect 170742 -960 170854 480
rect 171938 354 172050 480
rect 172256 354 172284 3726
rect 173176 480 173204 3726
rect 174280 480 174308 3726
rect 171938 326 172284 354
rect 171938 -960 172050 326
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 354 175546 480
rect 175752 354 175780 3726
rect 176672 480 176700 3726
rect 175434 326 175780 354
rect 175434 -960 175546 326
rect 176630 -960 176742 480
rect 177826 354 177938 480
rect 178052 354 178080 3726
rect 179064 480 179092 3726
rect 177826 326 178080 354
rect 177826 -960 177938 326
rect 179022 -960 179134 480
rect 180218 218 180330 480
rect 180444 218 180472 3726
rect 181456 3726 181620 3754
rect 182560 3726 182724 3754
rect 183892 3754 183920 4012
rect 184996 3754 185024 4012
rect 186192 3754 186220 4012
rect 187388 3754 187416 4012
rect 183892 3726 183968 3754
rect 181456 480 181484 3726
rect 182560 480 182588 3726
rect 180218 190 180472 218
rect 180218 -960 180330 190
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 218 183826 480
rect 183940 218 183968 3726
rect 184952 3726 185024 3754
rect 186148 3726 186220 3754
rect 187344 3726 187416 3754
rect 188492 3754 188520 4012
rect 189688 3754 189716 4012
rect 190792 3754 190820 4012
rect 191988 3754 192016 4012
rect 193184 3754 193212 4012
rect 194288 3754 194316 4012
rect 195484 3754 195512 4012
rect 188492 3726 188568 3754
rect 189688 3726 189764 3754
rect 190792 3726 190868 3754
rect 191988 3726 192064 3754
rect 193184 3726 193260 3754
rect 194288 3726 194456 3754
rect 184952 480 184980 3726
rect 186148 480 186176 3726
rect 187344 480 187372 3726
rect 188540 480 188568 3726
rect 189736 480 189764 3726
rect 190840 480 190868 3726
rect 192036 480 192064 3726
rect 193232 480 193260 3726
rect 194428 480 194456 3726
rect 195440 3726 195512 3754
rect 196680 3754 196708 4012
rect 197784 3754 197812 4012
rect 198980 3754 199008 4012
rect 196680 3726 196848 3754
rect 197784 3726 197952 3754
rect 183714 190 183968 218
rect 183714 -960 183826 190
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195440 218 195468 3726
rect 196820 480 196848 3726
rect 197924 480 197952 3726
rect 198936 3726 199008 3754
rect 200084 3754 200112 4012
rect 201280 3754 201308 4012
rect 202476 3754 202504 4012
rect 203580 3754 203608 4012
rect 204776 3754 204804 4012
rect 205880 3754 205908 4012
rect 207076 3754 207104 4012
rect 208272 3754 208300 4012
rect 209376 3754 209404 4012
rect 210572 3754 210600 4012
rect 211676 3754 211704 4012
rect 212872 3754 212900 4012
rect 214068 3754 214096 4012
rect 215172 3754 215200 4012
rect 216368 3806 216396 4012
rect 216356 3800 216408 3806
rect 200084 3726 200344 3754
rect 201280 3726 201356 3754
rect 202476 3726 202736 3754
rect 203580 3726 203656 3754
rect 204776 3726 205128 3754
rect 205880 3726 206232 3754
rect 207076 3726 207152 3754
rect 208272 3726 208624 3754
rect 209376 3726 209728 3754
rect 210572 3726 211016 3754
rect 211676 3726 211752 3754
rect 212872 3726 213408 3754
rect 214068 3726 214512 3754
rect 215172 3726 215248 3754
rect 216356 3742 216408 3748
rect 216864 3800 216916 3806
rect 216864 3742 216916 3748
rect 217472 3754 217500 4012
rect 218668 3754 218696 4012
rect 219864 3754 219892 4012
rect 220968 3754 220996 4012
rect 222164 3806 222192 4012
rect 222152 3800 222204 3806
rect 195582 218 195694 480
rect 195440 190 195694 218
rect 195582 -960 195694 190
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198936 218 198964 3726
rect 200316 480 200344 3726
rect 199078 218 199190 480
rect 198936 190 199190 218
rect 199078 -960 199190 190
rect 200274 -960 200386 480
rect 201328 354 201356 3726
rect 202708 480 202736 3726
rect 201470 354 201582 480
rect 201328 326 201582 354
rect 201470 -960 201582 326
rect 202666 -960 202778 480
rect 203628 354 203656 3726
rect 205100 480 205128 3726
rect 206204 480 206232 3726
rect 203862 354 203974 480
rect 203628 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207124 354 207152 3726
rect 208596 480 208624 3726
rect 209700 626 209728 3726
rect 209700 598 209774 626
rect 209746 480 209774 598
rect 210988 480 211016 3726
rect 207358 354 207470 480
rect 207124 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209746 326 209862 480
rect 209750 -960 209862 326
rect 210946 -960 211058 480
rect 211724 354 211752 3726
rect 213380 480 213408 3726
rect 214484 480 214512 3726
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215220 354 215248 3726
rect 216876 480 216904 3742
rect 217472 3726 217640 3754
rect 218668 3726 219296 3754
rect 219864 3726 220032 3754
rect 220968 3726 221136 3754
rect 222152 3742 222204 3748
rect 222752 3800 222804 3806
rect 222752 3742 222804 3748
rect 223360 3754 223388 4012
rect 224464 3806 224492 4012
rect 224452 3800 224504 3806
rect 215638 354 215750 480
rect 215220 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 217612 354 217640 3726
rect 219268 480 219296 3726
rect 218030 354 218142 480
rect 217612 326 218142 354
rect 218030 -960 218142 326
rect 219226 -960 219338 480
rect 220004 354 220032 3726
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 3726
rect 222764 480 222792 3742
rect 223360 3726 223528 3754
rect 224452 3742 224504 3748
rect 225144 3800 225196 3806
rect 225144 3742 225196 3748
rect 225660 3754 225688 4012
rect 226764 3754 226792 4012
rect 227960 3754 227988 4012
rect 229156 3754 229184 4012
rect 230260 3806 230288 4012
rect 231456 3806 231484 4012
rect 232560 3806 232588 4012
rect 233756 3806 233784 4012
rect 230248 3800 230300 3806
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223500 354 223528 3726
rect 225156 480 225184 3742
rect 225660 3726 225920 3754
rect 226764 3726 227576 3754
rect 227960 3726 228312 3754
rect 229156 3726 229416 3754
rect 230248 3742 230300 3748
rect 231032 3800 231084 3806
rect 231032 3742 231084 3748
rect 231444 3800 231496 3806
rect 231444 3742 231496 3748
rect 232228 3800 232280 3806
rect 232228 3742 232280 3748
rect 232548 3800 232600 3806
rect 232548 3742 232600 3748
rect 233424 3800 233476 3806
rect 233424 3742 233476 3748
rect 233744 3800 233796 3806
rect 233744 3742 233796 3748
rect 234620 3800 234672 3806
rect 234620 3742 234672 3748
rect 234952 3754 234980 4012
rect 236056 3754 236084 4012
rect 237252 3806 237280 4012
rect 238356 3806 238384 4012
rect 239552 3806 239580 4012
rect 240748 3806 240776 4012
rect 241852 3806 241880 4012
rect 237240 3800 237292 3806
rect 223918 354 224030 480
rect 223500 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 225892 354 225920 3726
rect 227548 480 227576 3726
rect 226310 354 226422 480
rect 225892 326 226422 354
rect 226310 -960 226422 326
rect 227506 -960 227618 480
rect 228284 354 228312 3726
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 3726
rect 231044 480 231072 3742
rect 232240 480 232268 3742
rect 233436 480 233464 3742
rect 234632 480 234660 3742
rect 234952 3726 235856 3754
rect 236056 3726 236592 3754
rect 237240 3742 237292 3748
rect 238116 3800 238168 3806
rect 238116 3742 238168 3748
rect 238344 3800 238396 3806
rect 238344 3742 238396 3748
rect 239312 3800 239364 3806
rect 239312 3742 239364 3748
rect 239540 3800 239592 3806
rect 239540 3742 239592 3748
rect 240508 3800 240560 3806
rect 240508 3742 240560 3748
rect 240736 3800 240788 3806
rect 240736 3742 240788 3748
rect 241704 3800 241756 3806
rect 241704 3742 241756 3748
rect 241840 3800 241892 3806
rect 241840 3742 241892 3748
rect 242900 3800 242952 3806
rect 242900 3742 242952 3748
rect 243048 3754 243076 4012
rect 244152 3874 244180 4012
rect 244140 3868 244192 3874
rect 244140 3810 244192 3816
rect 245200 3868 245252 3874
rect 245200 3810 245252 3816
rect 235828 480 235856 3726
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 3726
rect 238128 480 238156 3742
rect 239324 480 239352 3742
rect 240520 480 240548 3742
rect 241716 480 241744 3742
rect 242912 480 242940 3742
rect 243048 3726 244136 3754
rect 244108 480 244136 3726
rect 245212 480 245240 3810
rect 245348 3806 245376 4012
rect 246544 3806 246572 4012
rect 247648 3942 247676 4012
rect 247636 3936 247688 3942
rect 247636 3878 247688 3884
rect 248604 3936 248656 3942
rect 248604 3878 248656 3884
rect 248844 3890 248872 4012
rect 245336 3800 245388 3806
rect 245336 3742 245388 3748
rect 246396 3800 246448 3806
rect 246396 3742 246448 3748
rect 246532 3800 246584 3806
rect 246532 3742 246584 3748
rect 247592 3800 247644 3806
rect 247592 3742 247644 3748
rect 246408 480 246436 3742
rect 247604 480 247632 3742
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 236982 -960 237094 326
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248616 354 248644 3878
rect 248844 3862 248920 3890
rect 248892 2854 248920 3862
rect 250040 3806 250068 4012
rect 251144 3890 251172 4012
rect 251100 3862 251172 3890
rect 250028 3800 250080 3806
rect 250028 3742 250080 3748
rect 251100 2854 251128 3862
rect 252340 3806 252368 4012
rect 253444 3890 253472 4012
rect 254640 3890 254668 4012
rect 253400 3862 253472 3890
rect 254596 3862 254668 3890
rect 251180 3800 251232 3806
rect 251180 3742 251232 3748
rect 252328 3800 252380 3806
rect 252328 3742 252380 3748
rect 248880 2848 248932 2854
rect 248880 2790 248932 2796
rect 249984 2848 250036 2854
rect 249984 2790 250036 2796
rect 251088 2848 251140 2854
rect 251088 2790 251140 2796
rect 249996 480 250024 2790
rect 251192 480 251220 3742
rect 253400 2922 253428 3862
rect 253480 3800 253532 3806
rect 253480 3742 253532 3748
rect 253388 2916 253440 2922
rect 253388 2858 253440 2864
rect 252376 2848 252428 2854
rect 252376 2790 252428 2796
rect 252388 480 252416 2790
rect 253492 480 253520 3742
rect 254596 2854 254624 3862
rect 255836 3806 255864 4012
rect 256940 3874 256968 4012
rect 256928 3868 256980 3874
rect 256928 3810 256980 3816
rect 258136 3806 258164 4012
rect 259240 3874 259268 4012
rect 258264 3868 258316 3874
rect 258264 3810 258316 3816
rect 259228 3868 259280 3874
rect 259228 3810 259280 3816
rect 255824 3800 255876 3806
rect 255824 3742 255876 3748
rect 257068 3800 257120 3806
rect 257068 3742 257120 3748
rect 258124 3800 258176 3806
rect 258124 3742 258176 3748
rect 254676 2916 254728 2922
rect 254676 2858 254728 2864
rect 254584 2848 254636 2854
rect 254584 2790 254636 2796
rect 254688 480 254716 2858
rect 255872 2848 255924 2854
rect 255872 2790 255924 2796
rect 255884 480 255912 2790
rect 257080 480 257108 3742
rect 258276 480 258304 3810
rect 260436 3806 260464 4012
rect 261632 3874 261660 4012
rect 260656 3868 260708 3874
rect 260656 3810 260708 3816
rect 261620 3868 261672 3874
rect 261620 3810 261672 3816
rect 259460 3800 259512 3806
rect 259460 3742 259512 3748
rect 260424 3800 260476 3806
rect 260424 3742 260476 3748
rect 259472 480 259500 3742
rect 260668 480 260696 3810
rect 262736 3806 262764 4012
rect 263932 3874 263960 4012
rect 262956 3868 263008 3874
rect 262956 3810 263008 3816
rect 263920 3868 263972 3874
rect 263920 3810 263972 3816
rect 261760 3800 261812 3806
rect 261760 3742 261812 3748
rect 262724 3800 262776 3806
rect 262724 3742 262776 3748
rect 261772 480 261800 3742
rect 262968 480 262996 3810
rect 265036 3806 265064 4012
rect 265348 3868 265400 3874
rect 265348 3810 265400 3816
rect 264152 3800 264204 3806
rect 264152 3742 264204 3748
rect 265024 3800 265076 3806
rect 265024 3742 265076 3748
rect 264164 480 264192 3742
rect 265360 480 265388 3810
rect 266232 3754 266260 4012
rect 267428 3806 267456 4012
rect 268532 3874 268560 4012
rect 268520 3868 268572 3874
rect 268520 3810 268572 3816
rect 269728 3806 269756 4012
rect 270832 3874 270860 4012
rect 270040 3868 270092 3874
rect 270040 3810 270092 3816
rect 270820 3868 270872 3874
rect 270820 3810 270872 3816
rect 266544 3800 266596 3806
rect 266232 3726 266308 3754
rect 266544 3742 266596 3748
rect 267416 3800 267468 3806
rect 267416 3742 267468 3748
rect 268844 3800 268896 3806
rect 268844 3742 268896 3748
rect 269716 3800 269768 3806
rect 269716 3742 269768 3748
rect 266280 1358 266308 3726
rect 266268 1352 266320 1358
rect 266268 1294 266320 1300
rect 266556 480 266584 3742
rect 267740 1352 267792 1358
rect 267740 1294 267792 1300
rect 267752 480 267780 1294
rect 268856 480 268884 3742
rect 270052 480 270080 3810
rect 272028 3806 272056 4012
rect 272432 3868 272484 3874
rect 272432 3810 272484 3816
rect 271236 3800 271288 3806
rect 271236 3742 271288 3748
rect 272016 3800 272068 3806
rect 272016 3742 272068 3748
rect 271248 480 271276 3742
rect 272444 480 272472 3810
rect 273224 3754 273252 4012
rect 273180 3726 273252 3754
rect 273628 3800 273680 3806
rect 273628 3742 273680 3748
rect 274328 3754 274356 4012
rect 275524 3874 275552 4012
rect 275512 3868 275564 3874
rect 275512 3810 275564 3816
rect 276720 3806 276748 4012
rect 277824 3874 277852 4012
rect 277124 3868 277176 3874
rect 277124 3810 277176 3816
rect 277812 3868 277864 3874
rect 277812 3810 277864 3816
rect 276708 3800 276760 3806
rect 273180 1358 273208 3726
rect 273168 1352 273220 1358
rect 273168 1294 273220 1300
rect 273640 480 273668 3742
rect 274328 3726 274404 3754
rect 276708 3742 276760 3748
rect 274376 746 274404 3726
rect 274824 1352 274876 1358
rect 274824 1294 274876 1300
rect 274364 740 274416 746
rect 274364 682 274416 688
rect 274836 480 274864 1294
rect 276020 740 276072 746
rect 276020 682 276072 688
rect 276032 480 276060 682
rect 277136 480 277164 3810
rect 279020 3806 279048 4012
rect 279516 3868 279568 3874
rect 279516 3810 279568 3816
rect 278320 3800 278372 3806
rect 278320 3742 278372 3748
rect 279008 3800 279060 3806
rect 279008 3742 279060 3748
rect 278332 480 278360 3742
rect 279528 480 279556 3810
rect 280124 3754 280152 4012
rect 280080 3726 280152 3754
rect 280712 3800 280764 3806
rect 280712 3742 280764 3748
rect 281320 3754 281348 4012
rect 282516 3754 282544 4012
rect 283620 3806 283648 4012
rect 284816 3874 284844 4012
rect 285920 3942 285948 4012
rect 285908 3936 285960 3942
rect 285908 3878 285960 3884
rect 284804 3868 284856 3874
rect 284804 3810 284856 3816
rect 286600 3868 286652 3874
rect 286600 3810 286652 3816
rect 283608 3800 283660 3806
rect 280080 1358 280108 3726
rect 280068 1352 280120 1358
rect 280068 1294 280120 1300
rect 280724 480 280752 3742
rect 281320 3726 281396 3754
rect 282516 3726 282592 3754
rect 283608 3742 283660 3748
rect 285404 3800 285456 3806
rect 285404 3742 285456 3748
rect 281368 1290 281396 3726
rect 282564 1358 282592 3726
rect 281908 1352 281960 1358
rect 281908 1294 281960 1300
rect 282552 1352 282604 1358
rect 282552 1294 282604 1300
rect 284300 1352 284352 1358
rect 284300 1294 284352 1300
rect 281356 1284 281408 1290
rect 281356 1226 281408 1232
rect 281920 480 281948 1294
rect 283104 1284 283156 1290
rect 283104 1226 283156 1232
rect 283116 480 283144 1226
rect 284312 480 284340 1294
rect 285416 480 285444 3742
rect 286612 480 286640 3810
rect 287116 3806 287144 4012
rect 287796 3936 287848 3942
rect 287796 3878 287848 3884
rect 287104 3800 287156 3806
rect 287104 3742 287156 3748
rect 287808 480 287836 3878
rect 288312 3754 288340 4012
rect 288992 3800 289044 3806
rect 288312 3726 288388 3754
rect 288992 3742 289044 3748
rect 289416 3754 289444 4012
rect 290612 3754 290640 4012
rect 291716 3806 291744 4012
rect 292912 3874 292940 4012
rect 292900 3868 292952 3874
rect 292900 3810 292952 3816
rect 294108 3806 294136 4012
rect 294880 3868 294932 3874
rect 294880 3810 294932 3816
rect 291704 3800 291756 3806
rect 288360 1358 288388 3726
rect 288348 1352 288400 1358
rect 288348 1294 288400 1300
rect 289004 480 289032 3742
rect 289416 3726 289492 3754
rect 290612 3726 290688 3754
rect 291704 3742 291756 3748
rect 293684 3800 293736 3806
rect 293684 3742 293736 3748
rect 294096 3800 294148 3806
rect 294096 3742 294148 3748
rect 289464 1290 289492 3726
rect 290188 1352 290240 1358
rect 290188 1294 290240 1300
rect 289452 1284 289504 1290
rect 289452 1226 289504 1232
rect 290200 480 290228 1294
rect 290660 610 290688 3726
rect 291384 1284 291436 1290
rect 291384 1226 291436 1232
rect 290648 604 290700 610
rect 290648 546 290700 552
rect 291396 480 291424 1226
rect 292580 604 292632 610
rect 292580 546 292632 552
rect 292592 480 292620 546
rect 293696 480 293724 3742
rect 294892 480 294920 3810
rect 295212 3754 295240 4012
rect 296076 3800 296128 3806
rect 295212 3726 295288 3754
rect 296076 3742 296128 3748
rect 296408 3754 296436 4012
rect 297512 3754 297540 4012
rect 298708 3806 298736 4012
rect 299904 3874 299932 4012
rect 299892 3868 299944 3874
rect 299892 3810 299944 3816
rect 301008 3806 301036 4012
rect 301964 3868 302016 3874
rect 301964 3810 302016 3816
rect 298696 3800 298748 3806
rect 295260 1358 295288 3726
rect 295248 1352 295300 1358
rect 295248 1294 295300 1300
rect 296088 480 296116 3742
rect 296408 3726 296484 3754
rect 297512 3726 297588 3754
rect 298696 3742 298748 3748
rect 300768 3800 300820 3806
rect 300768 3742 300820 3748
rect 300996 3800 301048 3806
rect 300996 3742 301048 3748
rect 296456 1290 296484 3726
rect 297560 1358 297588 3726
rect 297272 1352 297324 1358
rect 297272 1294 297324 1300
rect 297548 1352 297600 1358
rect 297548 1294 297600 1300
rect 299664 1352 299716 1358
rect 299664 1294 299716 1300
rect 296444 1284 296496 1290
rect 296444 1226 296496 1232
rect 297284 480 297312 1294
rect 298468 1284 298520 1290
rect 298468 1226 298520 1232
rect 298480 480 298508 1226
rect 299676 480 299704 1294
rect 300780 480 300808 3742
rect 301976 480 302004 3810
rect 302204 3754 302232 4012
rect 302160 3726 302232 3754
rect 303160 3800 303212 3806
rect 303160 3742 303212 3748
rect 303308 3754 303336 4012
rect 304504 3754 304532 4012
rect 305700 3754 305728 4012
rect 306804 3874 306832 4012
rect 306792 3868 306844 3874
rect 306792 3810 306844 3816
rect 308000 3806 308028 4012
rect 309048 3868 309100 3874
rect 309048 3810 309100 3816
rect 307988 3800 308040 3806
rect 302160 1358 302188 3726
rect 302148 1352 302200 1358
rect 302148 1294 302200 1300
rect 303172 480 303200 3742
rect 303308 3726 303384 3754
rect 304504 3726 304580 3754
rect 305700 3726 305776 3754
rect 307988 3742 308040 3748
rect 303356 1290 303384 3726
rect 304356 1352 304408 1358
rect 304356 1294 304408 1300
rect 303344 1284 303396 1290
rect 303344 1226 303396 1232
rect 304368 480 304396 1294
rect 304552 610 304580 3726
rect 305748 1358 305776 3726
rect 305736 1352 305788 1358
rect 305736 1294 305788 1300
rect 307944 1352 307996 1358
rect 307944 1294 307996 1300
rect 305552 1284 305604 1290
rect 305552 1226 305604 1232
rect 304540 604 304592 610
rect 304540 546 304592 552
rect 305564 480 305592 1226
rect 306748 604 306800 610
rect 306748 546 306800 552
rect 306760 480 306788 546
rect 307956 480 307984 1294
rect 309060 480 309088 3810
rect 309196 3754 309224 4012
rect 310300 3890 310328 4012
rect 311496 3890 311524 4012
rect 310300 3862 310376 3890
rect 311496 3862 311572 3890
rect 310244 3800 310296 3806
rect 309196 3726 309272 3754
rect 310244 3742 310296 3748
rect 309244 2854 309272 3726
rect 309232 2848 309284 2854
rect 309232 2790 309284 2796
rect 310256 480 310284 3742
rect 310348 1358 310376 3862
rect 311440 2848 311492 2854
rect 311440 2790 311492 2796
rect 310336 1352 310388 1358
rect 310336 1294 310388 1300
rect 311452 480 311480 2790
rect 311544 1222 311572 3862
rect 312600 3754 312628 4012
rect 312556 3726 312628 3754
rect 313796 3754 313824 4012
rect 314992 3754 315020 4012
rect 316096 3806 316124 4012
rect 316084 3800 316136 3806
rect 313796 3726 313872 3754
rect 314992 3726 315068 3754
rect 317292 3754 317320 4012
rect 316084 3742 316136 3748
rect 312556 1290 312584 3726
rect 313844 1358 313872 3726
rect 315040 2854 315068 3726
rect 317248 3726 317320 3754
rect 318396 3754 318424 4012
rect 318524 3800 318576 3806
rect 318396 3726 318472 3754
rect 318524 3742 318576 3748
rect 319592 3754 319620 4012
rect 320788 3754 320816 4012
rect 321892 3754 321920 4012
rect 323088 3806 323116 4012
rect 323076 3800 323128 3806
rect 315028 2848 315080 2854
rect 315028 2790 315080 2796
rect 317248 1358 317276 3726
rect 317328 2848 317380 2854
rect 317328 2790 317380 2796
rect 312636 1352 312688 1358
rect 312636 1294 312688 1300
rect 313832 1352 313884 1358
rect 313832 1294 313884 1300
rect 316224 1352 316276 1358
rect 316224 1294 316276 1300
rect 317236 1352 317288 1358
rect 317236 1294 317288 1300
rect 312544 1284 312596 1290
rect 312544 1226 312596 1232
rect 311532 1216 311584 1222
rect 311532 1158 311584 1164
rect 312648 480 312676 1294
rect 315028 1284 315080 1290
rect 315028 1226 315080 1232
rect 313832 1216 313884 1222
rect 313832 1158 313884 1164
rect 313844 480 313872 1158
rect 315040 480 315068 1226
rect 316236 480 316264 1294
rect 317340 480 317368 2790
rect 318444 1290 318472 3726
rect 318432 1284 318484 1290
rect 318432 1226 318484 1232
rect 318536 480 318564 3742
rect 319592 3726 319668 3754
rect 320788 3726 320864 3754
rect 321892 3726 321968 3754
rect 323076 3742 323128 3748
rect 324192 3754 324220 4012
rect 325388 3754 325416 4012
rect 325608 3800 325660 3806
rect 324192 3726 324268 3754
rect 325388 3726 325464 3754
rect 325608 3742 325660 3748
rect 326584 3754 326612 4012
rect 327688 3754 327716 4012
rect 328884 3754 328912 4012
rect 329988 3754 330016 4012
rect 331184 3754 331212 4012
rect 319640 1222 319668 3726
rect 319720 1352 319772 1358
rect 319720 1294 319772 1300
rect 319628 1216 319680 1222
rect 319628 1158 319680 1164
rect 319732 480 319760 1294
rect 320836 1154 320864 3726
rect 321940 1358 321968 3726
rect 321928 1352 321980 1358
rect 321928 1294 321980 1300
rect 324240 1290 324268 3726
rect 325436 1358 325464 3726
rect 324412 1352 324464 1358
rect 324412 1294 324464 1300
rect 325424 1352 325476 1358
rect 325424 1294 325476 1300
rect 320916 1284 320968 1290
rect 320916 1226 320968 1232
rect 324228 1284 324280 1290
rect 324228 1226 324280 1232
rect 320824 1148 320876 1154
rect 320824 1090 320876 1096
rect 320928 480 320956 1226
rect 322112 1216 322164 1222
rect 322112 1158 322164 1164
rect 322124 480 322152 1158
rect 323308 1148 323360 1154
rect 323308 1090 323360 1096
rect 323320 480 323348 1090
rect 324424 480 324452 1294
rect 325620 480 325648 3742
rect 326584 3726 326660 3754
rect 327688 3726 327764 3754
rect 328884 3726 328960 3754
rect 329988 3726 330064 3754
rect 326632 1222 326660 3726
rect 326804 1284 326856 1290
rect 326804 1226 326856 1232
rect 326620 1216 326672 1222
rect 326620 1158 326672 1164
rect 326816 480 326844 1226
rect 327736 1154 327764 3726
rect 328932 1358 328960 3726
rect 328000 1352 328052 1358
rect 328000 1294 328052 1300
rect 328920 1352 328972 1358
rect 328920 1294 328972 1300
rect 327724 1148 327776 1154
rect 327724 1090 327776 1096
rect 328012 480 328040 1294
rect 330036 1290 330064 3726
rect 331140 3726 331212 3754
rect 332380 3754 332408 4012
rect 333484 3754 333512 4012
rect 334680 3754 334708 4012
rect 335876 3754 335904 4012
rect 336980 3754 337008 4012
rect 338176 3754 338204 4012
rect 339280 3754 339308 4012
rect 340476 3754 340504 4012
rect 341672 3754 341700 4012
rect 342776 3754 342804 4012
rect 343972 3754 344000 4012
rect 345076 3754 345104 4012
rect 346272 3754 346300 4012
rect 347468 3754 347496 4012
rect 348572 3754 348600 4012
rect 349768 3754 349796 4012
rect 350872 3754 350900 4012
rect 352068 3754 352096 4012
rect 353264 3754 353292 4012
rect 332380 3726 332456 3754
rect 333484 3726 333560 3754
rect 334680 3726 334756 3754
rect 335876 3726 335952 3754
rect 336980 3726 337056 3754
rect 338176 3726 338252 3754
rect 339280 3726 339356 3754
rect 340476 3726 340552 3754
rect 341672 3726 341748 3754
rect 342776 3726 342852 3754
rect 343972 3726 344048 3754
rect 345076 3726 345152 3754
rect 346272 3726 346348 3754
rect 347468 3726 347544 3754
rect 348572 3726 348648 3754
rect 349768 3726 349844 3754
rect 350872 3726 350948 3754
rect 352068 3726 352144 3754
rect 330024 1284 330076 1290
rect 330024 1226 330076 1232
rect 331140 1222 331168 3726
rect 332428 1358 332456 3726
rect 331588 1352 331640 1358
rect 331588 1294 331640 1300
rect 332416 1352 332468 1358
rect 332416 1294 332468 1300
rect 329196 1216 329248 1222
rect 329196 1158 329248 1164
rect 331128 1216 331180 1222
rect 331128 1158 331180 1164
rect 329208 480 329236 1158
rect 330392 1148 330444 1154
rect 330392 1090 330444 1096
rect 330404 480 330432 1090
rect 331600 480 331628 1294
rect 332692 1284 332744 1290
rect 332692 1226 332744 1232
rect 332704 480 332732 1226
rect 333532 746 333560 3726
rect 334728 1290 334756 3726
rect 335924 1358 335952 3726
rect 335084 1352 335136 1358
rect 335084 1294 335136 1300
rect 335912 1352 335964 1358
rect 335912 1294 335964 1300
rect 334716 1284 334768 1290
rect 334716 1226 334768 1232
rect 333888 1216 333940 1222
rect 333888 1158 333940 1164
rect 333520 740 333572 746
rect 333520 682 333572 688
rect 333900 480 333928 1158
rect 335096 480 335124 1294
rect 337028 1222 337056 3726
rect 337476 1284 337528 1290
rect 337476 1226 337528 1232
rect 337016 1216 337068 1222
rect 337016 1158 337068 1164
rect 336280 740 336332 746
rect 336280 682 336332 688
rect 336292 480 336320 682
rect 337488 480 337516 1226
rect 338224 746 338252 3726
rect 339328 1358 339356 3726
rect 338672 1352 338724 1358
rect 338672 1294 338724 1300
rect 339316 1352 339368 1358
rect 339316 1294 339368 1300
rect 338212 740 338264 746
rect 338212 682 338264 688
rect 338684 480 338712 1294
rect 340524 1290 340552 3726
rect 340512 1284 340564 1290
rect 340512 1226 340564 1232
rect 341720 1222 341748 3726
rect 342168 1352 342220 1358
rect 342168 1294 342220 1300
rect 339868 1216 339920 1222
rect 339868 1158 339920 1164
rect 341708 1216 341760 1222
rect 341708 1158 341760 1164
rect 339880 480 339908 1158
rect 340972 740 341024 746
rect 340972 682 341024 688
rect 340984 480 341012 682
rect 342180 480 342208 1294
rect 342824 746 342852 3726
rect 344020 1290 344048 3726
rect 345124 1358 345152 3726
rect 345112 1352 345164 1358
rect 345112 1294 345164 1300
rect 343364 1284 343416 1290
rect 343364 1226 343416 1232
rect 344008 1284 344060 1290
rect 344008 1226 344060 1232
rect 342812 740 342864 746
rect 342812 682 342864 688
rect 343376 480 343404 1226
rect 344560 1216 344612 1222
rect 344560 1158 344612 1164
rect 344572 480 344600 1158
rect 346320 746 346348 3726
rect 346952 1284 347004 1290
rect 346952 1226 347004 1232
rect 345756 740 345808 746
rect 345756 682 345808 688
rect 346308 740 346360 746
rect 346308 682 346360 688
rect 345768 480 345796 682
rect 346964 480 346992 1226
rect 347516 882 347544 3726
rect 348056 1352 348108 1358
rect 348056 1294 348108 1300
rect 347504 876 347556 882
rect 347504 818 347556 824
rect 348068 480 348096 1294
rect 348620 1290 348648 3726
rect 349816 1358 349844 3726
rect 349804 1352 349856 1358
rect 349804 1294 349856 1300
rect 348608 1284 348660 1290
rect 348608 1226 348660 1232
rect 350448 876 350500 882
rect 350448 818 350500 824
rect 349252 740 349304 746
rect 349252 682 349304 688
rect 349264 480 349292 682
rect 350460 480 350488 818
rect 350920 746 350948 3726
rect 352116 1290 352144 3726
rect 353220 3726 353292 3754
rect 354368 3754 354396 4012
rect 355564 3754 355592 4012
rect 356668 3754 356696 4012
rect 357864 3754 357892 4012
rect 359060 3754 359088 4012
rect 360164 3754 360192 4012
rect 354368 3726 354444 3754
rect 355564 3726 355640 3754
rect 356668 3726 356744 3754
rect 357864 3726 357940 3754
rect 359060 3726 359136 3754
rect 353220 1358 353248 3726
rect 352840 1352 352892 1358
rect 352840 1294 352892 1300
rect 353208 1352 353260 1358
rect 353208 1294 353260 1300
rect 351644 1284 351696 1290
rect 351644 1226 351696 1232
rect 352104 1284 352156 1290
rect 352104 1226 352156 1232
rect 350908 740 350960 746
rect 350908 682 350960 688
rect 351656 480 351684 1226
rect 352852 480 352880 1294
rect 354036 740 354088 746
rect 354036 682 354088 688
rect 354048 480 354076 682
rect 248758 354 248870 480
rect 248616 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 354416 66 354444 3726
rect 355612 1290 355640 3726
rect 356716 1358 356744 3726
rect 356336 1352 356388 1358
rect 356336 1294 356388 1300
rect 356704 1352 356756 1358
rect 356704 1294 356756 1300
rect 355232 1284 355284 1290
rect 355232 1226 355284 1232
rect 355600 1284 355652 1290
rect 355600 1226 355652 1232
rect 355244 480 355272 1226
rect 356348 480 356376 1294
rect 357912 1222 357940 3726
rect 359108 1290 359136 3726
rect 360120 3726 360192 3754
rect 361360 3754 361388 4012
rect 362556 3754 362584 4012
rect 363660 3754 363688 4012
rect 364856 3754 364884 4012
rect 365960 3754 365988 4012
rect 367156 3754 367184 4012
rect 368352 3754 368380 4012
rect 369456 3754 369484 4012
rect 370652 3754 370680 4012
rect 371756 3754 371784 4012
rect 372952 3754 372980 4012
rect 374148 3754 374176 4012
rect 375252 3754 375280 4012
rect 376448 3754 376476 4012
rect 361360 3726 361436 3754
rect 362556 3726 362632 3754
rect 363660 3726 363736 3754
rect 364856 3726 364932 3754
rect 365960 3726 366036 3754
rect 367156 3726 367232 3754
rect 368352 3726 368428 3754
rect 369456 3726 369532 3754
rect 370652 3726 370728 3754
rect 371756 3726 371832 3754
rect 372952 3726 373028 3754
rect 374148 3726 374224 3754
rect 375252 3726 375328 3754
rect 359924 1352 359976 1358
rect 359924 1294 359976 1300
rect 358728 1284 358780 1290
rect 358728 1226 358780 1232
rect 359096 1284 359148 1290
rect 359096 1226 359148 1232
rect 357900 1216 357952 1222
rect 357900 1158 357952 1164
rect 358740 480 358768 1226
rect 359936 480 359964 1294
rect 360120 1154 360148 3726
rect 361120 1216 361172 1222
rect 361120 1158 361172 1164
rect 360108 1148 360160 1154
rect 360108 1090 360160 1096
rect 361132 480 361160 1158
rect 361408 882 361436 3726
rect 362604 1358 362632 3726
rect 362592 1352 362644 1358
rect 362592 1294 362644 1300
rect 363708 1290 363736 3726
rect 362316 1284 362368 1290
rect 362316 1226 362368 1232
rect 363696 1284 363748 1290
rect 363696 1226 363748 1232
rect 361396 876 361448 882
rect 361396 818 361448 824
rect 362328 480 362356 1226
rect 364904 1222 364932 3726
rect 365812 1352 365864 1358
rect 365812 1294 365864 1300
rect 364892 1216 364944 1222
rect 364892 1158 364944 1164
rect 363512 1148 363564 1154
rect 363512 1090 363564 1096
rect 363524 480 363552 1090
rect 364616 876 364668 882
rect 364616 818 364668 824
rect 364628 480 364656 818
rect 365824 480 365852 1294
rect 366008 746 366036 3726
rect 367204 1358 367232 3726
rect 367192 1352 367244 1358
rect 367192 1294 367244 1300
rect 367008 1284 367060 1290
rect 367008 1226 367060 1232
rect 365996 740 366048 746
rect 365996 682 366048 688
rect 367020 480 367048 1226
rect 368204 1216 368256 1222
rect 368204 1158 368256 1164
rect 368216 480 368244 1158
rect 368400 882 368428 3726
rect 368388 876 368440 882
rect 368388 818 368440 824
rect 369504 746 369532 3726
rect 370700 1358 370728 3726
rect 370596 1352 370648 1358
rect 370596 1294 370648 1300
rect 370688 1352 370740 1358
rect 370688 1294 370740 1300
rect 369400 740 369452 746
rect 369400 682 369452 688
rect 369492 740 369544 746
rect 369492 682 369544 688
rect 369412 480 369440 682
rect 370608 480 370636 1294
rect 371804 882 371832 3726
rect 373000 1290 373028 3726
rect 374092 1352 374144 1358
rect 374092 1294 374144 1300
rect 372988 1284 373040 1290
rect 372988 1226 373040 1232
rect 371700 876 371752 882
rect 371700 818 371752 824
rect 371792 876 371844 882
rect 371792 818 371844 824
rect 371712 480 371740 818
rect 372896 740 372948 746
rect 372896 682 372948 688
rect 372908 480 372936 682
rect 374104 480 374132 1294
rect 374196 1018 374224 3726
rect 375300 1222 375328 3726
rect 376404 3726 376476 3754
rect 377552 3754 377580 4012
rect 378748 3754 378776 4012
rect 379944 3754 379972 4012
rect 377552 3726 377628 3754
rect 378748 3726 378824 3754
rect 376404 1358 376432 3726
rect 376392 1352 376444 1358
rect 376392 1294 376444 1300
rect 377600 1290 377628 3726
rect 376484 1284 376536 1290
rect 376484 1226 376536 1232
rect 377588 1284 377640 1290
rect 377588 1226 377640 1232
rect 375288 1216 375340 1222
rect 375288 1158 375340 1164
rect 374184 1012 374236 1018
rect 374184 954 374236 960
rect 375288 876 375340 882
rect 375288 818 375340 824
rect 375300 480 375328 818
rect 376496 480 376524 1226
rect 378796 1086 378824 3726
rect 379900 3726 379972 3754
rect 381048 3754 381076 4012
rect 382244 3754 382272 4012
rect 381048 3726 381124 3754
rect 378876 1216 378928 1222
rect 378876 1158 378928 1164
rect 378784 1080 378836 1086
rect 378784 1022 378836 1028
rect 377680 1012 377732 1018
rect 377680 954 377732 960
rect 377692 480 377720 954
rect 378888 480 378916 1158
rect 379900 1018 379928 3726
rect 379980 1352 380032 1358
rect 379980 1294 380032 1300
rect 379888 1012 379940 1018
rect 379888 954 379940 960
rect 379992 480 380020 1294
rect 381096 1222 381124 3726
rect 382200 3726 382272 3754
rect 383348 3754 383376 4012
rect 384544 3754 384572 4012
rect 385740 3754 385768 4012
rect 386844 3754 386872 4012
rect 388040 3754 388068 4012
rect 389236 3754 389264 4012
rect 390340 3754 390368 4012
rect 391536 3754 391564 4012
rect 392640 3754 392668 4012
rect 393836 3754 393864 4012
rect 395032 3754 395060 4012
rect 396136 3754 396164 4012
rect 397332 3754 397360 4012
rect 398436 3754 398464 4012
rect 399632 3754 399660 4012
rect 400828 3754 400856 4012
rect 401932 3754 401960 4012
rect 403128 3754 403156 4012
rect 404232 3754 404260 4012
rect 405428 3754 405456 4012
rect 406624 3754 406652 4012
rect 407728 3754 407756 4012
rect 408924 3754 408952 4012
rect 410028 3754 410056 4012
rect 411224 3754 411252 4012
rect 383348 3726 383424 3754
rect 384544 3726 384620 3754
rect 385740 3726 385816 3754
rect 386844 3726 386920 3754
rect 388040 3726 388116 3754
rect 389236 3726 389312 3754
rect 390340 3726 390416 3754
rect 391536 3726 391612 3754
rect 392640 3726 392716 3754
rect 393836 3726 393912 3754
rect 395032 3726 395108 3754
rect 396136 3726 396212 3754
rect 397332 3726 397408 3754
rect 398436 3726 398512 3754
rect 399632 3726 399708 3754
rect 400828 3726 400904 3754
rect 401932 3726 402008 3754
rect 403128 3726 403204 3754
rect 404232 3726 404308 3754
rect 405428 3726 405504 3754
rect 406624 3726 406700 3754
rect 407728 3726 407804 3754
rect 408924 3726 409000 3754
rect 410028 3726 410104 3754
rect 381176 1284 381228 1290
rect 381176 1226 381228 1232
rect 381084 1216 381136 1222
rect 381084 1158 381136 1164
rect 381188 480 381216 1226
rect 382200 1154 382228 3726
rect 382188 1148 382240 1154
rect 382188 1090 382240 1096
rect 382372 1080 382424 1086
rect 382372 1022 382424 1028
rect 382384 480 382412 1022
rect 354404 60 354456 66
rect 354404 2 354456 8
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 82 357614 480
rect 357360 66 357614 82
rect 357348 60 357614 66
rect 357400 54 357614 60
rect 357348 2 357400 8
rect 357502 -960 357614 54
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383396 406 383424 3726
rect 383568 1012 383620 1018
rect 383568 954 383620 960
rect 383580 480 383608 954
rect 384592 882 384620 3726
rect 385788 1358 385816 3726
rect 385776 1352 385828 1358
rect 385776 1294 385828 1300
rect 384764 1216 384816 1222
rect 384764 1158 384816 1164
rect 384580 876 384632 882
rect 384580 818 384632 824
rect 384776 480 384804 1158
rect 385960 1148 386012 1154
rect 385960 1090 386012 1096
rect 385972 480 386000 1090
rect 386892 1086 386920 3726
rect 388088 1290 388116 3726
rect 388076 1284 388128 1290
rect 388076 1226 388128 1232
rect 389284 1154 389312 3726
rect 389456 1352 389508 1358
rect 389456 1294 389508 1300
rect 389272 1148 389324 1154
rect 389272 1090 389324 1096
rect 386880 1080 386932 1086
rect 386880 1022 386932 1028
rect 388260 876 388312 882
rect 388260 818 388312 824
rect 388272 480 388300 818
rect 389468 480 389496 1294
rect 390388 1222 390416 3726
rect 390376 1216 390428 1222
rect 390376 1158 390428 1164
rect 390652 1080 390704 1086
rect 390652 1022 390704 1028
rect 390664 480 390692 1022
rect 391584 882 391612 3726
rect 391848 1284 391900 1290
rect 391848 1226 391900 1232
rect 391572 876 391624 882
rect 391572 818 391624 824
rect 391860 480 391888 1226
rect 383384 400 383436 406
rect 383384 342 383436 348
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 386788 400 386840 406
rect 387126 354 387238 480
rect 386840 348 387238 354
rect 386788 342 387238 348
rect 386800 326 387238 342
rect 387126 -960 387238 326
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392688 270 392716 3726
rect 393884 1290 393912 3726
rect 395080 1358 395108 3726
rect 395068 1352 395120 1358
rect 395068 1294 395120 1300
rect 393872 1284 393924 1290
rect 393872 1226 393924 1232
rect 394240 1216 394292 1222
rect 394240 1158 394292 1164
rect 393044 1148 393096 1154
rect 393044 1090 393096 1096
rect 393056 480 393084 1090
rect 394252 480 394280 1158
rect 396184 882 396212 3726
rect 397380 1154 397408 3726
rect 398484 1290 398512 3726
rect 399680 1358 399708 3726
rect 398932 1352 398984 1358
rect 398932 1294 398984 1300
rect 399668 1352 399720 1358
rect 399668 1294 399720 1300
rect 397736 1284 397788 1290
rect 397736 1226 397788 1232
rect 398472 1284 398524 1290
rect 398472 1226 398524 1232
rect 397368 1148 397420 1154
rect 397368 1090 397420 1096
rect 395344 876 395396 882
rect 395344 818 395396 824
rect 396172 876 396224 882
rect 396172 818 396224 824
rect 395356 480 395384 818
rect 397748 480 397776 1226
rect 398944 480 398972 1294
rect 400876 1222 400904 3726
rect 400864 1216 400916 1222
rect 400864 1158 400916 1164
rect 401324 1148 401376 1154
rect 401324 1090 401376 1096
rect 400128 876 400180 882
rect 400128 818 400180 824
rect 400140 480 400168 818
rect 401336 480 401364 1090
rect 392676 264 392728 270
rect 392676 206 392728 212
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396172 264 396224 270
rect 396510 218 396622 480
rect 396224 212 396622 218
rect 396172 206 396622 212
rect 396184 190 396622 206
rect 396510 -960 396622 190
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 401980 66 402008 3726
rect 403176 1290 403204 3726
rect 403624 1352 403676 1358
rect 403624 1294 403676 1300
rect 402520 1284 402572 1290
rect 402520 1226 402572 1232
rect 403164 1284 403216 1290
rect 403164 1226 403216 1232
rect 402532 480 402560 1226
rect 403636 480 403664 1294
rect 404280 1154 404308 3726
rect 405476 1358 405504 3726
rect 405464 1352 405516 1358
rect 405464 1294 405516 1300
rect 404820 1216 404872 1222
rect 404820 1158 404872 1164
rect 404268 1148 404320 1154
rect 404268 1090 404320 1096
rect 404832 480 404860 1158
rect 406672 882 406700 3726
rect 407212 1284 407264 1290
rect 407212 1226 407264 1232
rect 406660 876 406712 882
rect 406660 818 406712 824
rect 407224 480 407252 1226
rect 407776 1222 407804 3726
rect 407764 1216 407816 1222
rect 407764 1158 407816 1164
rect 408972 1154 409000 3726
rect 409604 1352 409656 1358
rect 409604 1294 409656 1300
rect 408408 1148 408460 1154
rect 408408 1090 408460 1096
rect 408960 1148 409012 1154
rect 408960 1090 409012 1096
rect 408420 480 408448 1090
rect 409616 480 409644 1294
rect 410076 1290 410104 3726
rect 411180 3726 411252 3754
rect 412420 3754 412448 4012
rect 413524 3754 413552 4012
rect 414720 3754 414748 4012
rect 415916 3754 415944 4012
rect 417020 3754 417048 4012
rect 418216 3754 418244 4012
rect 419320 3754 419348 4012
rect 420516 3754 420544 4012
rect 421712 3754 421740 4012
rect 422816 3754 422844 4012
rect 424012 3754 424040 4012
rect 425116 3754 425144 4012
rect 426312 3754 426340 4012
rect 427508 3754 427536 4012
rect 428612 3754 428640 4012
rect 429808 3754 429836 4012
rect 430912 3754 430940 4012
rect 432108 3754 432136 4012
rect 433304 3754 433332 4012
rect 434408 3754 434436 4012
rect 412420 3726 412496 3754
rect 413524 3726 413600 3754
rect 414720 3726 414796 3754
rect 415916 3726 415992 3754
rect 417020 3726 417096 3754
rect 418216 3726 418292 3754
rect 419320 3726 419396 3754
rect 420516 3726 420592 3754
rect 421712 3726 421788 3754
rect 422816 3726 422892 3754
rect 424012 3726 424088 3754
rect 425116 3726 425192 3754
rect 426312 3726 426388 3754
rect 427508 3726 427584 3754
rect 428612 3726 428688 3754
rect 429808 3726 429884 3754
rect 430912 3726 431080 3754
rect 432108 3726 432184 3754
rect 411180 2854 411208 3726
rect 411168 2848 411220 2854
rect 411168 2790 411220 2796
rect 410064 1284 410116 1290
rect 410064 1226 410116 1232
rect 411904 1216 411956 1222
rect 411904 1158 411956 1164
rect 410800 876 410852 882
rect 410800 818 410852 824
rect 410812 480 410840 818
rect 411916 480 411944 1158
rect 401968 60 402020 66
rect 401968 2 402020 8
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 82 406098 480
rect 405986 66 406240 82
rect 405986 60 406252 66
rect 405986 54 406200 60
rect 405986 -960 406098 54
rect 406200 2 406252 8
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412468 270 412496 3726
rect 413572 1222 413600 3726
rect 414296 1284 414348 1290
rect 414296 1226 414348 1232
rect 413560 1216 413612 1222
rect 413560 1158 413612 1164
rect 413100 1148 413152 1154
rect 413100 1090 413152 1096
rect 413112 480 413140 1090
rect 414308 480 414336 1226
rect 414768 1018 414796 3726
rect 415492 2848 415544 2854
rect 415492 2790 415544 2796
rect 414756 1012 414808 1018
rect 414756 954 414808 960
rect 415504 480 415532 2790
rect 415964 1358 415992 3726
rect 415952 1352 416004 1358
rect 415952 1294 416004 1300
rect 417068 882 417096 3726
rect 418264 1290 418292 3726
rect 418252 1284 418304 1290
rect 418252 1226 418304 1232
rect 419368 1222 419396 3726
rect 420184 1352 420236 1358
rect 420184 1294 420236 1300
rect 417884 1216 417936 1222
rect 417884 1158 417936 1164
rect 419356 1216 419408 1222
rect 419356 1158 419408 1164
rect 417056 876 417108 882
rect 417056 818 417108 824
rect 417896 480 417924 1158
rect 418988 1012 419040 1018
rect 418988 954 419040 960
rect 419000 480 419028 954
rect 420196 480 420224 1294
rect 420564 1154 420592 3726
rect 420552 1148 420604 1154
rect 420552 1090 420604 1096
rect 421380 876 421432 882
rect 421380 818 421432 824
rect 421392 480 421420 818
rect 412456 264 412508 270
rect 412456 206 412508 212
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 218 416770 480
rect 416872 264 416924 270
rect 416658 212 416872 218
rect 416658 206 416924 212
rect 416658 190 416912 206
rect 416658 -960 416770 190
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 421760 270 421788 3726
rect 422576 1284 422628 1290
rect 422576 1226 422628 1232
rect 422588 480 422616 1226
rect 422864 1018 422892 3726
rect 424060 1290 424088 3726
rect 424048 1284 424100 1290
rect 424048 1226 424100 1232
rect 423404 1216 423456 1222
rect 423404 1158 423456 1164
rect 422852 1012 422904 1018
rect 422852 954 422904 960
rect 421748 264 421800 270
rect 421748 206 421800 212
rect 422546 -960 422658 480
rect 423416 354 423444 1158
rect 424968 1148 425020 1154
rect 424968 1090 425020 1096
rect 424980 480 425008 1090
rect 425164 1086 425192 3726
rect 426360 1222 426388 3726
rect 427556 1358 427584 3726
rect 427544 1352 427596 1358
rect 427544 1294 427596 1300
rect 428464 1284 428516 1290
rect 428464 1226 428516 1232
rect 426348 1216 426400 1222
rect 426348 1158 426400 1164
rect 425152 1080 425204 1086
rect 425152 1022 425204 1028
rect 427268 1012 427320 1018
rect 427268 954 427320 960
rect 427280 480 427308 954
rect 428476 480 428504 1226
rect 428660 1154 428688 3726
rect 428648 1148 428700 1154
rect 428648 1090 428700 1096
rect 429660 1080 429712 1086
rect 429660 1022 429712 1028
rect 429672 480 429700 1022
rect 429856 882 429884 3726
rect 430856 1216 430908 1222
rect 430856 1158 430908 1164
rect 429844 876 429896 882
rect 429844 818 429896 824
rect 430868 480 430896 1158
rect 423742 354 423854 480
rect 423416 326 423854 354
rect 423742 -960 423854 326
rect 424938 -960 425050 480
rect 425796 264 425848 270
rect 426134 218 426246 480
rect 425848 212 426246 218
rect 425796 206 426246 212
rect 425808 190 426246 206
rect 426134 -960 426246 190
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 431052 134 431080 3726
rect 431868 1352 431920 1358
rect 431868 1294 431920 1300
rect 431880 354 431908 1294
rect 432156 1018 432184 3726
rect 433260 3726 433332 3754
rect 434364 3726 434436 3754
rect 435604 3754 435632 4012
rect 436708 3754 436736 4012
rect 437904 3754 437932 4012
rect 439100 3754 439128 4012
rect 440204 3754 440232 4012
rect 435604 3726 435680 3754
rect 436708 3726 436784 3754
rect 437904 3726 437980 3754
rect 439100 3726 439176 3754
rect 433260 1358 433288 3726
rect 433248 1352 433300 1358
rect 433248 1294 433300 1300
rect 433248 1148 433300 1154
rect 433248 1090 433300 1096
rect 432144 1012 432196 1018
rect 432144 954 432196 960
rect 433260 480 433288 1090
rect 434364 814 434392 3726
rect 435652 1290 435680 3726
rect 435640 1284 435692 1290
rect 435640 1226 435692 1232
rect 436756 1154 436784 3726
rect 437848 1352 437900 1358
rect 437848 1294 437900 1300
rect 436744 1148 436796 1154
rect 436744 1090 436796 1096
rect 436744 1012 436796 1018
rect 436744 954 436796 960
rect 434444 876 434496 882
rect 434444 818 434496 824
rect 434352 808 434404 814
rect 434352 750 434404 756
rect 434456 480 434484 818
rect 436756 480 436784 954
rect 437860 762 437888 1294
rect 437952 950 437980 3726
rect 439148 1086 439176 3726
rect 440160 3726 440232 3754
rect 441400 3754 441428 4012
rect 442596 3754 442624 4012
rect 443700 3754 443728 4012
rect 444896 3754 444924 4012
rect 446000 3754 446028 4012
rect 447196 3754 447224 4012
rect 448392 3754 448420 4012
rect 449496 3754 449524 4012
rect 450692 3754 450720 4012
rect 451796 3754 451824 4012
rect 452992 3754 453020 4012
rect 454188 3754 454216 4012
rect 455292 3754 455320 4012
rect 456488 3754 456516 4012
rect 457592 3754 457620 4012
rect 458788 3754 458816 4012
rect 459984 3754 460012 4012
rect 461088 3754 461116 4012
rect 462284 3754 462312 4012
rect 441400 3726 441476 3754
rect 442596 3726 442672 3754
rect 443700 3726 443776 3754
rect 444896 3726 444972 3754
rect 446000 3726 446076 3754
rect 447196 3726 447272 3754
rect 448392 3726 448468 3754
rect 449496 3726 449572 3754
rect 450692 3726 450768 3754
rect 451796 3726 451872 3754
rect 452992 3726 453068 3754
rect 454188 3726 454264 3754
rect 455292 3726 455368 3754
rect 456488 3726 456564 3754
rect 457592 3726 457668 3754
rect 458788 3726 458864 3754
rect 459984 3726 460060 3754
rect 461088 3726 461164 3754
rect 440160 2854 440188 3726
rect 440148 2848 440200 2854
rect 440148 2790 440200 2796
rect 439964 1284 440016 1290
rect 439964 1226 440016 1232
rect 439136 1080 439188 1086
rect 439136 1022 439188 1028
rect 437940 944 437992 950
rect 437940 886 437992 892
rect 439136 808 439188 814
rect 437860 734 437980 762
rect 439136 750 439188 756
rect 437952 480 437980 734
rect 439148 480 439176 750
rect 432022 354 432134 480
rect 431880 326 432134 354
rect 431040 128 431092 134
rect 431040 70 431092 76
rect 432022 -960 432134 326
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435180 128 435232 134
rect 435518 82 435630 480
rect 435232 76 435630 82
rect 435180 70 435630 76
rect 435192 54 435630 70
rect 435518 -960 435630 54
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 439976 354 440004 1226
rect 441448 1222 441476 3726
rect 442644 1358 442672 3726
rect 442632 1352 442684 1358
rect 442632 1294 442684 1300
rect 441436 1216 441488 1222
rect 441436 1158 441488 1164
rect 441528 1148 441580 1154
rect 441528 1090 441580 1096
rect 441540 480 441568 1090
rect 442632 944 442684 950
rect 442632 886 442684 892
rect 442644 480 442672 886
rect 443748 882 443776 3726
rect 444944 1290 444972 3726
rect 445024 2848 445076 2854
rect 445024 2790 445076 2796
rect 444932 1284 444984 1290
rect 444932 1226 444984 1232
rect 443828 1080 443880 1086
rect 443828 1022 443880 1028
rect 443736 876 443788 882
rect 443736 818 443788 824
rect 443840 480 443868 1022
rect 445036 480 445064 2790
rect 446048 1222 446076 3726
rect 445852 1216 445904 1222
rect 445852 1158 445904 1164
rect 446036 1216 446088 1222
rect 446036 1158 446088 1164
rect 440302 354 440414 480
rect 439976 326 440414 354
rect 440302 -960 440414 326
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445864 354 445892 1158
rect 447244 1086 447272 3726
rect 448440 1358 448468 3726
rect 449544 2854 449572 3726
rect 449532 2848 449584 2854
rect 449532 2790 449584 2796
rect 447416 1352 447468 1358
rect 447416 1294 447468 1300
rect 448428 1352 448480 1358
rect 448428 1294 448480 1300
rect 447232 1080 447284 1086
rect 447232 1022 447284 1028
rect 447428 480 447456 1294
rect 450740 1290 450768 3726
rect 449808 1284 449860 1290
rect 449808 1226 449860 1232
rect 450728 1284 450780 1290
rect 450728 1226 450780 1232
rect 448244 876 448296 882
rect 448244 818 448296 824
rect 446190 354 446302 480
rect 445864 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448256 354 448284 818
rect 449820 480 449848 1226
rect 450912 1216 450964 1222
rect 450912 1158 450964 1164
rect 450924 480 450952 1158
rect 451844 882 451872 3726
rect 452108 1080 452160 1086
rect 452108 1022 452160 1028
rect 451832 876 451884 882
rect 451832 818 451884 824
rect 452120 480 452148 1022
rect 453040 1018 453068 3726
rect 453304 1352 453356 1358
rect 453304 1294 453356 1300
rect 453028 1012 453080 1018
rect 453028 954 453080 960
rect 453316 480 453344 1294
rect 454236 1154 454264 3726
rect 454500 2848 454552 2854
rect 454500 2790 454552 2796
rect 454224 1148 454276 1154
rect 454224 1090 454276 1096
rect 454512 480 454540 2790
rect 455340 1086 455368 3726
rect 456536 1290 456564 3726
rect 455696 1284 455748 1290
rect 455696 1226 455748 1232
rect 456524 1284 456576 1290
rect 456524 1226 456576 1232
rect 455328 1080 455380 1086
rect 455328 1022 455380 1028
rect 455708 480 455736 1226
rect 457640 1222 457668 3726
rect 458836 1358 458864 3726
rect 458824 1352 458876 1358
rect 458824 1294 458876 1300
rect 457628 1216 457680 1222
rect 457628 1158 457680 1164
rect 459192 1148 459244 1154
rect 459192 1090 459244 1096
rect 458088 1012 458140 1018
rect 458088 954 458140 960
rect 456524 876 456576 882
rect 456524 818 456576 824
rect 448582 354 448694 480
rect 448256 326 448694 354
rect 448582 -960 448694 326
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456536 354 456564 818
rect 458100 480 458128 954
rect 459204 480 459232 1090
rect 456862 354 456974 480
rect 456536 326 456974 354
rect 456862 -960 456974 326
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460032 134 460060 3726
rect 461136 1154 461164 3726
rect 462240 3726 462312 3754
rect 463388 3754 463416 4012
rect 464584 3754 464612 4012
rect 465780 3754 465808 4012
rect 466884 3754 466912 4012
rect 468080 3754 468108 4012
rect 469276 3754 469304 4012
rect 470380 3754 470408 4012
rect 471576 3754 471604 4012
rect 472680 3754 472708 4012
rect 473876 3754 473904 4012
rect 475072 3754 475100 4012
rect 476176 3754 476204 4012
rect 477372 3754 477400 4012
rect 478476 3754 478504 4012
rect 479672 3754 479700 4012
rect 480868 3754 480896 4012
rect 481972 3754 482000 4012
rect 483168 3754 483196 4012
rect 484272 3754 484300 4012
rect 485468 3754 485496 4012
rect 486664 3754 486692 4012
rect 487768 3754 487796 4012
rect 488964 3754 488992 4012
rect 490068 3754 490096 4012
rect 491264 3754 491292 4012
rect 463388 3726 463464 3754
rect 464584 3726 464660 3754
rect 465780 3726 465856 3754
rect 466884 3726 466960 3754
rect 468080 3726 468156 3754
rect 469276 3726 469352 3754
rect 470380 3726 470456 3754
rect 471576 3726 471652 3754
rect 472680 3726 472756 3754
rect 473876 3726 473952 3754
rect 475072 3726 475148 3754
rect 476176 3726 476252 3754
rect 477372 3726 477448 3754
rect 478476 3726 478552 3754
rect 479672 3726 479748 3754
rect 480868 3726 480944 3754
rect 481972 3726 482048 3754
rect 483168 3726 483244 3754
rect 484272 3726 484348 3754
rect 485468 3726 485544 3754
rect 486664 3726 486740 3754
rect 487768 3726 487844 3754
rect 488964 3726 489040 3754
rect 490068 3726 490144 3754
rect 462240 1290 462268 3726
rect 461584 1284 461636 1290
rect 461584 1226 461636 1232
rect 462228 1284 462280 1290
rect 462228 1226 462280 1232
rect 461124 1148 461176 1154
rect 461124 1090 461176 1096
rect 460112 1080 460164 1086
rect 460112 1022 460164 1028
rect 460124 354 460152 1022
rect 461596 480 461624 1226
rect 462412 1216 462464 1222
rect 462412 1158 462464 1164
rect 460358 354 460470 480
rect 460124 326 460470 354
rect 460020 128 460072 134
rect 460020 70 460072 76
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462424 354 462452 1158
rect 463436 882 463464 3726
rect 463976 1352 464028 1358
rect 463976 1294 464028 1300
rect 463424 876 463476 882
rect 463424 818 463476 824
rect 463988 480 464016 1294
rect 464632 1018 464660 3726
rect 465828 1222 465856 3726
rect 465816 1216 465868 1222
rect 465816 1158 465868 1164
rect 466276 1148 466328 1154
rect 466276 1090 466328 1096
rect 464620 1012 464672 1018
rect 464620 954 464672 960
rect 466288 480 466316 1090
rect 466932 1086 466960 3726
rect 468128 1358 468156 3726
rect 468116 1352 468168 1358
rect 468116 1294 468168 1300
rect 467472 1284 467524 1290
rect 467472 1226 467524 1232
rect 466920 1080 466972 1086
rect 466920 1022 466972 1028
rect 467484 480 467512 1226
rect 468668 876 468720 882
rect 468668 818 468720 824
rect 468680 480 468708 818
rect 462750 354 462862 480
rect 462424 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 464988 128 465040 134
rect 465142 82 465254 480
rect 465040 76 465254 82
rect 464988 70 465254 76
rect 465000 54 465254 70
rect 465142 -960 465254 54
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469324 270 469352 3726
rect 469864 1012 469916 1018
rect 469864 954 469916 960
rect 469876 480 469904 954
rect 469312 264 469364 270
rect 469312 206 469364 212
rect 469834 -960 469946 480
rect 470428 134 470456 3726
rect 471624 1290 471652 3726
rect 471612 1284 471664 1290
rect 471612 1226 471664 1232
rect 470692 1216 470744 1222
rect 470692 1158 470744 1164
rect 470704 354 470732 1158
rect 472728 1154 472756 3726
rect 473084 1352 473136 1358
rect 473084 1294 473136 1300
rect 472716 1148 472768 1154
rect 472716 1090 472768 1096
rect 472256 1080 472308 1086
rect 472256 1022 472308 1028
rect 472268 480 472296 1022
rect 471030 354 471142 480
rect 470704 326 471142 354
rect 470416 128 470468 134
rect 470416 70 470468 76
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473096 354 473124 1294
rect 473924 1018 473952 3726
rect 475120 1222 475148 3726
rect 475108 1216 475160 1222
rect 475108 1158 475160 1164
rect 473912 1012 473964 1018
rect 473912 954 473964 960
rect 476224 882 476252 3726
rect 476580 1284 476632 1290
rect 476580 1226 476632 1232
rect 476212 876 476264 882
rect 476212 818 476264 824
rect 473422 354 473534 480
rect 473096 326 473534 354
rect 473422 -960 473534 326
rect 474188 264 474240 270
rect 474526 218 474638 480
rect 474240 212 474638 218
rect 474188 206 474638 212
rect 474200 190 474638 206
rect 474526 -960 474638 190
rect 475722 82 475834 480
rect 476592 354 476620 1226
rect 477420 1086 477448 3726
rect 478524 2854 478552 3726
rect 478512 2848 478564 2854
rect 478512 2790 478564 2796
rect 479720 1290 479748 3726
rect 480916 1358 480944 3726
rect 480904 1352 480956 1358
rect 480904 1294 480956 1300
rect 479708 1284 479760 1290
rect 479708 1226 479760 1232
rect 482020 1222 482048 3726
rect 480536 1216 480588 1222
rect 480536 1158 480588 1164
rect 482008 1216 482060 1222
rect 482008 1158 482060 1164
rect 478144 1148 478196 1154
rect 478144 1090 478196 1096
rect 477408 1080 477460 1086
rect 477408 1022 477460 1028
rect 478156 480 478184 1090
rect 479340 1012 479392 1018
rect 479340 954 479392 960
rect 479352 480 479380 954
rect 480548 480 480576 1158
rect 482468 1080 482520 1086
rect 482468 1022 482520 1028
rect 481364 876 481416 882
rect 481364 818 481416 824
rect 476918 354 477030 480
rect 476592 326 477030 354
rect 475936 128 475988 134
rect 475722 76 475936 82
rect 475722 70 475988 76
rect 475722 54 475976 70
rect 475722 -960 475834 54
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481376 354 481404 818
rect 481702 354 481814 480
rect 481376 326 481814 354
rect 482480 354 482508 1022
rect 483216 950 483244 3726
rect 484032 2848 484084 2854
rect 484032 2790 484084 2796
rect 483204 944 483256 950
rect 483204 886 483256 892
rect 484044 480 484072 2790
rect 484320 1018 484348 3726
rect 484860 1284 484912 1290
rect 484860 1226 484912 1232
rect 484308 1012 484360 1018
rect 484308 954 484360 960
rect 482806 354 482918 480
rect 482480 326 482918 354
rect 481702 -960 481814 326
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484872 354 484900 1226
rect 485516 1086 485544 3726
rect 486424 1352 486476 1358
rect 486424 1294 486476 1300
rect 485504 1080 485556 1086
rect 485504 1022 485556 1028
rect 486436 480 486464 1294
rect 486712 1154 486740 3726
rect 487816 1358 487844 3726
rect 487804 1352 487856 1358
rect 487804 1294 487856 1300
rect 489012 1290 489040 3726
rect 489000 1284 489052 1290
rect 489000 1226 489052 1232
rect 487252 1216 487304 1222
rect 487252 1158 487304 1164
rect 486700 1148 486752 1154
rect 486700 1090 486752 1096
rect 485198 354 485310 480
rect 484872 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487264 354 487292 1158
rect 490116 1018 490144 3726
rect 491220 3726 491292 3754
rect 492460 3754 492488 4012
rect 493564 3754 493592 4012
rect 494760 3754 494788 4012
rect 495956 3754 495984 4012
rect 497060 3754 497088 4012
rect 498256 3754 498284 4012
rect 499360 3754 499388 4012
rect 500556 3754 500584 4012
rect 501752 3754 501780 4012
rect 492460 3726 492536 3754
rect 493564 3726 493640 3754
rect 494760 3726 494836 3754
rect 495956 3726 496032 3754
rect 497060 3726 497136 3754
rect 498256 3726 498332 3754
rect 490748 1080 490800 1086
rect 490748 1022 490800 1028
rect 489920 1012 489972 1018
rect 489920 954 489972 960
rect 490104 1012 490156 1018
rect 490104 954 490156 960
rect 488816 944 488868 950
rect 488816 886 488868 892
rect 488828 480 488856 886
rect 489932 480 489960 954
rect 487590 354 487702 480
rect 487264 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 1022
rect 491220 950 491248 3726
rect 492508 1222 492536 3726
rect 493140 1352 493192 1358
rect 493140 1294 493192 1300
rect 492496 1216 492548 1222
rect 492496 1158 492548 1164
rect 492312 1148 492364 1154
rect 492312 1090 492364 1096
rect 491208 944 491260 950
rect 491208 886 491260 892
rect 492324 480 492352 1090
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493152 354 493180 1294
rect 493612 1154 493640 3726
rect 494704 1284 494756 1290
rect 494704 1226 494756 1232
rect 493600 1148 493652 1154
rect 493600 1090 493652 1096
rect 494716 480 494744 1226
rect 494808 1086 494836 3726
rect 494796 1080 494848 1086
rect 494796 1022 494848 1028
rect 496004 1018 496032 3726
rect 497108 1358 497136 3726
rect 497096 1352 497148 1358
rect 497096 1294 497148 1300
rect 498304 1290 498332 3726
rect 499224 3726 499388 3754
rect 500512 3726 500584 3754
rect 501708 3726 501780 3754
rect 502856 3754 502884 4012
rect 504052 3754 504080 4012
rect 505156 3754 505184 4012
rect 506352 3754 506380 4012
rect 507548 3754 507576 4012
rect 502856 3726 502932 3754
rect 504052 3726 504128 3754
rect 505156 3726 505232 3754
rect 498292 1284 498344 1290
rect 498292 1226 498344 1232
rect 498200 1216 498252 1222
rect 498200 1158 498252 1164
rect 495532 1012 495584 1018
rect 495532 954 495584 960
rect 495992 1012 496044 1018
rect 495992 954 496044 960
rect 493478 354 493590 480
rect 493152 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495544 354 495572 954
rect 497096 944 497148 950
rect 497096 886 497148 892
rect 497108 480 497136 886
rect 498212 480 498240 1158
rect 495870 354 495982 480
rect 495544 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499224 66 499252 3726
rect 500512 1154 500540 3726
rect 499396 1148 499448 1154
rect 499396 1090 499448 1096
rect 500500 1148 500552 1154
rect 500500 1090 500552 1096
rect 499408 480 499436 1090
rect 501708 1086 501736 3726
rect 500592 1080 500644 1086
rect 500592 1022 500644 1028
rect 501696 1080 501748 1086
rect 501696 1022 501748 1028
rect 500604 480 500632 1022
rect 502904 1018 502932 3726
rect 504100 1358 504128 3726
rect 502984 1352 503036 1358
rect 502984 1294 503036 1300
rect 504088 1352 504140 1358
rect 504088 1294 504140 1300
rect 501788 1012 501840 1018
rect 501788 954 501840 960
rect 502892 1012 502944 1018
rect 502892 954 502944 960
rect 501800 480 501828 954
rect 502996 480 503024 1294
rect 503812 1284 503864 1290
rect 503812 1226 503864 1232
rect 499212 60 499264 66
rect 499212 2 499264 8
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503824 354 503852 1226
rect 505204 1222 505232 3726
rect 506308 3726 506380 3754
rect 507504 3726 507576 3754
rect 508652 3754 508680 4012
rect 509848 3754 509876 4012
rect 510952 3754 510980 4012
rect 512148 3754 512176 4012
rect 513344 3754 513372 4012
rect 508652 3726 508728 3754
rect 509848 3726 509924 3754
rect 510952 3726 511028 3754
rect 512148 3726 512224 3754
rect 505192 1216 505244 1222
rect 505192 1158 505244 1164
rect 504150 354 504262 480
rect 503824 326 504262 354
rect 504150 -960 504262 326
rect 505346 82 505458 480
rect 505346 66 505600 82
rect 506308 66 506336 3726
rect 506480 1148 506532 1154
rect 506480 1090 506532 1096
rect 506492 480 506520 1090
rect 507308 1080 507360 1086
rect 507308 1022 507360 1028
rect 505346 60 505612 66
rect 505346 54 505560 60
rect 505346 -960 505458 54
rect 505560 2 505612 8
rect 506296 60 506348 66
rect 506296 2 506348 8
rect 506450 -960 506562 480
rect 507320 354 507348 1022
rect 507504 474 507532 3726
rect 507492 468 507544 474
rect 507492 410 507544 416
rect 507646 354 507758 480
rect 507320 326 507758 354
rect 507646 -960 507758 326
rect 508700 270 508728 3726
rect 509896 1358 509924 3726
rect 509700 1352 509752 1358
rect 509700 1294 509752 1300
rect 509884 1352 509936 1358
rect 509884 1294 509936 1300
rect 508872 1012 508924 1018
rect 508872 954 508924 960
rect 508884 480 508912 954
rect 508688 264 508740 270
rect 508688 206 508740 212
rect 508842 -960 508954 480
rect 509712 354 509740 1294
rect 511000 1290 511028 3726
rect 510988 1284 511040 1290
rect 510988 1226 511040 1232
rect 511264 1216 511316 1222
rect 511264 1158 511316 1164
rect 511276 480 511304 1158
rect 512196 1154 512224 3726
rect 513300 3726 513372 3754
rect 514448 3754 514476 4012
rect 515644 3754 515672 4012
rect 516748 3754 516776 4012
rect 517944 3754 517972 4012
rect 519140 3754 519168 4012
rect 520244 3754 520272 4012
rect 514448 3726 514524 3754
rect 515644 3726 515720 3754
rect 516748 3726 516824 3754
rect 517944 3726 518020 3754
rect 519140 3726 519216 3754
rect 513300 1222 513328 3726
rect 513288 1216 513340 1222
rect 513288 1158 513340 1164
rect 512184 1148 512236 1154
rect 512184 1090 512236 1096
rect 514496 1086 514524 3726
rect 514484 1080 514536 1086
rect 514484 1022 514536 1028
rect 510038 354 510150 480
rect 509712 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512430 82 512542 480
rect 513380 468 513432 474
rect 513380 410 513432 416
rect 513392 354 513420 410
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512104 66 512542 82
rect 512092 60 512542 66
rect 512144 54 512542 60
rect 512092 2 512144 8
rect 512430 -960 512542 54
rect 513534 -960 513646 326
rect 514730 218 514842 480
rect 514944 264 514996 270
rect 514730 212 514944 218
rect 514730 206 514996 212
rect 514730 190 514984 206
rect 514730 -960 514842 190
rect 515692 134 515720 3726
rect 515772 1352 515824 1358
rect 515772 1294 515824 1300
rect 515784 354 515812 1294
rect 515926 354 516038 480
rect 515784 326 516038 354
rect 515680 128 515732 134
rect 515680 70 515732 76
rect 515926 -960 516038 326
rect 516796 66 516824 3726
rect 517992 1290 518020 3726
rect 519188 1358 519216 3726
rect 520200 3726 520272 3754
rect 521440 3754 521468 4012
rect 522636 3754 522664 4012
rect 523740 3754 523768 4012
rect 524936 3754 524964 4012
rect 526040 3754 526068 4012
rect 527236 3754 527264 4012
rect 528432 3754 528460 4012
rect 529536 3754 529564 4012
rect 530732 3754 530760 4012
rect 531836 3754 531864 4012
rect 533032 3754 533060 4012
rect 534228 3754 534256 4012
rect 535332 3754 535360 4012
rect 536528 3754 536556 4012
rect 537632 3754 537660 4012
rect 538828 3754 538856 4012
rect 540024 3754 540052 4012
rect 541128 3754 541156 4012
rect 542324 3754 542352 4012
rect 521440 3726 521516 3754
rect 522636 3726 522712 3754
rect 523740 3726 523816 3754
rect 524936 3726 525012 3754
rect 526040 3726 526116 3754
rect 527236 3726 527312 3754
rect 528432 3726 528508 3754
rect 529536 3726 529612 3754
rect 530732 3726 530808 3754
rect 531836 3726 531912 3754
rect 533032 3726 533108 3754
rect 534228 3726 534304 3754
rect 535332 3726 535408 3754
rect 536528 3726 536604 3754
rect 537632 3726 537708 3754
rect 538828 3726 538904 3754
rect 540024 3726 540100 3754
rect 541128 3726 541204 3754
rect 519176 1352 519228 1358
rect 519176 1294 519228 1300
rect 517152 1284 517204 1290
rect 517152 1226 517204 1232
rect 517980 1284 518032 1290
rect 517980 1226 518032 1232
rect 517164 480 517192 1226
rect 519544 1216 519596 1222
rect 519544 1158 519596 1164
rect 517980 1148 518032 1154
rect 517980 1090 518032 1096
rect 516784 60 516836 66
rect 516784 2 516836 8
rect 517122 -960 517234 480
rect 517992 354 518020 1090
rect 519556 480 519584 1158
rect 520200 1018 520228 3726
rect 521488 1086 521516 3726
rect 522684 1222 522712 3726
rect 522672 1216 522724 1222
rect 522672 1158 522724 1164
rect 523788 1154 523816 3726
rect 523868 1284 523920 1290
rect 523868 1226 523920 1232
rect 523776 1148 523828 1154
rect 523776 1090 523828 1096
rect 520740 1080 520792 1086
rect 520740 1022 520792 1028
rect 521476 1080 521528 1086
rect 521476 1022 521528 1028
rect 520188 1012 520240 1018
rect 520188 954 520240 960
rect 520752 480 520780 1022
rect 518318 354 518430 480
rect 517992 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521660 128 521712 134
rect 521814 82 521926 480
rect 521712 76 521926 82
rect 521660 70 521926 76
rect 521672 54 521926 70
rect 521814 -960 521926 54
rect 523010 82 523122 480
rect 523880 354 523908 1226
rect 524206 354 524318 480
rect 523880 326 524318 354
rect 523010 66 523264 82
rect 523010 60 523276 66
rect 523010 54 523224 60
rect 523010 -960 523122 54
rect 523224 2 523276 8
rect 524206 -960 524318 326
rect 524984 134 525012 3726
rect 526088 1358 526116 3726
rect 525432 1352 525484 1358
rect 525432 1294 525484 1300
rect 526076 1352 526128 1358
rect 526076 1294 526128 1300
rect 525444 480 525472 1294
rect 527284 1290 527312 3726
rect 527272 1284 527324 1290
rect 527272 1226 527324 1232
rect 527824 1080 527876 1086
rect 527824 1022 527876 1028
rect 526628 1012 526680 1018
rect 526628 954 526680 960
rect 526640 480 526668 954
rect 527836 480 527864 1022
rect 524972 128 525024 134
rect 524972 70 525024 76
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528480 270 528508 3726
rect 529020 1216 529072 1222
rect 529020 1158 529072 1164
rect 529032 480 529060 1158
rect 529584 1086 529612 3726
rect 530780 1154 530808 3726
rect 531884 1222 531912 3726
rect 532148 1352 532200 1358
rect 532148 1294 532200 1300
rect 531872 1216 531924 1222
rect 531872 1158 531924 1164
rect 530124 1148 530176 1154
rect 530124 1090 530176 1096
rect 530768 1148 530820 1154
rect 530768 1090 530820 1096
rect 529572 1080 529624 1086
rect 529572 1022 529624 1028
rect 530136 480 530164 1090
rect 528468 264 528520 270
rect 528468 206 528520 212
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 82 531402 480
rect 532160 354 532188 1294
rect 533080 1018 533108 3726
rect 534276 1358 534304 3726
rect 534264 1352 534316 1358
rect 534264 1294 534316 1300
rect 533712 1284 533764 1290
rect 533712 1226 533764 1232
rect 533068 1012 533120 1018
rect 533068 954 533120 960
rect 533724 480 533752 1226
rect 532486 354 532598 480
rect 532160 326 532598 354
rect 531504 128 531556 134
rect 531290 76 531504 82
rect 531290 70 531556 76
rect 531290 54 531544 70
rect 531290 -960 531402 54
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534540 264 534592 270
rect 534878 218 534990 480
rect 535380 406 535408 3726
rect 536104 1080 536156 1086
rect 536104 1022 536156 1028
rect 536116 480 536144 1022
rect 535368 400 535420 406
rect 535368 342 535420 348
rect 534592 212 534990 218
rect 534540 206 534990 212
rect 534552 190 534990 206
rect 534878 -960 534990 190
rect 536074 -960 536186 480
rect 536576 474 536604 3726
rect 537208 1148 537260 1154
rect 537208 1090 537260 1096
rect 537220 480 537248 1090
rect 536564 468 536616 474
rect 536564 410 536616 416
rect 537178 -960 537290 480
rect 537680 338 537708 3726
rect 538404 1216 538456 1222
rect 538404 1158 538456 1164
rect 538416 480 538444 1158
rect 538876 1154 538904 3726
rect 540072 1222 540100 3726
rect 540428 1352 540480 1358
rect 540428 1294 540480 1300
rect 540060 1216 540112 1222
rect 540060 1158 540112 1164
rect 538864 1148 538916 1154
rect 538864 1090 538916 1096
rect 539600 1012 539652 1018
rect 539600 954 539652 960
rect 539612 480 539640 954
rect 537668 332 537720 338
rect 537668 274 537720 280
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540440 354 540468 1294
rect 541176 746 541204 3726
rect 542280 3726 542352 3754
rect 543428 3754 543456 4012
rect 544624 3754 544652 4012
rect 545820 3754 545848 4012
rect 546924 3754 546952 4012
rect 548120 3754 548148 4012
rect 549316 3754 549344 4012
rect 550420 3754 550448 4012
rect 551616 3754 551644 4012
rect 552720 3754 552748 4012
rect 553916 3754 553944 4012
rect 555112 3754 555140 4012
rect 556216 3754 556244 4012
rect 557412 3754 557440 4012
rect 558516 3754 558544 4012
rect 559712 3754 559740 4012
rect 543428 3726 543504 3754
rect 544624 3726 544700 3754
rect 545820 3726 545896 3754
rect 546924 3726 547000 3754
rect 548120 3726 548196 3754
rect 549316 3726 549392 3754
rect 550420 3726 550496 3754
rect 551616 3726 551692 3754
rect 552720 3726 552796 3754
rect 553916 3726 553992 3754
rect 555112 3726 555188 3754
rect 556216 3726 556292 3754
rect 557412 3726 557488 3754
rect 542280 1358 542308 3726
rect 542268 1352 542320 1358
rect 542268 1294 542320 1300
rect 543476 1290 543504 3726
rect 543464 1284 543516 1290
rect 543464 1226 543516 1232
rect 541164 740 541216 746
rect 541164 682 541216 688
rect 540766 354 540878 480
rect 540440 326 540878 354
rect 540766 -960 540878 326
rect 541962 354 542074 480
rect 542820 468 542872 474
rect 542820 410 542872 416
rect 542176 400 542228 406
rect 541962 348 542176 354
rect 541962 342 542228 348
rect 542832 354 542860 410
rect 543158 354 543270 480
rect 541962 326 542216 342
rect 542832 326 543270 354
rect 541962 -960 542074 326
rect 543158 -960 543270 326
rect 544354 354 544466 480
rect 544672 474 544700 3726
rect 545488 1148 545540 1154
rect 545488 1090 545540 1096
rect 545500 480 545528 1090
rect 544660 468 544712 474
rect 544660 410 544712 416
rect 544354 338 544608 354
rect 544354 332 544620 338
rect 544354 326 544568 332
rect 544354 -960 544466 326
rect 544568 274 544620 280
rect 545458 -960 545570 480
rect 545868 338 545896 3726
rect 546684 1216 546736 1222
rect 546684 1158 546736 1164
rect 546696 480 546724 1158
rect 545856 332 545908 338
rect 545856 274 545908 280
rect 546654 -960 546766 480
rect 546972 406 547000 3726
rect 548168 1222 548196 3726
rect 549076 1352 549128 1358
rect 549076 1294 549128 1300
rect 548156 1216 548208 1222
rect 548156 1158 548208 1164
rect 547880 740 547932 746
rect 547880 682 547932 688
rect 547892 480 547920 682
rect 549088 480 549116 1294
rect 549364 1086 549392 3726
rect 550468 1290 550496 3726
rect 551664 1358 551692 3726
rect 551652 1352 551704 1358
rect 551652 1294 551704 1300
rect 550272 1284 550324 1290
rect 550272 1226 550324 1232
rect 550456 1284 550508 1290
rect 550456 1226 550508 1232
rect 549352 1080 549404 1086
rect 549352 1022 549404 1028
rect 550284 480 550312 1226
rect 552768 1154 552796 3726
rect 552756 1148 552808 1154
rect 552756 1090 552808 1096
rect 553964 678 553992 3726
rect 554964 1216 555016 1222
rect 554964 1158 555016 1164
rect 553952 672 554004 678
rect 552400 598 552704 626
rect 553952 614 554004 620
rect 546960 400 547012 406
rect 546960 342 547012 348
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551100 468 551152 474
rect 551100 410 551152 416
rect 551112 354 551140 410
rect 551438 354 551550 480
rect 551112 326 551550 354
rect 552400 338 552428 598
rect 552676 480 552704 598
rect 554976 480 555004 1158
rect 551438 -960 551550 326
rect 552388 332 552440 338
rect 552388 274 552440 280
rect 552634 -960 552746 480
rect 553738 354 553850 480
rect 553952 400 554004 406
rect 553738 348 553952 354
rect 553738 342 554004 348
rect 553738 326 553992 342
rect 553738 -960 553850 326
rect 554934 -960 555046 480
rect 555160 134 555188 3726
rect 556160 1080 556212 1086
rect 556160 1022 556212 1028
rect 556172 480 556200 1022
rect 556264 610 556292 3726
rect 557356 1284 557408 1290
rect 557356 1226 557408 1232
rect 556252 604 556304 610
rect 556252 546 556304 552
rect 557368 480 557396 1226
rect 557460 626 557488 3726
rect 558472 3726 558544 3754
rect 559668 3726 559740 3754
rect 560908 3754 560936 4012
rect 562012 3754 562040 4012
rect 563208 3754 563236 4012
rect 564312 3754 564340 4012
rect 565508 3754 565536 4012
rect 566704 3754 566732 4012
rect 560908 3726 560984 3754
rect 562012 3726 562088 3754
rect 558472 1222 558500 3726
rect 558552 1352 558604 1358
rect 558552 1294 558604 1300
rect 558460 1216 558512 1222
rect 558460 1158 558512 1164
rect 557540 740 557592 746
rect 557540 682 557592 688
rect 557552 626 557580 682
rect 557460 598 557580 626
rect 558564 480 558592 1294
rect 559668 1086 559696 3726
rect 560956 1358 560984 3726
rect 560944 1352 560996 1358
rect 560944 1294 560996 1300
rect 562060 1290 562088 3726
rect 563164 3726 563236 3754
rect 564268 3726 564340 3754
rect 565464 3726 565536 3754
rect 566660 3726 566732 3754
rect 567808 3754 567836 4012
rect 569004 3754 569032 4012
rect 570108 3754 570136 4012
rect 571304 3754 571332 4012
rect 567808 3726 567884 3754
rect 569004 3726 569080 3754
rect 570108 3726 570184 3754
rect 562048 1284 562100 1290
rect 562048 1226 562100 1232
rect 559748 1148 559800 1154
rect 559748 1090 559800 1096
rect 559656 1080 559708 1086
rect 559656 1022 559708 1028
rect 559760 480 559788 1090
rect 563164 678 563192 3726
rect 563152 672 563204 678
rect 563152 614 563204 620
rect 560852 604 560904 610
rect 560852 546 560904 552
rect 563244 604 563296 610
rect 563244 546 563296 552
rect 560864 480 560892 546
rect 563256 480 563284 546
rect 555148 128 555200 134
rect 555148 70 555200 76
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 82 562130 480
rect 562232 128 562284 134
rect 562018 76 562232 82
rect 562018 70 562284 76
rect 562018 54 562272 70
rect 562018 -960 562130 54
rect 563214 -960 563326 480
rect 564268 202 564296 3726
rect 564440 740 564492 746
rect 564440 682 564492 688
rect 564452 480 564480 682
rect 564256 196 564308 202
rect 564256 138 564308 144
rect 564410 -960 564522 480
rect 565464 134 565492 3726
rect 565636 1216 565688 1222
rect 565636 1158 565688 1164
rect 565648 480 565676 1158
rect 565452 128 565504 134
rect 565452 70 565504 76
rect 565606 -960 565718 480
rect 566660 474 566688 3726
rect 567856 1154 567884 3726
rect 568028 1352 568080 1358
rect 568028 1294 568080 1300
rect 567844 1148 567896 1154
rect 567844 1090 567896 1096
rect 566832 1080 566884 1086
rect 566832 1022 566884 1028
rect 566844 480 566872 1022
rect 568040 480 568068 1294
rect 569052 1222 569080 3726
rect 570156 1290 570184 3726
rect 571260 3726 571332 3754
rect 572500 3754 572528 4012
rect 573604 3754 573632 4012
rect 574800 3754 574828 4012
rect 575918 3998 576164 4026
rect 572500 3726 572576 3754
rect 573604 3726 573680 3754
rect 574800 3726 574876 3754
rect 571260 1358 571288 3726
rect 571248 1352 571300 1358
rect 571248 1294 571300 1300
rect 569132 1284 569184 1290
rect 569132 1226 569184 1232
rect 570144 1284 570196 1290
rect 570144 1226 570196 1232
rect 569040 1216 569092 1222
rect 569040 1158 569092 1164
rect 569144 480 569172 1226
rect 570328 672 570380 678
rect 570328 614 570380 620
rect 570340 480 570368 614
rect 566648 468 566700 474
rect 566648 410 566700 416
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 218 571606 480
rect 571352 202 571606 218
rect 571340 196 571606 202
rect 571392 190 571606 196
rect 571340 138 571392 144
rect 571494 -960 571606 190
rect 572548 66 572576 3726
rect 572690 82 572802 480
rect 573652 338 573680 3726
rect 573732 468 573784 474
rect 573732 410 573784 416
rect 573744 354 573772 410
rect 573886 354 573998 480
rect 573640 332 573692 338
rect 573744 326 573998 354
rect 573640 274 573692 280
rect 572904 128 572956 134
rect 572690 76 572904 82
rect 572690 70 572956 76
rect 572536 60 572588 66
rect 572536 2 572588 8
rect 572690 54 572944 70
rect 572690 -960 572802 54
rect 573886 -960 573998 326
rect 574848 202 574876 3726
rect 575112 1148 575164 1154
rect 575112 1090 575164 1096
rect 575124 480 575152 1090
rect 574836 196 574888 202
rect 574836 138 574888 144
rect 575082 -960 575194 480
rect 576136 134 576164 3998
rect 578608 1352 578660 1358
rect 578608 1294 578660 1300
rect 577412 1284 577464 1290
rect 577412 1226 577464 1232
rect 576308 1216 576360 1222
rect 576308 1158 576360 1164
rect 576320 480 576348 1158
rect 577424 480 577452 1226
rect 578620 480 578648 1294
rect 576124 128 576176 134
rect 576124 70 576176 76
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 82 579886 480
rect 579632 66 579886 82
rect 579620 60 579886 66
rect 579672 54 579886 60
rect 579620 2 579672 8
rect 579774 -960 579886 54
rect 580970 354 581082 480
rect 580970 338 581224 354
rect 580970 332 581236 338
rect 580970 326 581184 332
rect 580970 -960 581082 326
rect 581184 274 581236 280
rect 582166 218 582278 480
rect 581840 202 582278 218
rect 581828 196 582278 202
rect 581880 190 582278 196
rect 581828 138 581880 144
rect 582166 -960 582278 190
rect 583362 82 583474 480
rect 583576 128 583628 134
rect 583362 76 583576 82
rect 583362 70 583628 76
rect 583362 54 583616 70
rect 583362 -960 583474 54
<< via2 >>
rect 3514 697920 3570 697976
rect 576766 698128 576822 698184
rect 3514 697312 3570 697368
rect 580170 697176 580226 697232
rect 579526 684664 579582 684720
rect 579618 683848 579674 683904
rect 578330 644564 578386 644600
rect 578330 644544 578332 644564
rect 578332 644544 578384 644564
rect 578384 644544 578386 644564
rect 580906 644000 580962 644056
rect 3422 436600 3478 436656
rect 3422 435986 3478 436042
rect 3422 423544 3478 423600
rect 3422 422932 3478 422988
rect 3422 410488 3478 410544
rect 3422 409878 3478 409934
rect 3422 397432 3478 397488
rect 3422 396824 3478 396880
rect 3422 384376 3478 384432
rect 3422 383648 3478 383704
rect 3422 371320 3478 371376
rect 3422 370594 3478 370650
rect 3422 358400 3478 358456
rect 3422 357540 3478 357596
rect 579526 351872 579582 351928
rect 579526 351056 579582 351112
rect 3422 345344 3478 345400
rect 3422 344364 3478 344420
rect 579618 338544 579674 338600
rect 579526 337864 579582 337920
rect 3422 332288 3478 332344
rect 3422 331310 3478 331366
rect 580170 325216 580226 325272
rect 580170 324400 580226 324456
rect 3422 319232 3478 319288
rect 3422 318256 3478 318312
rect 579618 312024 579674 312080
rect 579526 311072 579582 311128
rect 3422 306176 3478 306232
rect 3422 305080 3478 305136
rect 579618 298696 579674 298752
rect 579526 297744 579582 297800
rect 3422 293120 3478 293176
rect 3422 292026 3478 292082
rect 580170 285368 580226 285424
rect 580170 284416 580226 284472
rect 3422 280064 3478 280120
rect 3422 278972 3478 279028
rect 579618 272176 579674 272232
rect 579526 271088 579582 271144
rect 3422 267144 3478 267200
rect 3422 265918 3478 265974
rect 580906 258848 580962 258904
rect 578882 257624 578938 257680
rect 3422 254088 3478 254144
rect 3422 252742 3478 252798
rect 580170 245520 580226 245576
rect 580170 244432 580226 244488
rect 3422 241032 3478 241088
rect 3422 239688 3478 239744
rect 579618 232328 579674 232384
rect 579526 231104 579582 231160
rect 3422 227976 3478 228032
rect 3422 226634 3478 226690
rect 579618 219000 579674 219056
rect 579526 217640 579582 217696
rect 3422 214920 3478 214976
rect 3422 213458 3478 213514
rect 579618 205672 579674 205728
rect 579526 204312 579582 204368
rect 3422 201864 3478 201920
rect 3422 200404 3478 200460
rect 579618 192480 579674 192536
rect 579526 190984 579582 191040
rect 3606 188808 3662 188864
rect 3606 187350 3662 187406
rect 579618 179152 579674 179208
rect 579526 177656 579582 177712
rect 3422 175888 3478 175944
rect 3422 174174 3478 174230
rect 579618 165824 579674 165880
rect 579526 164328 579582 164384
rect 2134 162832 2190 162888
rect 2134 161064 2190 161120
rect 580906 152632 580962 152688
rect 578514 151000 578570 151056
rect 3422 149776 3478 149832
rect 3422 148066 3478 148122
rect 579618 139304 579674 139360
rect 579526 137536 579582 137592
rect 2134 136720 2190 136776
rect 2134 134952 2190 135008
rect 579618 125976 579674 126032
rect 579526 124344 579582 124400
rect 3422 123664 3478 123720
rect 3422 121836 3478 121892
rect 579618 112784 579674 112840
rect 579526 110880 579582 110936
rect 2134 110608 2190 110664
rect 2134 108840 2190 108896
rect 579618 99456 579674 99512
rect 3422 97552 3478 97608
rect 579526 97552 579582 97608
rect 3422 95728 3478 95784
rect 579618 86128 579674 86184
rect 2134 84632 2190 84688
rect 579526 84224 579582 84280
rect 2134 82592 2190 82648
rect 579618 72936 579674 72992
rect 3422 71576 3478 71632
rect 579526 70896 579582 70952
rect 3422 69498 3478 69554
rect 579618 59608 579674 59664
rect 2134 58520 2190 58576
rect 579526 57568 579582 57624
rect 2134 56480 2190 56536
rect 579986 46280 580042 46336
rect 3422 45464 3478 45520
rect 578330 44240 578386 44296
rect 3422 43268 3478 43324
rect 579618 33088 579674 33144
rect 2134 32408 2190 32464
rect 579526 30912 579582 30968
rect 2134 30232 2190 30288
rect 579618 19760 579674 19816
rect 2042 19352 2098 19408
rect 579526 17584 579582 17640
rect 2042 17176 2098 17232
rect 579618 6568 579674 6624
rect 2778 6432 2834 6488
rect 2778 4120 2834 4176
rect 576766 4120 576822 4176
<< metal3 >>
rect 576761 698186 576827 698189
rect 575890 698184 576827 698186
rect 575890 698128 576766 698184
rect 576822 698128 576827 698184
rect 575890 698126 576827 698128
rect 3509 697978 3575 697981
rect 3509 697976 4048 697978
rect 3509 697920 3514 697976
rect 3570 697920 4048 697976
rect 575890 697948 575950 698126
rect 576761 698123 576827 698126
rect 3509 697918 4048 697920
rect 3509 697915 3575 697918
rect -960 697370 480 697460
rect 3509 697370 3575 697373
rect -960 697368 3575 697370
rect -960 697312 3514 697368
rect 3570 697312 3575 697368
rect -960 697310 3575 697312
rect -960 697220 480 697310
rect 3509 697307 3575 697310
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect 3374 684742 4048 684802
rect -960 684314 480 684404
rect 3374 684314 3434 684742
rect 579521 684722 579587 684725
rect 576350 684720 579587 684722
rect 576350 684680 579526 684720
rect 575920 684664 579526 684680
rect 579582 684664 579587 684720
rect 575920 684662 579587 684664
rect 575920 684620 576410 684662
rect 579521 684659 579587 684662
rect -960 684254 3434 684314
rect -960 684164 480 684254
rect 579613 683906 579679 683909
rect 583520 683906 584960 683996
rect 579613 683904 584960 683906
rect 579613 683848 579618 683904
rect 579674 683848 584960 683904
rect 579613 683846 584960 683848
rect 579613 683843 579679 683846
rect 583520 683756 584960 683846
rect 3374 671688 4048 671748
rect -960 671258 480 671348
rect 3374 671258 3434 671688
rect 576350 671382 583586 671394
rect 575920 671334 583586 671382
rect 575920 671322 576410 671334
rect -960 671198 3434 671258
rect -960 671108 480 671198
rect 583526 670850 583586 671334
rect 583342 670804 583586 670850
rect 583342 670790 584960 670804
rect 583342 670714 583402 670790
rect 583520 670714 584960 670790
rect 583342 670654 584960 670714
rect 583520 670564 584960 670654
rect 3374 658634 4048 658694
rect -960 658202 480 658292
rect 3374 658202 3434 658634
rect -960 658142 3434 658202
rect -960 658052 480 658142
rect 575920 657930 576410 657962
rect 575920 657902 583586 657930
rect 576350 657870 583586 657902
rect 583526 657522 583586 657870
rect 583342 657476 583586 657522
rect 583342 657462 584960 657476
rect 583342 657386 583402 657462
rect 583520 657386 584960 657462
rect 583342 657326 584960 657386
rect 583520 657236 584960 657326
rect 3374 645458 4048 645518
rect -960 645146 480 645236
rect 3374 645146 3434 645458
rect -960 645086 3434 645146
rect -960 644996 480 645086
rect 575920 644604 576410 644664
rect 576350 644602 576410 644604
rect 578325 644602 578391 644605
rect 576350 644600 578391 644602
rect 576350 644544 578330 644600
rect 578386 644544 578391 644600
rect 576350 644542 578391 644544
rect 578325 644539 578391 644542
rect 580901 644058 580967 644061
rect 583520 644058 584960 644148
rect 580901 644056 584960 644058
rect 580901 644000 580906 644056
rect 580962 644000 584960 644056
rect 580901 643998 584960 644000
rect 580901 643995 580967 643998
rect 583520 643908 584960 643998
rect 3374 632404 4048 632464
rect -960 632090 480 632180
rect 3374 632090 3434 632404
rect -960 632030 3434 632090
rect -960 631940 480 632030
rect 575920 631306 576410 631366
rect 576350 631274 576410 631306
rect 576350 631214 583586 631274
rect 583526 631002 583586 631214
rect 583342 630956 583586 631002
rect 583342 630942 584960 630956
rect 583342 630866 583402 630942
rect 583520 630866 584960 630942
rect 583342 630806 584960 630866
rect 583520 630716 584960 630806
rect 3374 619350 4048 619410
rect -960 619170 480 619260
rect 3374 619170 3434 619350
rect -960 619110 3434 619170
rect -960 619020 480 619110
rect 575920 617886 583586 617946
rect 583526 617674 583586 617886
rect 583342 617628 583586 617674
rect 583342 617614 584960 617628
rect 583342 617538 583402 617614
rect 583520 617538 584960 617614
rect 583342 617478 584960 617538
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3374 606174 4048 606234
rect 3374 606114 3434 606174
rect -960 606054 3434 606114
rect -960 605964 480 606054
rect 575920 604618 576410 604648
rect 575920 604588 576870 604618
rect 576350 604558 576870 604588
rect 576810 604482 576870 604558
rect 576810 604422 579722 604482
rect 579662 604210 579722 604422
rect 583520 604210 584960 604300
rect 579662 604150 584960 604210
rect 583520 604060 584960 604150
rect -960 593058 480 593148
rect 3374 593120 4048 593180
rect 3374 593058 3434 593120
rect -960 592998 3434 593058
rect -960 592908 480 592998
rect 575920 591290 576410 591350
rect 576350 591230 576870 591290
rect 576810 591018 576870 591230
rect 583520 591018 584960 591108
rect 576810 590958 584960 591018
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3374 580066 4048 580126
rect 3374 580002 3434 580066
rect -960 579942 3434 580002
rect -960 579852 480 579942
rect 575920 577870 576410 577930
rect 576350 577826 576410 577870
rect 576350 577766 576870 577826
rect 576810 577690 576870 577766
rect 583520 577690 584960 577780
rect 576810 577630 584960 577690
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3374 566946 4048 566950
rect -960 566890 4048 566946
rect -960 566886 3434 566890
rect -960 566796 480 566886
rect 575920 564572 576410 564632
rect 576350 564498 576410 564572
rect 576350 564438 579722 564498
rect 579662 564362 579722 564438
rect 583520 564362 584960 564452
rect 579662 564302 584960 564362
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3374 553890 4048 553896
rect -960 553836 4048 553890
rect -960 553830 3434 553836
rect -960 553740 480 553830
rect 575920 551170 576410 551212
rect 583520 551170 584960 551260
rect 575920 551152 584960 551170
rect 576350 551110 584960 551152
rect 583520 551020 584960 551110
rect -960 540834 480 540924
rect 3374 540834 4048 540842
rect -960 540782 4048 540834
rect -960 540774 3434 540782
rect -960 540684 480 540774
rect 575920 537854 576410 537914
rect 576350 537842 576410 537854
rect 583520 537842 584960 537932
rect 576350 537782 584960 537842
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect -960 527854 3434 527914
rect -960 527764 480 527854
rect 3374 527788 3434 527854
rect 3374 527728 4048 527788
rect 575920 524556 576410 524616
rect 576350 524514 576410 524556
rect 583520 524514 584960 524604
rect 576350 524454 584960 524514
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect -960 514798 3434 514858
rect -960 514708 480 514798
rect 3374 514612 3434 514798
rect 3374 514552 4048 514612
rect 583520 511322 584960 511412
rect 576350 511262 584960 511322
rect 576350 511196 576410 511262
rect 575920 511136 576410 511196
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect -960 501742 3434 501802
rect -960 501652 480 501742
rect 3374 501558 3434 501742
rect 3374 501498 4048 501558
rect 583520 497994 584960 498084
rect 576350 497934 584960 497994
rect 576350 497898 576410 497934
rect 575920 497838 576410 497898
rect 583520 497844 584960 497934
rect -960 488746 480 488836
rect -960 488686 3434 488746
rect -960 488596 480 488686
rect 3374 488504 3434 488686
rect 3374 488444 4048 488504
rect 583520 484666 584960 484756
rect 576350 484606 584960 484666
rect 576350 484600 576410 484606
rect 575920 484540 576410 484600
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect -960 475630 3434 475690
rect -960 475540 480 475630
rect 3374 475328 3434 475630
rect 3374 475268 4048 475328
rect 583520 471474 584960 471564
rect 576810 471414 584960 471474
rect 576810 471202 576870 471414
rect 583520 471324 584960 471414
rect 576350 471180 576870 471202
rect 575920 471142 576870 471180
rect 575920 471120 576410 471142
rect -960 462634 480 462724
rect -960 462574 3434 462634
rect -960 462484 480 462574
rect 3374 462274 3434 462574
rect 3374 462214 4048 462274
rect 583520 458146 584960 458236
rect 576810 458086 584960 458146
rect 576810 458010 576870 458086
rect 576350 457950 576870 458010
rect 583520 457996 584960 458086
rect 576350 457882 576410 457950
rect 575920 457822 576410 457882
rect -960 449578 480 449668
rect -960 449518 3434 449578
rect -960 449428 480 449518
rect 3374 449220 3434 449518
rect 3374 449160 4048 449220
rect 583520 444818 584960 444908
rect 576810 444758 584960 444818
rect 576810 444682 576870 444758
rect 576350 444622 576870 444682
rect 583520 444668 584960 444758
rect 576350 444584 576410 444622
rect 575920 444524 576410 444584
rect -960 436658 480 436748
rect 3417 436658 3483 436661
rect -960 436656 3483 436658
rect -960 436600 3422 436656
rect 3478 436600 3483 436656
rect -960 436598 3483 436600
rect -960 436508 480 436598
rect 3417 436595 3483 436598
rect 3417 436044 3483 436047
rect 3417 436042 4048 436044
rect 3417 435986 3422 436042
rect 3478 435986 4048 436042
rect 3417 435984 4048 435986
rect 3417 435981 3483 435984
rect 583520 431626 584960 431716
rect 583342 431566 584960 431626
rect 583342 431490 583402 431566
rect 583520 431490 584960 431566
rect 583342 431476 584960 431490
rect 583342 431430 583586 431476
rect 583526 431218 583586 431430
rect 576350 431164 583586 431218
rect 575920 431158 583586 431164
rect 575920 431104 576410 431158
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 3417 422990 3483 422993
rect 3417 422988 4048 422990
rect 3417 422932 3422 422988
rect 3478 422932 4048 422988
rect 3417 422930 4048 422932
rect 3417 422927 3483 422930
rect 583520 418298 584960 418388
rect 579662 418238 584960 418298
rect 579662 418162 579722 418238
rect 576810 418102 579722 418162
rect 583520 418148 584960 418238
rect 576810 417890 576870 418102
rect 576350 417866 576870 417890
rect 575920 417830 576870 417866
rect 575920 417806 576410 417830
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 3417 409936 3483 409939
rect 3417 409934 4048 409936
rect 3417 409878 3422 409934
rect 3478 409878 4048 409934
rect 3417 409876 4048 409878
rect 3417 409873 3483 409876
rect 583520 404970 584960 405060
rect 583342 404910 584960 404970
rect 583342 404834 583402 404910
rect 583520 404834 584960 404910
rect 583342 404820 584960 404834
rect 583342 404774 583586 404820
rect 583526 404562 583586 404774
rect 576350 404502 583586 404562
rect 576350 404446 576410 404502
rect 575920 404386 576410 404446
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 3417 396882 3483 396885
rect 3417 396880 4048 396882
rect 3417 396824 3422 396880
rect 3478 396824 4048 396880
rect 3417 396822 4048 396824
rect 3417 396819 3483 396822
rect 583520 391778 584960 391868
rect 583342 391718 584960 391778
rect 583342 391642 583402 391718
rect 583520 391642 584960 391718
rect 583342 391628 584960 391642
rect 583342 391582 583586 391628
rect 583526 391234 583586 391582
rect 576350 391174 583586 391234
rect 576350 391148 576410 391174
rect 575920 391088 576410 391148
rect -960 384434 480 384524
rect 3417 384434 3483 384437
rect -960 384432 3483 384434
rect -960 384376 3422 384432
rect 3478 384376 3483 384432
rect -960 384374 3483 384376
rect -960 384284 480 384374
rect 3417 384371 3483 384374
rect 3417 383706 3483 383709
rect 3417 383704 4048 383706
rect 3417 383648 3422 383704
rect 3478 383648 4048 383704
rect 3417 383646 4048 383648
rect 3417 383643 3483 383646
rect 583520 378450 584960 378540
rect 579662 378390 584960 378450
rect 579662 378178 579722 378390
rect 583520 378300 584960 378390
rect 579478 378118 579722 378178
rect 579478 377906 579538 378118
rect 576350 377850 579538 377906
rect 575920 377846 579538 377850
rect 575920 377790 576410 377846
rect -960 371378 480 371468
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 3417 370652 3483 370655
rect 3417 370650 4048 370652
rect 3417 370594 3422 370650
rect 3478 370594 4048 370650
rect 3417 370592 4048 370594
rect 3417 370589 3483 370592
rect 583520 365122 584960 365212
rect 583342 365062 584960 365122
rect 583342 364986 583402 365062
rect 583520 364986 584960 365062
rect 583342 364972 584960 364986
rect 583342 364926 583586 364972
rect 583526 364442 583586 364926
rect 576350 364430 583586 364442
rect 575920 364382 583586 364430
rect 575920 364370 576410 364382
rect -960 358458 480 358548
rect 3417 358458 3483 358461
rect -960 358456 3483 358458
rect -960 358400 3422 358456
rect 3478 358400 3483 358456
rect -960 358398 3483 358400
rect -960 358308 480 358398
rect 3417 358395 3483 358398
rect 3417 357598 3483 357601
rect 3417 357596 4048 357598
rect 3417 357540 3422 357596
rect 3478 357540 4048 357596
rect 3417 357538 4048 357540
rect 3417 357535 3483 357538
rect 579521 351930 579587 351933
rect 583520 351930 584960 352020
rect 579521 351928 584960 351930
rect 579521 351872 579526 351928
rect 579582 351872 584960 351928
rect 579521 351870 584960 351872
rect 579521 351867 579587 351870
rect 583520 351780 584960 351870
rect 575920 351114 576410 351132
rect 579521 351114 579587 351117
rect 575920 351112 579587 351114
rect 575920 351072 579526 351112
rect 576350 351056 579526 351072
rect 579582 351056 579587 351112
rect 576350 351054 579587 351056
rect 579521 351051 579587 351054
rect -960 345402 480 345492
rect 3417 345402 3483 345405
rect -960 345400 3483 345402
rect -960 345344 3422 345400
rect 3478 345344 3483 345400
rect -960 345342 3483 345344
rect -960 345252 480 345342
rect 3417 345339 3483 345342
rect 3417 344422 3483 344425
rect 3417 344420 4048 344422
rect 3417 344364 3422 344420
rect 3478 344364 4048 344420
rect 3417 344362 4048 344364
rect 3417 344359 3483 344362
rect 579613 338602 579679 338605
rect 583520 338602 584960 338692
rect 579613 338600 584960 338602
rect 579613 338544 579618 338600
rect 579674 338544 584960 338600
rect 579613 338542 584960 338544
rect 579613 338539 579679 338542
rect 583520 338452 584960 338542
rect 579521 337922 579587 337925
rect 576350 337920 579587 337922
rect 576350 337864 579526 337920
rect 579582 337864 579587 337920
rect 576350 337862 579587 337864
rect 576350 337834 576410 337862
rect 579521 337859 579587 337862
rect 575920 337774 576410 337834
rect -960 332346 480 332436
rect 3417 332346 3483 332349
rect -960 332344 3483 332346
rect -960 332288 3422 332344
rect 3478 332288 3483 332344
rect -960 332286 3483 332288
rect -960 332196 480 332286
rect 3417 332283 3483 332286
rect 3417 331368 3483 331371
rect 3417 331366 4048 331368
rect 3417 331310 3422 331366
rect 3478 331310 4048 331366
rect 3417 331308 4048 331310
rect 3417 331305 3483 331308
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 580165 324458 580231 324461
rect 576350 324456 580231 324458
rect 576350 324414 580170 324456
rect 575920 324400 580170 324414
rect 580226 324400 580231 324456
rect 575920 324398 580231 324400
rect 575920 324354 576410 324398
rect 580165 324395 580231 324398
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 3417 318314 3483 318317
rect 3417 318312 4048 318314
rect 3417 318256 3422 318312
rect 3478 318256 4048 318312
rect 3417 318254 4048 318256
rect 3417 318251 3483 318254
rect 579613 312082 579679 312085
rect 583520 312082 584960 312172
rect 579613 312080 584960 312082
rect 579613 312024 579618 312080
rect 579674 312024 584960 312080
rect 579613 312022 584960 312024
rect 579613 312019 579679 312022
rect 583520 311932 584960 312022
rect 579521 311130 579587 311133
rect 576350 311128 579587 311130
rect 576350 311116 579526 311128
rect 575920 311072 579526 311116
rect 579582 311072 579587 311128
rect 575920 311070 579587 311072
rect 575920 311056 576410 311070
rect 579521 311067 579587 311070
rect -960 306234 480 306324
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 3417 305138 3483 305141
rect 3417 305136 4048 305138
rect 3417 305080 3422 305136
rect 3478 305080 4048 305136
rect 3417 305078 4048 305080
rect 3417 305075 3483 305078
rect 579613 298754 579679 298757
rect 583520 298754 584960 298844
rect 579613 298752 584960 298754
rect 579613 298696 579618 298752
rect 579674 298696 584960 298752
rect 579613 298694 584960 298696
rect 579613 298691 579679 298694
rect 583520 298604 584960 298694
rect 575920 297802 576410 297818
rect 579521 297802 579587 297805
rect 575920 297800 579587 297802
rect 575920 297758 579526 297800
rect 576350 297744 579526 297758
rect 579582 297744 579587 297800
rect 576350 297742 579587 297744
rect 579521 297739 579587 297742
rect -960 293178 480 293268
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 3417 292084 3483 292087
rect 3417 292082 4048 292084
rect 3417 292026 3422 292082
rect 3478 292026 4048 292082
rect 3417 292024 4048 292026
rect 3417 292021 3483 292024
rect 580165 285426 580231 285429
rect 583520 285426 584960 285516
rect 580165 285424 584960 285426
rect 580165 285368 580170 285424
rect 580226 285368 584960 285424
rect 580165 285366 584960 285368
rect 580165 285363 580231 285366
rect 583520 285276 584960 285366
rect 580165 284474 580231 284477
rect 576350 284472 580231 284474
rect 576350 284416 580170 284472
rect 580226 284416 580231 284472
rect 576350 284414 580231 284416
rect 576350 284398 576410 284414
rect 580165 284411 580231 284414
rect 575920 284338 576410 284398
rect -960 280122 480 280212
rect 3417 280122 3483 280125
rect -960 280120 3483 280122
rect -960 280064 3422 280120
rect 3478 280064 3483 280120
rect -960 280062 3483 280064
rect -960 279972 480 280062
rect 3417 280059 3483 280062
rect 3417 279030 3483 279033
rect 3417 279028 4048 279030
rect 3417 278972 3422 279028
rect 3478 278972 4048 279028
rect 3417 278970 4048 278972
rect 3417 278967 3483 278970
rect 579613 272234 579679 272237
rect 583520 272234 584960 272324
rect 579613 272232 584960 272234
rect 579613 272176 579618 272232
rect 579674 272176 584960 272232
rect 579613 272174 584960 272176
rect 579613 272171 579679 272174
rect 583520 272084 584960 272174
rect 579521 271146 579587 271149
rect 576350 271144 579587 271146
rect 576350 271100 579526 271144
rect 575920 271088 579526 271100
rect 579582 271088 579587 271144
rect 575920 271086 579587 271088
rect 575920 271040 576410 271086
rect 579521 271083 579587 271086
rect -960 267202 480 267292
rect 3417 267202 3483 267205
rect -960 267200 3483 267202
rect -960 267144 3422 267200
rect 3478 267144 3483 267200
rect -960 267142 3483 267144
rect -960 267052 480 267142
rect 3417 267139 3483 267142
rect 3417 265976 3483 265979
rect 3417 265974 4048 265976
rect 3417 265918 3422 265974
rect 3478 265918 4048 265974
rect 3417 265916 4048 265918
rect 3417 265913 3483 265916
rect 580901 258906 580967 258909
rect 583520 258906 584960 258996
rect 580901 258904 584960 258906
rect 580901 258848 580906 258904
rect 580962 258848 584960 258904
rect 580901 258846 584960 258848
rect 580901 258843 580967 258846
rect 583520 258756 584960 258846
rect 578877 257682 578943 257685
rect 576350 257680 578943 257682
rect 575920 257624 578882 257680
rect 578938 257624 578943 257680
rect 575920 257622 578943 257624
rect 575920 257620 576410 257622
rect 578877 257619 578943 257622
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 3417 252800 3483 252803
rect 3417 252798 4048 252800
rect 3417 252742 3422 252798
rect 3478 252742 4048 252798
rect 3417 252740 4048 252742
rect 3417 252737 3483 252740
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 580165 244490 580231 244493
rect 576350 244488 580231 244490
rect 576350 244432 580170 244488
rect 580226 244432 580231 244488
rect 576350 244430 580231 244432
rect 576350 244382 576410 244430
rect 580165 244427 580231 244430
rect 575920 244322 576410 244382
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 3417 239746 3483 239749
rect 3417 239744 4048 239746
rect 3417 239688 3422 239744
rect 3478 239688 4048 239744
rect 3417 239686 4048 239688
rect 3417 239683 3483 239686
rect 579613 232386 579679 232389
rect 583520 232386 584960 232476
rect 579613 232384 584960 232386
rect 579613 232328 579618 232384
rect 579674 232328 584960 232384
rect 579613 232326 584960 232328
rect 579613 232323 579679 232326
rect 583520 232236 584960 232326
rect 579521 231162 579587 231165
rect 576350 231160 579587 231162
rect 576350 231104 579526 231160
rect 579582 231104 579587 231160
rect 576350 231102 579587 231104
rect 576350 231084 576410 231102
rect 579521 231099 579587 231102
rect 575920 231024 576410 231084
rect -960 228034 480 228124
rect 3417 228034 3483 228037
rect -960 228032 3483 228034
rect -960 227976 3422 228032
rect 3478 227976 3483 228032
rect -960 227974 3483 227976
rect -960 227884 480 227974
rect 3417 227971 3483 227974
rect 3417 226692 3483 226695
rect 3417 226690 4048 226692
rect 3417 226634 3422 226690
rect 3478 226634 4048 226690
rect 3417 226632 4048 226634
rect 3417 226629 3483 226632
rect 579613 219058 579679 219061
rect 583520 219058 584960 219148
rect 579613 219056 584960 219058
rect 579613 219000 579618 219056
rect 579674 219000 584960 219056
rect 579613 218998 584960 219000
rect 579613 218995 579679 218998
rect 583520 218908 584960 218998
rect 579521 217698 579587 217701
rect 576350 217696 579587 217698
rect 576350 217664 579526 217696
rect 575920 217640 579526 217664
rect 579582 217640 579587 217696
rect 575920 217638 579587 217640
rect 575920 217604 576410 217638
rect 579521 217635 579587 217638
rect -960 214978 480 215068
rect 3417 214978 3483 214981
rect -960 214976 3483 214978
rect -960 214920 3422 214976
rect 3478 214920 3483 214976
rect -960 214918 3483 214920
rect -960 214828 480 214918
rect 3417 214915 3483 214918
rect 3417 213516 3483 213519
rect 3417 213514 4048 213516
rect 3417 213458 3422 213514
rect 3478 213458 4048 213514
rect 3417 213456 4048 213458
rect 3417 213453 3483 213456
rect 579613 205730 579679 205733
rect 583520 205730 584960 205820
rect 579613 205728 584960 205730
rect 579613 205672 579618 205728
rect 579674 205672 584960 205728
rect 579613 205670 584960 205672
rect 579613 205667 579679 205670
rect 583520 205580 584960 205670
rect 579521 204370 579587 204373
rect 576350 204368 579587 204370
rect 576350 204366 579526 204368
rect 575920 204312 579526 204366
rect 579582 204312 579587 204368
rect 575920 204310 579587 204312
rect 575920 204306 576410 204310
rect 579521 204307 579587 204310
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 3417 200462 3483 200465
rect 3417 200460 4048 200462
rect 3417 200404 3422 200460
rect 3478 200404 4048 200460
rect 3417 200402 4048 200404
rect 3417 200399 3483 200402
rect 579613 192538 579679 192541
rect 583520 192538 584960 192628
rect 579613 192536 584960 192538
rect 579613 192480 579618 192536
rect 579674 192480 584960 192536
rect 579613 192478 584960 192480
rect 579613 192475 579679 192478
rect 583520 192388 584960 192478
rect 575920 191042 576410 191068
rect 579521 191042 579587 191045
rect 575920 191040 579587 191042
rect 575920 191008 579526 191040
rect 576350 190984 579526 191008
rect 579582 190984 579587 191040
rect 576350 190982 579587 190984
rect 579521 190979 579587 190982
rect -960 188866 480 188956
rect 3601 188866 3667 188869
rect -960 188864 3667 188866
rect -960 188808 3606 188864
rect 3662 188808 3667 188864
rect -960 188806 3667 188808
rect -960 188716 480 188806
rect 3601 188803 3667 188806
rect 3601 187408 3667 187411
rect 3601 187406 4048 187408
rect 3601 187350 3606 187406
rect 3662 187350 4048 187406
rect 3601 187348 4048 187350
rect 3601 187345 3667 187348
rect 579613 179210 579679 179213
rect 583520 179210 584960 179300
rect 579613 179208 584960 179210
rect 579613 179152 579618 179208
rect 579674 179152 584960 179208
rect 579613 179150 584960 179152
rect 579613 179147 579679 179150
rect 583520 179060 584960 179150
rect 579521 177714 579587 177717
rect 576350 177712 579587 177714
rect 576350 177656 579526 177712
rect 579582 177656 579587 177712
rect 576350 177654 579587 177656
rect 576350 177648 576410 177654
rect 579521 177651 579587 177654
rect 575920 177588 576410 177648
rect -960 175946 480 176036
rect 3417 175946 3483 175949
rect -960 175944 3483 175946
rect -960 175888 3422 175944
rect 3478 175888 3483 175944
rect -960 175886 3483 175888
rect -960 175796 480 175886
rect 3417 175883 3483 175886
rect 3417 174232 3483 174235
rect 3417 174230 4048 174232
rect 3417 174174 3422 174230
rect 3478 174174 4048 174230
rect 3417 174172 4048 174174
rect 3417 174169 3483 174172
rect 579613 165882 579679 165885
rect 583520 165882 584960 165972
rect 579613 165880 584960 165882
rect 579613 165824 579618 165880
rect 579674 165824 584960 165880
rect 579613 165822 584960 165824
rect 579613 165819 579679 165822
rect 583520 165732 584960 165822
rect 579521 164386 579587 164389
rect 576350 164384 579587 164386
rect 576350 164350 579526 164384
rect 575920 164328 579526 164350
rect 579582 164328 579587 164384
rect 575920 164326 579587 164328
rect 575920 164290 576410 164326
rect 579521 164323 579587 164326
rect -960 162890 480 162980
rect 2129 162890 2195 162893
rect -960 162888 2195 162890
rect -960 162832 2134 162888
rect 2190 162832 2195 162888
rect -960 162830 2195 162832
rect -960 162740 480 162830
rect 2129 162827 2195 162830
rect 2129 161122 2195 161125
rect 3374 161122 4048 161178
rect 2129 161120 4048 161122
rect 2129 161064 2134 161120
rect 2190 161118 4048 161120
rect 2190 161064 3434 161118
rect 2129 161062 3434 161064
rect 2129 161059 2195 161062
rect 580901 152690 580967 152693
rect 583520 152690 584960 152780
rect 580901 152688 584960 152690
rect 580901 152632 580906 152688
rect 580962 152632 584960 152688
rect 580901 152630 584960 152632
rect 580901 152627 580967 152630
rect 583520 152540 584960 152630
rect 578509 151058 578575 151061
rect 576350 151056 578575 151058
rect 576350 151052 578514 151056
rect 575920 151000 578514 151052
rect 578570 151000 578575 151056
rect 575920 150998 578575 151000
rect 575920 150992 576410 150998
rect 578509 150995 578575 150998
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 3417 148124 3483 148127
rect 3417 148122 4048 148124
rect 3417 148066 3422 148122
rect 3478 148066 4048 148122
rect 3417 148064 4048 148066
rect 3417 148061 3483 148064
rect 579613 139362 579679 139365
rect 583520 139362 584960 139452
rect 579613 139360 584960 139362
rect 579613 139304 579618 139360
rect 579674 139304 584960 139360
rect 579613 139302 584960 139304
rect 579613 139299 579679 139302
rect 583520 139212 584960 139302
rect 575920 137594 576410 137632
rect 579521 137594 579587 137597
rect 575920 137592 579587 137594
rect 575920 137572 579526 137592
rect 576350 137536 579526 137572
rect 579582 137536 579587 137592
rect 576350 137534 579587 137536
rect 579521 137531 579587 137534
rect -960 136778 480 136868
rect 2129 136778 2195 136781
rect -960 136776 2195 136778
rect -960 136720 2134 136776
rect 2190 136720 2195 136776
rect -960 136718 2195 136720
rect -960 136628 480 136718
rect 2129 136715 2195 136718
rect 2129 135010 2195 135013
rect 3374 135010 4048 135070
rect 2129 135008 3434 135010
rect 2129 134952 2134 135008
rect 2190 134952 3434 135008
rect 2129 134950 3434 134952
rect 2129 134947 2195 134950
rect 579613 126034 579679 126037
rect 583520 126034 584960 126124
rect 579613 126032 584960 126034
rect 579613 125976 579618 126032
rect 579674 125976 584960 126032
rect 579613 125974 584960 125976
rect 579613 125971 579679 125974
rect 583520 125884 584960 125974
rect 579521 124402 579587 124405
rect 576350 124400 579587 124402
rect 576350 124344 579526 124400
rect 579582 124344 579587 124400
rect 576350 124342 579587 124344
rect 576350 124334 576410 124342
rect 579521 124339 579587 124342
rect 575920 124274 576410 124334
rect -960 123722 480 123812
rect 3417 123722 3483 123725
rect -960 123720 3483 123722
rect -960 123664 3422 123720
rect 3478 123664 3483 123720
rect -960 123662 3483 123664
rect -960 123572 480 123662
rect 3417 123659 3483 123662
rect 3417 121894 3483 121897
rect 3417 121892 4048 121894
rect 3417 121836 3422 121892
rect 3478 121836 4048 121892
rect 3417 121834 4048 121836
rect 3417 121831 3483 121834
rect 579613 112842 579679 112845
rect 583520 112842 584960 112932
rect 579613 112840 584960 112842
rect 579613 112784 579618 112840
rect 579674 112784 584960 112840
rect 579613 112782 584960 112784
rect 579613 112779 579679 112782
rect 583520 112692 584960 112782
rect 579521 110938 579587 110941
rect 576350 110936 579587 110938
rect 576350 110914 579526 110936
rect 575920 110880 579526 110914
rect 579582 110880 579587 110936
rect 575920 110878 579587 110880
rect 575920 110854 576410 110878
rect 579521 110875 579587 110878
rect -960 110666 480 110756
rect 2129 110666 2195 110669
rect -960 110664 2195 110666
rect -960 110608 2134 110664
rect 2190 110608 2195 110664
rect -960 110606 2195 110608
rect -960 110516 480 110606
rect 2129 110603 2195 110606
rect 2129 108898 2195 108901
rect 2129 108896 3434 108898
rect 2129 108840 2134 108896
rect 2190 108840 3434 108896
rect 2129 108838 4048 108840
rect 2129 108835 2195 108838
rect 3374 108780 4048 108838
rect 579613 99514 579679 99517
rect 583520 99514 584960 99604
rect 579613 99512 584960 99514
rect 579613 99456 579618 99512
rect 579674 99456 584960 99512
rect 579613 99454 584960 99456
rect 579613 99451 579679 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect 575920 97610 576410 97616
rect 579521 97610 579587 97613
rect 575920 97608 579587 97610
rect 575920 97556 579526 97608
rect -960 97550 3483 97552
rect 576350 97552 579526 97556
rect 579582 97552 579587 97608
rect 576350 97550 579587 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 579521 97547 579587 97550
rect 3417 95786 3483 95789
rect 3417 95784 4048 95786
rect 3417 95728 3422 95784
rect 3478 95728 4048 95784
rect 3417 95726 4048 95728
rect 3417 95723 3483 95726
rect 579613 86186 579679 86189
rect 583520 86186 584960 86276
rect 579613 86184 584960 86186
rect 579613 86128 579618 86184
rect 579674 86128 584960 86184
rect 579613 86126 584960 86128
rect 579613 86123 579679 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 2129 84690 2195 84693
rect -960 84688 2195 84690
rect -960 84632 2134 84688
rect 2190 84632 2195 84688
rect -960 84630 2195 84632
rect -960 84540 480 84630
rect 2129 84627 2195 84630
rect 575920 84282 576410 84318
rect 579521 84282 579587 84285
rect 575920 84280 579587 84282
rect 575920 84258 579526 84280
rect 576350 84224 579526 84258
rect 579582 84224 579587 84280
rect 576350 84222 579587 84224
rect 579521 84219 579587 84222
rect 2129 82650 2195 82653
rect 2129 82648 3434 82650
rect 2129 82592 2134 82648
rect 2190 82610 3434 82648
rect 2190 82592 4048 82610
rect 2129 82590 4048 82592
rect 2129 82587 2195 82590
rect 3374 82550 4048 82590
rect 579613 72994 579679 72997
rect 583520 72994 584960 73084
rect 579613 72992 584960 72994
rect 579613 72936 579618 72992
rect 579674 72936 584960 72992
rect 579613 72934 584960 72936
rect 579613 72931 579679 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 579521 70954 579587 70957
rect 576350 70952 579587 70954
rect 576350 70898 579526 70952
rect 575920 70896 579526 70898
rect 579582 70896 579587 70952
rect 575920 70894 579587 70896
rect 575920 70838 576410 70894
rect 579521 70891 579587 70894
rect 3417 69556 3483 69559
rect 3417 69554 4048 69556
rect 3417 69498 3422 69554
rect 3478 69498 4048 69554
rect 3417 69496 4048 69498
rect 3417 69493 3483 69496
rect 579613 59666 579679 59669
rect 583520 59666 584960 59756
rect 579613 59664 584960 59666
rect 579613 59608 579618 59664
rect 579674 59608 584960 59664
rect 579613 59606 584960 59608
rect 579613 59603 579679 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 2129 58578 2195 58581
rect -960 58576 2195 58578
rect -960 58520 2134 58576
rect 2190 58520 2195 58576
rect -960 58518 2195 58520
rect -960 58428 480 58518
rect 2129 58515 2195 58518
rect 579521 57626 579587 57629
rect 576350 57624 579587 57626
rect 576350 57600 579526 57624
rect 575920 57568 579526 57600
rect 579582 57568 579587 57624
rect 575920 57566 579587 57568
rect 575920 57540 576410 57566
rect 579521 57563 579587 57566
rect 2129 56538 2195 56541
rect 2129 56536 3434 56538
rect 2129 56480 2134 56536
rect 2190 56502 3434 56536
rect 2190 56480 4048 56502
rect 2129 56478 4048 56480
rect 2129 56475 2195 56478
rect 3374 56442 4048 56478
rect 579981 46338 580047 46341
rect 583520 46338 584960 46428
rect 579981 46336 584960 46338
rect 579981 46280 579986 46336
rect 580042 46280 584960 46336
rect 579981 46278 584960 46280
rect 579981 46275 580047 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 575920 44298 576410 44302
rect 578325 44298 578391 44301
rect 575920 44296 578391 44298
rect 575920 44242 578330 44296
rect 576350 44240 578330 44242
rect 578386 44240 578391 44296
rect 576350 44238 578391 44240
rect 578325 44235 578391 44238
rect 3417 43326 3483 43329
rect 3417 43324 4048 43326
rect 3417 43268 3422 43324
rect 3478 43268 4048 43324
rect 3417 43266 4048 43268
rect 3417 43263 3483 43266
rect 579613 33146 579679 33149
rect 583520 33146 584960 33236
rect 579613 33144 584960 33146
rect 579613 33088 579618 33144
rect 579674 33088 584960 33144
rect 579613 33086 584960 33088
rect 579613 33083 579679 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2129 32466 2195 32469
rect -960 32464 2195 32466
rect -960 32408 2134 32464
rect 2190 32408 2195 32464
rect -960 32406 2195 32408
rect -960 32316 480 32406
rect 2129 32403 2195 32406
rect 579521 30970 579587 30973
rect 576350 30968 579587 30970
rect 576350 30912 579526 30968
rect 579582 30912 579587 30968
rect 576350 30910 579587 30912
rect 576350 30882 576410 30910
rect 579521 30907 579587 30910
rect 575920 30822 576410 30882
rect 2129 30290 2195 30293
rect 2129 30288 3434 30290
rect 2129 30232 2134 30288
rect 2190 30272 3434 30288
rect 2190 30232 4048 30272
rect 2129 30230 4048 30232
rect 2129 30227 2195 30230
rect 3374 30212 4048 30230
rect 579613 19818 579679 19821
rect 583520 19818 584960 19908
rect 579613 19816 584960 19818
rect 579613 19760 579618 19816
rect 579674 19760 584960 19816
rect 579613 19758 584960 19760
rect 579613 19755 579679 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 2037 19410 2103 19413
rect -960 19408 2103 19410
rect -960 19352 2042 19408
rect 2098 19352 2103 19408
rect -960 19350 2103 19352
rect -960 19260 480 19350
rect 2037 19347 2103 19350
rect 579521 17642 579587 17645
rect 576350 17640 579587 17642
rect 576350 17584 579526 17640
rect 579582 17584 579587 17640
rect 575920 17582 579587 17584
rect 575920 17524 576410 17582
rect 579521 17579 579587 17582
rect 2037 17234 2103 17237
rect 2037 17232 3434 17234
rect 2037 17176 2042 17232
rect 2098 17218 3434 17232
rect 2098 17176 4048 17218
rect 2037 17174 4048 17176
rect 2037 17171 2103 17174
rect 3374 17158 4048 17174
rect 579613 6626 579679 6629
rect 583520 6626 584960 6716
rect 579613 6624 584960 6626
rect -960 6490 480 6580
rect 579613 6568 579618 6624
rect 579674 6568 584960 6624
rect 579613 6566 584960 6568
rect 579613 6563 579679 6566
rect 2773 6490 2839 6493
rect -960 6488 2839 6490
rect -960 6432 2778 6488
rect 2834 6432 2839 6488
rect 583520 6476 584960 6566
rect -960 6430 2839 6432
rect -960 6340 480 6430
rect 2773 6427 2839 6430
rect 2773 4178 2839 4181
rect 576761 4178 576827 4181
rect 2773 4176 3802 4178
rect 2773 4120 2778 4176
rect 2834 4164 3802 4176
rect 576350 4176 576827 4178
rect 576350 4164 576766 4176
rect 2834 4120 4048 4164
rect 2773 4118 4048 4120
rect 2773 4115 2839 4118
rect 3742 4104 4048 4118
rect 575920 4120 576766 4164
rect 576822 4120 576827 4176
rect 575920 4118 576827 4120
rect 575920 4104 576410 4118
rect 576761 4115 576827 4118
<< metal4 >>
rect -23776 726608 -23156 726640
rect -23776 726372 -23744 726608
rect -23508 726372 -23424 726608
rect -23188 726372 -23156 726608
rect -23776 726288 -23156 726372
rect -23776 726052 -23744 726288
rect -23508 726052 -23424 726288
rect -23188 726052 -23156 726288
rect -23776 677494 -23156 726052
rect -23776 677258 -23744 677494
rect -23508 677258 -23424 677494
rect -23188 677258 -23156 677494
rect -23776 677174 -23156 677258
rect -23776 676938 -23744 677174
rect -23508 676938 -23424 677174
rect -23188 676938 -23156 677174
rect -23776 641494 -23156 676938
rect -23776 641258 -23744 641494
rect -23508 641258 -23424 641494
rect -23188 641258 -23156 641494
rect -23776 641174 -23156 641258
rect -23776 640938 -23744 641174
rect -23508 640938 -23424 641174
rect -23188 640938 -23156 641174
rect -23776 605494 -23156 640938
rect -23776 605258 -23744 605494
rect -23508 605258 -23424 605494
rect -23188 605258 -23156 605494
rect -23776 605174 -23156 605258
rect -23776 604938 -23744 605174
rect -23508 604938 -23424 605174
rect -23188 604938 -23156 605174
rect -23776 569494 -23156 604938
rect -23776 569258 -23744 569494
rect -23508 569258 -23424 569494
rect -23188 569258 -23156 569494
rect -23776 569174 -23156 569258
rect -23776 568938 -23744 569174
rect -23508 568938 -23424 569174
rect -23188 568938 -23156 569174
rect -23776 533494 -23156 568938
rect -23776 533258 -23744 533494
rect -23508 533258 -23424 533494
rect -23188 533258 -23156 533494
rect -23776 533174 -23156 533258
rect -23776 532938 -23744 533174
rect -23508 532938 -23424 533174
rect -23188 532938 -23156 533174
rect -23776 497494 -23156 532938
rect -23776 497258 -23744 497494
rect -23508 497258 -23424 497494
rect -23188 497258 -23156 497494
rect -23776 497174 -23156 497258
rect -23776 496938 -23744 497174
rect -23508 496938 -23424 497174
rect -23188 496938 -23156 497174
rect -23776 461494 -23156 496938
rect -23776 461258 -23744 461494
rect -23508 461258 -23424 461494
rect -23188 461258 -23156 461494
rect -23776 461174 -23156 461258
rect -23776 460938 -23744 461174
rect -23508 460938 -23424 461174
rect -23188 460938 -23156 461174
rect -23776 425494 -23156 460938
rect -23776 425258 -23744 425494
rect -23508 425258 -23424 425494
rect -23188 425258 -23156 425494
rect -23776 425174 -23156 425258
rect -23776 424938 -23744 425174
rect -23508 424938 -23424 425174
rect -23188 424938 -23156 425174
rect -23776 389494 -23156 424938
rect -23776 389258 -23744 389494
rect -23508 389258 -23424 389494
rect -23188 389258 -23156 389494
rect -23776 389174 -23156 389258
rect -23776 388938 -23744 389174
rect -23508 388938 -23424 389174
rect -23188 388938 -23156 389174
rect -23776 353494 -23156 388938
rect -23776 353258 -23744 353494
rect -23508 353258 -23424 353494
rect -23188 353258 -23156 353494
rect -23776 353174 -23156 353258
rect -23776 352938 -23744 353174
rect -23508 352938 -23424 353174
rect -23188 352938 -23156 353174
rect -23776 317494 -23156 352938
rect -23776 317258 -23744 317494
rect -23508 317258 -23424 317494
rect -23188 317258 -23156 317494
rect -23776 317174 -23156 317258
rect -23776 316938 -23744 317174
rect -23508 316938 -23424 317174
rect -23188 316938 -23156 317174
rect -23776 281494 -23156 316938
rect -23776 281258 -23744 281494
rect -23508 281258 -23424 281494
rect -23188 281258 -23156 281494
rect -23776 281174 -23156 281258
rect -23776 280938 -23744 281174
rect -23508 280938 -23424 281174
rect -23188 280938 -23156 281174
rect -23776 245494 -23156 280938
rect -23776 245258 -23744 245494
rect -23508 245258 -23424 245494
rect -23188 245258 -23156 245494
rect -23776 245174 -23156 245258
rect -23776 244938 -23744 245174
rect -23508 244938 -23424 245174
rect -23188 244938 -23156 245174
rect -23776 209494 -23156 244938
rect -23776 209258 -23744 209494
rect -23508 209258 -23424 209494
rect -23188 209258 -23156 209494
rect -23776 209174 -23156 209258
rect -23776 208938 -23744 209174
rect -23508 208938 -23424 209174
rect -23188 208938 -23156 209174
rect -23776 173494 -23156 208938
rect -23776 173258 -23744 173494
rect -23508 173258 -23424 173494
rect -23188 173258 -23156 173494
rect -23776 173174 -23156 173258
rect -23776 172938 -23744 173174
rect -23508 172938 -23424 173174
rect -23188 172938 -23156 173174
rect -23776 137494 -23156 172938
rect -23776 137258 -23744 137494
rect -23508 137258 -23424 137494
rect -23188 137258 -23156 137494
rect -23776 137174 -23156 137258
rect -23776 136938 -23744 137174
rect -23508 136938 -23424 137174
rect -23188 136938 -23156 137174
rect -23776 101494 -23156 136938
rect -23776 101258 -23744 101494
rect -23508 101258 -23424 101494
rect -23188 101258 -23156 101494
rect -23776 101174 -23156 101258
rect -23776 100938 -23744 101174
rect -23508 100938 -23424 101174
rect -23188 100938 -23156 101174
rect -23776 65494 -23156 100938
rect -23776 65258 -23744 65494
rect -23508 65258 -23424 65494
rect -23188 65258 -23156 65494
rect -23776 65174 -23156 65258
rect -23776 64938 -23744 65174
rect -23508 64938 -23424 65174
rect -23188 64938 -23156 65174
rect -23776 29494 -23156 64938
rect -23776 29258 -23744 29494
rect -23508 29258 -23424 29494
rect -23188 29258 -23156 29494
rect -23776 29174 -23156 29258
rect -23776 28938 -23744 29174
rect -23508 28938 -23424 29174
rect -23188 28938 -23156 29174
rect -23776 -22116 -23156 28938
rect -20666 723498 -20046 723530
rect -20666 723262 -20634 723498
rect -20398 723262 -20314 723498
rect -20078 723262 -20046 723498
rect -20666 723178 -20046 723262
rect -20666 722942 -20634 723178
rect -20398 722942 -20314 723178
rect -20078 722942 -20046 723178
rect -20666 673774 -20046 722942
rect -20666 673538 -20634 673774
rect -20398 673538 -20314 673774
rect -20078 673538 -20046 673774
rect -20666 673454 -20046 673538
rect -20666 673218 -20634 673454
rect -20398 673218 -20314 673454
rect -20078 673218 -20046 673454
rect -20666 637774 -20046 673218
rect -20666 637538 -20634 637774
rect -20398 637538 -20314 637774
rect -20078 637538 -20046 637774
rect -20666 637454 -20046 637538
rect -20666 637218 -20634 637454
rect -20398 637218 -20314 637454
rect -20078 637218 -20046 637454
rect -20666 601774 -20046 637218
rect -20666 601538 -20634 601774
rect -20398 601538 -20314 601774
rect -20078 601538 -20046 601774
rect -20666 601454 -20046 601538
rect -20666 601218 -20634 601454
rect -20398 601218 -20314 601454
rect -20078 601218 -20046 601454
rect -20666 565774 -20046 601218
rect -20666 565538 -20634 565774
rect -20398 565538 -20314 565774
rect -20078 565538 -20046 565774
rect -20666 565454 -20046 565538
rect -20666 565218 -20634 565454
rect -20398 565218 -20314 565454
rect -20078 565218 -20046 565454
rect -20666 529774 -20046 565218
rect -20666 529538 -20634 529774
rect -20398 529538 -20314 529774
rect -20078 529538 -20046 529774
rect -20666 529454 -20046 529538
rect -20666 529218 -20634 529454
rect -20398 529218 -20314 529454
rect -20078 529218 -20046 529454
rect -20666 493774 -20046 529218
rect -20666 493538 -20634 493774
rect -20398 493538 -20314 493774
rect -20078 493538 -20046 493774
rect -20666 493454 -20046 493538
rect -20666 493218 -20634 493454
rect -20398 493218 -20314 493454
rect -20078 493218 -20046 493454
rect -20666 457774 -20046 493218
rect -20666 457538 -20634 457774
rect -20398 457538 -20314 457774
rect -20078 457538 -20046 457774
rect -20666 457454 -20046 457538
rect -20666 457218 -20634 457454
rect -20398 457218 -20314 457454
rect -20078 457218 -20046 457454
rect -20666 421774 -20046 457218
rect -20666 421538 -20634 421774
rect -20398 421538 -20314 421774
rect -20078 421538 -20046 421774
rect -20666 421454 -20046 421538
rect -20666 421218 -20634 421454
rect -20398 421218 -20314 421454
rect -20078 421218 -20046 421454
rect -20666 385774 -20046 421218
rect -20666 385538 -20634 385774
rect -20398 385538 -20314 385774
rect -20078 385538 -20046 385774
rect -20666 385454 -20046 385538
rect -20666 385218 -20634 385454
rect -20398 385218 -20314 385454
rect -20078 385218 -20046 385454
rect -20666 349774 -20046 385218
rect -20666 349538 -20634 349774
rect -20398 349538 -20314 349774
rect -20078 349538 -20046 349774
rect -20666 349454 -20046 349538
rect -20666 349218 -20634 349454
rect -20398 349218 -20314 349454
rect -20078 349218 -20046 349454
rect -20666 313774 -20046 349218
rect -20666 313538 -20634 313774
rect -20398 313538 -20314 313774
rect -20078 313538 -20046 313774
rect -20666 313454 -20046 313538
rect -20666 313218 -20634 313454
rect -20398 313218 -20314 313454
rect -20078 313218 -20046 313454
rect -20666 277774 -20046 313218
rect -20666 277538 -20634 277774
rect -20398 277538 -20314 277774
rect -20078 277538 -20046 277774
rect -20666 277454 -20046 277538
rect -20666 277218 -20634 277454
rect -20398 277218 -20314 277454
rect -20078 277218 -20046 277454
rect -20666 241774 -20046 277218
rect -20666 241538 -20634 241774
rect -20398 241538 -20314 241774
rect -20078 241538 -20046 241774
rect -20666 241454 -20046 241538
rect -20666 241218 -20634 241454
rect -20398 241218 -20314 241454
rect -20078 241218 -20046 241454
rect -20666 205774 -20046 241218
rect -20666 205538 -20634 205774
rect -20398 205538 -20314 205774
rect -20078 205538 -20046 205774
rect -20666 205454 -20046 205538
rect -20666 205218 -20634 205454
rect -20398 205218 -20314 205454
rect -20078 205218 -20046 205454
rect -20666 169774 -20046 205218
rect -20666 169538 -20634 169774
rect -20398 169538 -20314 169774
rect -20078 169538 -20046 169774
rect -20666 169454 -20046 169538
rect -20666 169218 -20634 169454
rect -20398 169218 -20314 169454
rect -20078 169218 -20046 169454
rect -20666 133774 -20046 169218
rect -20666 133538 -20634 133774
rect -20398 133538 -20314 133774
rect -20078 133538 -20046 133774
rect -20666 133454 -20046 133538
rect -20666 133218 -20634 133454
rect -20398 133218 -20314 133454
rect -20078 133218 -20046 133454
rect -20666 97774 -20046 133218
rect -20666 97538 -20634 97774
rect -20398 97538 -20314 97774
rect -20078 97538 -20046 97774
rect -20666 97454 -20046 97538
rect -20666 97218 -20634 97454
rect -20398 97218 -20314 97454
rect -20078 97218 -20046 97454
rect -20666 61774 -20046 97218
rect -20666 61538 -20634 61774
rect -20398 61538 -20314 61774
rect -20078 61538 -20046 61774
rect -20666 61454 -20046 61538
rect -20666 61218 -20634 61454
rect -20398 61218 -20314 61454
rect -20078 61218 -20046 61454
rect -20666 25774 -20046 61218
rect -20666 25538 -20634 25774
rect -20398 25538 -20314 25774
rect -20078 25538 -20046 25774
rect -20666 25454 -20046 25538
rect -20666 25218 -20634 25454
rect -20398 25218 -20314 25454
rect -20078 25218 -20046 25454
rect -20666 -19006 -20046 25218
rect -17556 720388 -16936 720420
rect -17556 720152 -17524 720388
rect -17288 720152 -17204 720388
rect -16968 720152 -16936 720388
rect -17556 720068 -16936 720152
rect -17556 719832 -17524 720068
rect -17288 719832 -17204 720068
rect -16968 719832 -16936 720068
rect -17556 670054 -16936 719832
rect -17556 669818 -17524 670054
rect -17288 669818 -17204 670054
rect -16968 669818 -16936 670054
rect -17556 669734 -16936 669818
rect -17556 669498 -17524 669734
rect -17288 669498 -17204 669734
rect -16968 669498 -16936 669734
rect -17556 634054 -16936 669498
rect -17556 633818 -17524 634054
rect -17288 633818 -17204 634054
rect -16968 633818 -16936 634054
rect -17556 633734 -16936 633818
rect -17556 633498 -17524 633734
rect -17288 633498 -17204 633734
rect -16968 633498 -16936 633734
rect -17556 598054 -16936 633498
rect -17556 597818 -17524 598054
rect -17288 597818 -17204 598054
rect -16968 597818 -16936 598054
rect -17556 597734 -16936 597818
rect -17556 597498 -17524 597734
rect -17288 597498 -17204 597734
rect -16968 597498 -16936 597734
rect -17556 562054 -16936 597498
rect -17556 561818 -17524 562054
rect -17288 561818 -17204 562054
rect -16968 561818 -16936 562054
rect -17556 561734 -16936 561818
rect -17556 561498 -17524 561734
rect -17288 561498 -17204 561734
rect -16968 561498 -16936 561734
rect -17556 526054 -16936 561498
rect -17556 525818 -17524 526054
rect -17288 525818 -17204 526054
rect -16968 525818 -16936 526054
rect -17556 525734 -16936 525818
rect -17556 525498 -17524 525734
rect -17288 525498 -17204 525734
rect -16968 525498 -16936 525734
rect -17556 490054 -16936 525498
rect -17556 489818 -17524 490054
rect -17288 489818 -17204 490054
rect -16968 489818 -16936 490054
rect -17556 489734 -16936 489818
rect -17556 489498 -17524 489734
rect -17288 489498 -17204 489734
rect -16968 489498 -16936 489734
rect -17556 454054 -16936 489498
rect -17556 453818 -17524 454054
rect -17288 453818 -17204 454054
rect -16968 453818 -16936 454054
rect -17556 453734 -16936 453818
rect -17556 453498 -17524 453734
rect -17288 453498 -17204 453734
rect -16968 453498 -16936 453734
rect -17556 418054 -16936 453498
rect -17556 417818 -17524 418054
rect -17288 417818 -17204 418054
rect -16968 417818 -16936 418054
rect -17556 417734 -16936 417818
rect -17556 417498 -17524 417734
rect -17288 417498 -17204 417734
rect -16968 417498 -16936 417734
rect -17556 382054 -16936 417498
rect -17556 381818 -17524 382054
rect -17288 381818 -17204 382054
rect -16968 381818 -16936 382054
rect -17556 381734 -16936 381818
rect -17556 381498 -17524 381734
rect -17288 381498 -17204 381734
rect -16968 381498 -16936 381734
rect -17556 346054 -16936 381498
rect -17556 345818 -17524 346054
rect -17288 345818 -17204 346054
rect -16968 345818 -16936 346054
rect -17556 345734 -16936 345818
rect -17556 345498 -17524 345734
rect -17288 345498 -17204 345734
rect -16968 345498 -16936 345734
rect -17556 310054 -16936 345498
rect -17556 309818 -17524 310054
rect -17288 309818 -17204 310054
rect -16968 309818 -16936 310054
rect -17556 309734 -16936 309818
rect -17556 309498 -17524 309734
rect -17288 309498 -17204 309734
rect -16968 309498 -16936 309734
rect -17556 274054 -16936 309498
rect -17556 273818 -17524 274054
rect -17288 273818 -17204 274054
rect -16968 273818 -16936 274054
rect -17556 273734 -16936 273818
rect -17556 273498 -17524 273734
rect -17288 273498 -17204 273734
rect -16968 273498 -16936 273734
rect -17556 238054 -16936 273498
rect -17556 237818 -17524 238054
rect -17288 237818 -17204 238054
rect -16968 237818 -16936 238054
rect -17556 237734 -16936 237818
rect -17556 237498 -17524 237734
rect -17288 237498 -17204 237734
rect -16968 237498 -16936 237734
rect -17556 202054 -16936 237498
rect -17556 201818 -17524 202054
rect -17288 201818 -17204 202054
rect -16968 201818 -16936 202054
rect -17556 201734 -16936 201818
rect -17556 201498 -17524 201734
rect -17288 201498 -17204 201734
rect -16968 201498 -16936 201734
rect -17556 166054 -16936 201498
rect -17556 165818 -17524 166054
rect -17288 165818 -17204 166054
rect -16968 165818 -16936 166054
rect -17556 165734 -16936 165818
rect -17556 165498 -17524 165734
rect -17288 165498 -17204 165734
rect -16968 165498 -16936 165734
rect -17556 130054 -16936 165498
rect -17556 129818 -17524 130054
rect -17288 129818 -17204 130054
rect -16968 129818 -16936 130054
rect -17556 129734 -16936 129818
rect -17556 129498 -17524 129734
rect -17288 129498 -17204 129734
rect -16968 129498 -16936 129734
rect -17556 94054 -16936 129498
rect -17556 93818 -17524 94054
rect -17288 93818 -17204 94054
rect -16968 93818 -16936 94054
rect -17556 93734 -16936 93818
rect -17556 93498 -17524 93734
rect -17288 93498 -17204 93734
rect -16968 93498 -16936 93734
rect -17556 58054 -16936 93498
rect -17556 57818 -17524 58054
rect -17288 57818 -17204 58054
rect -16968 57818 -16936 58054
rect -17556 57734 -16936 57818
rect -17556 57498 -17524 57734
rect -17288 57498 -17204 57734
rect -16968 57498 -16936 57734
rect -17556 -15896 -16936 57498
rect -14446 717278 -13826 717310
rect -14446 717042 -14414 717278
rect -14178 717042 -14094 717278
rect -13858 717042 -13826 717278
rect -14446 716958 -13826 717042
rect -14446 716722 -14414 716958
rect -14178 716722 -14094 716958
rect -13858 716722 -13826 716958
rect -14446 666334 -13826 716722
rect -14446 666098 -14414 666334
rect -14178 666098 -14094 666334
rect -13858 666098 -13826 666334
rect -14446 666014 -13826 666098
rect -14446 665778 -14414 666014
rect -14178 665778 -14094 666014
rect -13858 665778 -13826 666014
rect -14446 630334 -13826 665778
rect -14446 630098 -14414 630334
rect -14178 630098 -14094 630334
rect -13858 630098 -13826 630334
rect -14446 630014 -13826 630098
rect -14446 629778 -14414 630014
rect -14178 629778 -14094 630014
rect -13858 629778 -13826 630014
rect -14446 594334 -13826 629778
rect -14446 594098 -14414 594334
rect -14178 594098 -14094 594334
rect -13858 594098 -13826 594334
rect -14446 594014 -13826 594098
rect -14446 593778 -14414 594014
rect -14178 593778 -14094 594014
rect -13858 593778 -13826 594014
rect -14446 558334 -13826 593778
rect -14446 558098 -14414 558334
rect -14178 558098 -14094 558334
rect -13858 558098 -13826 558334
rect -14446 558014 -13826 558098
rect -14446 557778 -14414 558014
rect -14178 557778 -14094 558014
rect -13858 557778 -13826 558014
rect -14446 522334 -13826 557778
rect -14446 522098 -14414 522334
rect -14178 522098 -14094 522334
rect -13858 522098 -13826 522334
rect -14446 522014 -13826 522098
rect -14446 521778 -14414 522014
rect -14178 521778 -14094 522014
rect -13858 521778 -13826 522014
rect -14446 486334 -13826 521778
rect -14446 486098 -14414 486334
rect -14178 486098 -14094 486334
rect -13858 486098 -13826 486334
rect -14446 486014 -13826 486098
rect -14446 485778 -14414 486014
rect -14178 485778 -14094 486014
rect -13858 485778 -13826 486014
rect -14446 450334 -13826 485778
rect -14446 450098 -14414 450334
rect -14178 450098 -14094 450334
rect -13858 450098 -13826 450334
rect -14446 450014 -13826 450098
rect -14446 449778 -14414 450014
rect -14178 449778 -14094 450014
rect -13858 449778 -13826 450014
rect -14446 414334 -13826 449778
rect -14446 414098 -14414 414334
rect -14178 414098 -14094 414334
rect -13858 414098 -13826 414334
rect -14446 414014 -13826 414098
rect -14446 413778 -14414 414014
rect -14178 413778 -14094 414014
rect -13858 413778 -13826 414014
rect -14446 378334 -13826 413778
rect -14446 378098 -14414 378334
rect -14178 378098 -14094 378334
rect -13858 378098 -13826 378334
rect -14446 378014 -13826 378098
rect -14446 377778 -14414 378014
rect -14178 377778 -14094 378014
rect -13858 377778 -13826 378014
rect -14446 342334 -13826 377778
rect -14446 342098 -14414 342334
rect -14178 342098 -14094 342334
rect -13858 342098 -13826 342334
rect -14446 342014 -13826 342098
rect -14446 341778 -14414 342014
rect -14178 341778 -14094 342014
rect -13858 341778 -13826 342014
rect -14446 306334 -13826 341778
rect -14446 306098 -14414 306334
rect -14178 306098 -14094 306334
rect -13858 306098 -13826 306334
rect -14446 306014 -13826 306098
rect -14446 305778 -14414 306014
rect -14178 305778 -14094 306014
rect -13858 305778 -13826 306014
rect -14446 270334 -13826 305778
rect -14446 270098 -14414 270334
rect -14178 270098 -14094 270334
rect -13858 270098 -13826 270334
rect -14446 270014 -13826 270098
rect -14446 269778 -14414 270014
rect -14178 269778 -14094 270014
rect -13858 269778 -13826 270014
rect -14446 234334 -13826 269778
rect -14446 234098 -14414 234334
rect -14178 234098 -14094 234334
rect -13858 234098 -13826 234334
rect -14446 234014 -13826 234098
rect -14446 233778 -14414 234014
rect -14178 233778 -14094 234014
rect -13858 233778 -13826 234014
rect -14446 198334 -13826 233778
rect -14446 198098 -14414 198334
rect -14178 198098 -14094 198334
rect -13858 198098 -13826 198334
rect -14446 198014 -13826 198098
rect -14446 197778 -14414 198014
rect -14178 197778 -14094 198014
rect -13858 197778 -13826 198014
rect -14446 162334 -13826 197778
rect -14446 162098 -14414 162334
rect -14178 162098 -14094 162334
rect -13858 162098 -13826 162334
rect -14446 162014 -13826 162098
rect -14446 161778 -14414 162014
rect -14178 161778 -14094 162014
rect -13858 161778 -13826 162014
rect -14446 126334 -13826 161778
rect -14446 126098 -14414 126334
rect -14178 126098 -14094 126334
rect -13858 126098 -13826 126334
rect -14446 126014 -13826 126098
rect -14446 125778 -14414 126014
rect -14178 125778 -14094 126014
rect -13858 125778 -13826 126014
rect -14446 90334 -13826 125778
rect -14446 90098 -14414 90334
rect -14178 90098 -14094 90334
rect -13858 90098 -13826 90334
rect -14446 90014 -13826 90098
rect -14446 89778 -14414 90014
rect -14178 89778 -14094 90014
rect -13858 89778 -13826 90014
rect -14446 54334 -13826 89778
rect -14446 54098 -14414 54334
rect -14178 54098 -14094 54334
rect -13858 54098 -13826 54334
rect -14446 54014 -13826 54098
rect -14446 53778 -14414 54014
rect -14178 53778 -14094 54014
rect -13858 53778 -13826 54014
rect -14446 18334 -13826 53778
rect -14446 18098 -14414 18334
rect -14178 18098 -14094 18334
rect -13858 18098 -13826 18334
rect -14446 18014 -13826 18098
rect -14446 17778 -14414 18014
rect -14178 17778 -14094 18014
rect -13858 17778 -13826 18014
rect -14446 -12786 -13826 17778
rect -11336 714168 -10716 714200
rect -11336 713932 -11304 714168
rect -11068 713932 -10984 714168
rect -10748 713932 -10716 714168
rect -11336 713848 -10716 713932
rect -11336 713612 -11304 713848
rect -11068 713612 -10984 713848
rect -10748 713612 -10716 713848
rect -11336 698614 -10716 713612
rect -11336 698378 -11304 698614
rect -11068 698378 -10984 698614
rect -10748 698378 -10716 698614
rect -11336 698294 -10716 698378
rect -11336 698058 -11304 698294
rect -11068 698058 -10984 698294
rect -10748 698058 -10716 698294
rect -11336 662614 -10716 698058
rect -11336 662378 -11304 662614
rect -11068 662378 -10984 662614
rect -10748 662378 -10716 662614
rect -11336 662294 -10716 662378
rect -11336 662058 -11304 662294
rect -11068 662058 -10984 662294
rect -10748 662058 -10716 662294
rect -11336 626614 -10716 662058
rect -11336 626378 -11304 626614
rect -11068 626378 -10984 626614
rect -10748 626378 -10716 626614
rect -11336 626294 -10716 626378
rect -11336 626058 -11304 626294
rect -11068 626058 -10984 626294
rect -10748 626058 -10716 626294
rect -11336 590614 -10716 626058
rect -11336 590378 -11304 590614
rect -11068 590378 -10984 590614
rect -10748 590378 -10716 590614
rect -11336 590294 -10716 590378
rect -11336 590058 -11304 590294
rect -11068 590058 -10984 590294
rect -10748 590058 -10716 590294
rect -11336 554614 -10716 590058
rect -11336 554378 -11304 554614
rect -11068 554378 -10984 554614
rect -10748 554378 -10716 554614
rect -11336 554294 -10716 554378
rect -11336 554058 -11304 554294
rect -11068 554058 -10984 554294
rect -10748 554058 -10716 554294
rect -11336 518614 -10716 554058
rect -11336 518378 -11304 518614
rect -11068 518378 -10984 518614
rect -10748 518378 -10716 518614
rect -11336 518294 -10716 518378
rect -11336 518058 -11304 518294
rect -11068 518058 -10984 518294
rect -10748 518058 -10716 518294
rect -11336 482614 -10716 518058
rect -11336 482378 -11304 482614
rect -11068 482378 -10984 482614
rect -10748 482378 -10716 482614
rect -11336 482294 -10716 482378
rect -11336 482058 -11304 482294
rect -11068 482058 -10984 482294
rect -10748 482058 -10716 482294
rect -11336 446614 -10716 482058
rect -11336 446378 -11304 446614
rect -11068 446378 -10984 446614
rect -10748 446378 -10716 446614
rect -11336 446294 -10716 446378
rect -11336 446058 -11304 446294
rect -11068 446058 -10984 446294
rect -10748 446058 -10716 446294
rect -11336 410614 -10716 446058
rect -11336 410378 -11304 410614
rect -11068 410378 -10984 410614
rect -10748 410378 -10716 410614
rect -11336 410294 -10716 410378
rect -11336 410058 -11304 410294
rect -11068 410058 -10984 410294
rect -10748 410058 -10716 410294
rect -11336 374614 -10716 410058
rect -11336 374378 -11304 374614
rect -11068 374378 -10984 374614
rect -10748 374378 -10716 374614
rect -11336 374294 -10716 374378
rect -11336 374058 -11304 374294
rect -11068 374058 -10984 374294
rect -10748 374058 -10716 374294
rect -11336 338614 -10716 374058
rect -11336 338378 -11304 338614
rect -11068 338378 -10984 338614
rect -10748 338378 -10716 338614
rect -11336 338294 -10716 338378
rect -11336 338058 -11304 338294
rect -11068 338058 -10984 338294
rect -10748 338058 -10716 338294
rect -11336 302614 -10716 338058
rect -11336 302378 -11304 302614
rect -11068 302378 -10984 302614
rect -10748 302378 -10716 302614
rect -11336 302294 -10716 302378
rect -11336 302058 -11304 302294
rect -11068 302058 -10984 302294
rect -10748 302058 -10716 302294
rect -11336 266614 -10716 302058
rect -11336 266378 -11304 266614
rect -11068 266378 -10984 266614
rect -10748 266378 -10716 266614
rect -11336 266294 -10716 266378
rect -11336 266058 -11304 266294
rect -11068 266058 -10984 266294
rect -10748 266058 -10716 266294
rect -11336 230614 -10716 266058
rect -11336 230378 -11304 230614
rect -11068 230378 -10984 230614
rect -10748 230378 -10716 230614
rect -11336 230294 -10716 230378
rect -11336 230058 -11304 230294
rect -11068 230058 -10984 230294
rect -10748 230058 -10716 230294
rect -11336 194614 -10716 230058
rect -11336 194378 -11304 194614
rect -11068 194378 -10984 194614
rect -10748 194378 -10716 194614
rect -11336 194294 -10716 194378
rect -11336 194058 -11304 194294
rect -11068 194058 -10984 194294
rect -10748 194058 -10716 194294
rect -11336 158614 -10716 194058
rect -11336 158378 -11304 158614
rect -11068 158378 -10984 158614
rect -10748 158378 -10716 158614
rect -11336 158294 -10716 158378
rect -11336 158058 -11304 158294
rect -11068 158058 -10984 158294
rect -10748 158058 -10716 158294
rect -11336 122614 -10716 158058
rect -11336 122378 -11304 122614
rect -11068 122378 -10984 122614
rect -10748 122378 -10716 122614
rect -11336 122294 -10716 122378
rect -11336 122058 -11304 122294
rect -11068 122058 -10984 122294
rect -10748 122058 -10716 122294
rect -11336 86614 -10716 122058
rect -11336 86378 -11304 86614
rect -11068 86378 -10984 86614
rect -10748 86378 -10716 86614
rect -11336 86294 -10716 86378
rect -11336 86058 -11304 86294
rect -11068 86058 -10984 86294
rect -10748 86058 -10716 86294
rect -11336 50614 -10716 86058
rect -11336 50378 -11304 50614
rect -11068 50378 -10984 50614
rect -10748 50378 -10716 50614
rect -11336 50294 -10716 50378
rect -11336 50058 -11304 50294
rect -11068 50058 -10984 50294
rect -10748 50058 -10716 50294
rect -11336 14614 -10716 50058
rect -11336 14378 -11304 14614
rect -11068 14378 -10984 14614
rect -10748 14378 -10716 14614
rect -11336 14294 -10716 14378
rect -11336 14058 -11304 14294
rect -11068 14058 -10984 14294
rect -10748 14058 -10716 14294
rect -11336 -9676 -10716 14058
rect -8226 711058 -7606 711090
rect -8226 710822 -8194 711058
rect -7958 710822 -7874 711058
rect -7638 710822 -7606 711058
rect -8226 710738 -7606 710822
rect -8226 710502 -8194 710738
rect -7958 710502 -7874 710738
rect -7638 710502 -7606 710738
rect -8226 694894 -7606 710502
rect -8226 694658 -8194 694894
rect -7958 694658 -7874 694894
rect -7638 694658 -7606 694894
rect -8226 694574 -7606 694658
rect -8226 694338 -8194 694574
rect -7958 694338 -7874 694574
rect -7638 694338 -7606 694574
rect -8226 658894 -7606 694338
rect -8226 658658 -8194 658894
rect -7958 658658 -7874 658894
rect -7638 658658 -7606 658894
rect -8226 658574 -7606 658658
rect -8226 658338 -8194 658574
rect -7958 658338 -7874 658574
rect -7638 658338 -7606 658574
rect -8226 622894 -7606 658338
rect -8226 622658 -8194 622894
rect -7958 622658 -7874 622894
rect -7638 622658 -7606 622894
rect -8226 622574 -7606 622658
rect -8226 622338 -8194 622574
rect -7958 622338 -7874 622574
rect -7638 622338 -7606 622574
rect -8226 586894 -7606 622338
rect -8226 586658 -8194 586894
rect -7958 586658 -7874 586894
rect -7638 586658 -7606 586894
rect -8226 586574 -7606 586658
rect -8226 586338 -8194 586574
rect -7958 586338 -7874 586574
rect -7638 586338 -7606 586574
rect -8226 550894 -7606 586338
rect -8226 550658 -8194 550894
rect -7958 550658 -7874 550894
rect -7638 550658 -7606 550894
rect -8226 550574 -7606 550658
rect -8226 550338 -8194 550574
rect -7958 550338 -7874 550574
rect -7638 550338 -7606 550574
rect -8226 514894 -7606 550338
rect -8226 514658 -8194 514894
rect -7958 514658 -7874 514894
rect -7638 514658 -7606 514894
rect -8226 514574 -7606 514658
rect -8226 514338 -8194 514574
rect -7958 514338 -7874 514574
rect -7638 514338 -7606 514574
rect -8226 478894 -7606 514338
rect -8226 478658 -8194 478894
rect -7958 478658 -7874 478894
rect -7638 478658 -7606 478894
rect -8226 478574 -7606 478658
rect -8226 478338 -8194 478574
rect -7958 478338 -7874 478574
rect -7638 478338 -7606 478574
rect -8226 442894 -7606 478338
rect -8226 442658 -8194 442894
rect -7958 442658 -7874 442894
rect -7638 442658 -7606 442894
rect -8226 442574 -7606 442658
rect -8226 442338 -8194 442574
rect -7958 442338 -7874 442574
rect -7638 442338 -7606 442574
rect -8226 406894 -7606 442338
rect -8226 406658 -8194 406894
rect -7958 406658 -7874 406894
rect -7638 406658 -7606 406894
rect -8226 406574 -7606 406658
rect -8226 406338 -8194 406574
rect -7958 406338 -7874 406574
rect -7638 406338 -7606 406574
rect -8226 370894 -7606 406338
rect -8226 370658 -8194 370894
rect -7958 370658 -7874 370894
rect -7638 370658 -7606 370894
rect -8226 370574 -7606 370658
rect -8226 370338 -8194 370574
rect -7958 370338 -7874 370574
rect -7638 370338 -7606 370574
rect -8226 334894 -7606 370338
rect -8226 334658 -8194 334894
rect -7958 334658 -7874 334894
rect -7638 334658 -7606 334894
rect -8226 334574 -7606 334658
rect -8226 334338 -8194 334574
rect -7958 334338 -7874 334574
rect -7638 334338 -7606 334574
rect -8226 298894 -7606 334338
rect -8226 298658 -8194 298894
rect -7958 298658 -7874 298894
rect -7638 298658 -7606 298894
rect -8226 298574 -7606 298658
rect -8226 298338 -8194 298574
rect -7958 298338 -7874 298574
rect -7638 298338 -7606 298574
rect -8226 262894 -7606 298338
rect -8226 262658 -8194 262894
rect -7958 262658 -7874 262894
rect -7638 262658 -7606 262894
rect -8226 262574 -7606 262658
rect -8226 262338 -8194 262574
rect -7958 262338 -7874 262574
rect -7638 262338 -7606 262574
rect -8226 226894 -7606 262338
rect -8226 226658 -8194 226894
rect -7958 226658 -7874 226894
rect -7638 226658 -7606 226894
rect -8226 226574 -7606 226658
rect -8226 226338 -8194 226574
rect -7958 226338 -7874 226574
rect -7638 226338 -7606 226574
rect -8226 190894 -7606 226338
rect -8226 190658 -8194 190894
rect -7958 190658 -7874 190894
rect -7638 190658 -7606 190894
rect -8226 190574 -7606 190658
rect -8226 190338 -8194 190574
rect -7958 190338 -7874 190574
rect -7638 190338 -7606 190574
rect -8226 154894 -7606 190338
rect -8226 154658 -8194 154894
rect -7958 154658 -7874 154894
rect -7638 154658 -7606 154894
rect -8226 154574 -7606 154658
rect -8226 154338 -8194 154574
rect -7958 154338 -7874 154574
rect -7638 154338 -7606 154574
rect -8226 118894 -7606 154338
rect -8226 118658 -8194 118894
rect -7958 118658 -7874 118894
rect -7638 118658 -7606 118894
rect -8226 118574 -7606 118658
rect -8226 118338 -8194 118574
rect -7958 118338 -7874 118574
rect -7638 118338 -7606 118574
rect -8226 82894 -7606 118338
rect -8226 82658 -8194 82894
rect -7958 82658 -7874 82894
rect -7638 82658 -7606 82894
rect -8226 82574 -7606 82658
rect -8226 82338 -8194 82574
rect -7958 82338 -7874 82574
rect -7638 82338 -7606 82574
rect -8226 46894 -7606 82338
rect -8226 46658 -8194 46894
rect -7958 46658 -7874 46894
rect -7638 46658 -7606 46894
rect -8226 46574 -7606 46658
rect -8226 46338 -8194 46574
rect -7958 46338 -7874 46574
rect -7638 46338 -7606 46574
rect -8226 10894 -7606 46338
rect -8226 10658 -8194 10894
rect -7958 10658 -7874 10894
rect -7638 10658 -7606 10894
rect -8226 10574 -7606 10658
rect -8226 10338 -8194 10574
rect -7958 10338 -7874 10574
rect -7638 10338 -7606 10574
rect -8226 -6566 -7606 10338
rect -5116 707948 -4496 707980
rect -5116 707712 -5084 707948
rect -4848 707712 -4764 707948
rect -4528 707712 -4496 707948
rect -5116 707628 -4496 707712
rect -5116 707392 -5084 707628
rect -4848 707392 -4764 707628
rect -4528 707392 -4496 707628
rect -5116 691174 -4496 707392
rect 581514 707948 582134 726640
rect 607080 726608 607700 726640
rect 607080 726372 607112 726608
rect 607348 726372 607432 726608
rect 607668 726372 607700 726608
rect 607080 726288 607700 726372
rect 607080 726052 607112 726288
rect 607348 726052 607432 726288
rect 607668 726052 607700 726288
rect 603970 723498 604590 723530
rect 603970 723262 604002 723498
rect 604238 723262 604322 723498
rect 604558 723262 604590 723498
rect 603970 723178 604590 723262
rect 603970 722942 604002 723178
rect 604238 722942 604322 723178
rect 604558 722942 604590 723178
rect 600860 720388 601480 720420
rect 600860 720152 600892 720388
rect 601128 720152 601212 720388
rect 601448 720152 601480 720388
rect 600860 720068 601480 720152
rect 600860 719832 600892 720068
rect 601128 719832 601212 720068
rect 601448 719832 601480 720068
rect 597750 717278 598370 717310
rect 597750 717042 597782 717278
rect 598018 717042 598102 717278
rect 598338 717042 598370 717278
rect 597750 716958 598370 717042
rect 597750 716722 597782 716958
rect 598018 716722 598102 716958
rect 598338 716722 598370 716958
rect 594640 714168 595260 714200
rect 594640 713932 594672 714168
rect 594908 713932 594992 714168
rect 595228 713932 595260 714168
rect 594640 713848 595260 713932
rect 594640 713612 594672 713848
rect 594908 713612 594992 713848
rect 595228 713612 595260 713848
rect 591530 711058 592150 711090
rect 591530 710822 591562 711058
rect 591798 710822 591882 711058
rect 592118 710822 592150 711058
rect 591530 710738 592150 710822
rect 591530 710502 591562 710738
rect 591798 710502 591882 710738
rect 592118 710502 592150 710738
rect 581514 707712 581546 707948
rect 581782 707712 581866 707948
rect 582102 707712 582134 707948
rect 581514 707628 582134 707712
rect 581514 707392 581546 707628
rect 581782 707392 581866 707628
rect 582102 707392 582134 707628
rect -5116 690938 -5084 691174
rect -4848 690938 -4764 691174
rect -4528 690938 -4496 691174
rect -5116 690854 -4496 690938
rect -5116 690618 -5084 690854
rect -4848 690618 -4764 690854
rect -4528 690618 -4496 690854
rect -5116 655174 -4496 690618
rect -5116 654938 -5084 655174
rect -4848 654938 -4764 655174
rect -4528 654938 -4496 655174
rect -5116 654854 -4496 654938
rect -5116 654618 -5084 654854
rect -4848 654618 -4764 654854
rect -4528 654618 -4496 654854
rect -5116 619174 -4496 654618
rect -5116 618938 -5084 619174
rect -4848 618938 -4764 619174
rect -4528 618938 -4496 619174
rect -5116 618854 -4496 618938
rect -5116 618618 -5084 618854
rect -4848 618618 -4764 618854
rect -4528 618618 -4496 618854
rect -5116 583174 -4496 618618
rect -5116 582938 -5084 583174
rect -4848 582938 -4764 583174
rect -4528 582938 -4496 583174
rect -5116 582854 -4496 582938
rect -5116 582618 -5084 582854
rect -4848 582618 -4764 582854
rect -4528 582618 -4496 582854
rect -5116 547174 -4496 582618
rect -5116 546938 -5084 547174
rect -4848 546938 -4764 547174
rect -4528 546938 -4496 547174
rect -5116 546854 -4496 546938
rect -5116 546618 -5084 546854
rect -4848 546618 -4764 546854
rect -4528 546618 -4496 546854
rect -5116 511174 -4496 546618
rect -5116 510938 -5084 511174
rect -4848 510938 -4764 511174
rect -4528 510938 -4496 511174
rect -5116 510854 -4496 510938
rect -5116 510618 -5084 510854
rect -4848 510618 -4764 510854
rect -4528 510618 -4496 510854
rect -5116 475174 -4496 510618
rect -5116 474938 -5084 475174
rect -4848 474938 -4764 475174
rect -4528 474938 -4496 475174
rect -5116 474854 -4496 474938
rect -5116 474618 -5084 474854
rect -4848 474618 -4764 474854
rect -4528 474618 -4496 474854
rect -5116 439174 -4496 474618
rect -5116 438938 -5084 439174
rect -4848 438938 -4764 439174
rect -4528 438938 -4496 439174
rect -5116 438854 -4496 438938
rect -5116 438618 -5084 438854
rect -4848 438618 -4764 438854
rect -4528 438618 -4496 438854
rect -5116 403174 -4496 438618
rect -5116 402938 -5084 403174
rect -4848 402938 -4764 403174
rect -4528 402938 -4496 403174
rect -5116 402854 -4496 402938
rect -5116 402618 -5084 402854
rect -4848 402618 -4764 402854
rect -4528 402618 -4496 402854
rect -5116 367174 -4496 402618
rect -5116 366938 -5084 367174
rect -4848 366938 -4764 367174
rect -4528 366938 -4496 367174
rect -5116 366854 -4496 366938
rect -5116 366618 -5084 366854
rect -4848 366618 -4764 366854
rect -4528 366618 -4496 366854
rect -5116 331174 -4496 366618
rect -5116 330938 -5084 331174
rect -4848 330938 -4764 331174
rect -4528 330938 -4496 331174
rect -5116 330854 -4496 330938
rect -5116 330618 -5084 330854
rect -4848 330618 -4764 330854
rect -4528 330618 -4496 330854
rect -5116 295174 -4496 330618
rect -5116 294938 -5084 295174
rect -4848 294938 -4764 295174
rect -4528 294938 -4496 295174
rect -5116 294854 -4496 294938
rect -5116 294618 -5084 294854
rect -4848 294618 -4764 294854
rect -4528 294618 -4496 294854
rect -5116 259174 -4496 294618
rect -5116 258938 -5084 259174
rect -4848 258938 -4764 259174
rect -4528 258938 -4496 259174
rect -5116 258854 -4496 258938
rect -5116 258618 -5084 258854
rect -4848 258618 -4764 258854
rect -4528 258618 -4496 258854
rect -5116 223174 -4496 258618
rect -5116 222938 -5084 223174
rect -4848 222938 -4764 223174
rect -4528 222938 -4496 223174
rect -5116 222854 -4496 222938
rect -5116 222618 -5084 222854
rect -4848 222618 -4764 222854
rect -4528 222618 -4496 222854
rect -5116 187174 -4496 222618
rect -5116 186938 -5084 187174
rect -4848 186938 -4764 187174
rect -4528 186938 -4496 187174
rect -5116 186854 -4496 186938
rect -5116 186618 -5084 186854
rect -4848 186618 -4764 186854
rect -4528 186618 -4496 186854
rect -5116 151174 -4496 186618
rect -5116 150938 -5084 151174
rect -4848 150938 -4764 151174
rect -4528 150938 -4496 151174
rect -5116 150854 -4496 150938
rect -5116 150618 -5084 150854
rect -4848 150618 -4764 150854
rect -4528 150618 -4496 150854
rect -5116 115174 -4496 150618
rect -5116 114938 -5084 115174
rect -4848 114938 -4764 115174
rect -4528 114938 -4496 115174
rect -5116 114854 -4496 114938
rect -5116 114618 -5084 114854
rect -4848 114618 -4764 114854
rect -4528 114618 -4496 114854
rect -5116 79174 -4496 114618
rect -5116 78938 -5084 79174
rect -4848 78938 -4764 79174
rect -4528 78938 -4496 79174
rect -5116 78854 -4496 78938
rect -5116 78618 -5084 78854
rect -4848 78618 -4764 78854
rect -4528 78618 -4496 78854
rect -5116 43174 -4496 78618
rect -5116 42938 -5084 43174
rect -4848 42938 -4764 43174
rect -4528 42938 -4496 43174
rect -5116 42854 -4496 42938
rect -5116 42618 -5084 42854
rect -4848 42618 -4764 42854
rect -4528 42618 -4496 42854
rect -5116 7174 -4496 42618
rect -5116 6938 -5084 7174
rect -4848 6938 -4764 7174
rect -4528 6938 -4496 7174
rect -5116 6854 -4496 6938
rect -5116 6618 -5084 6854
rect -4848 6618 -4764 6854
rect -4528 6618 -4496 6854
rect -5116 -3456 -4496 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect 7844 693480 7876 693716
rect 8112 693480 8196 693716
rect 8432 693480 8464 693716
rect 7844 693396 8464 693480
rect 7844 693160 7876 693396
rect 8112 693160 8196 693396
rect 8432 693160 8464 693396
rect 38000 693480 38032 693716
rect 38268 693480 38352 693716
rect 38588 693480 38620 693716
rect 38000 693396 38620 693480
rect 38000 693160 38032 693396
rect 38268 693160 38352 693396
rect 38588 693160 38620 693396
rect 74000 693480 74032 693716
rect 74268 693480 74352 693716
rect 74588 693480 74620 693716
rect 74000 693396 74620 693480
rect 74000 693160 74032 693396
rect 74268 693160 74352 693396
rect 74588 693160 74620 693396
rect 110000 693480 110032 693716
rect 110268 693480 110352 693716
rect 110588 693480 110620 693716
rect 110000 693396 110620 693480
rect 110000 693160 110032 693396
rect 110268 693160 110352 693396
rect 110588 693160 110620 693396
rect 146000 693480 146032 693716
rect 146268 693480 146352 693716
rect 146588 693480 146620 693716
rect 146000 693396 146620 693480
rect 146000 693160 146032 693396
rect 146268 693160 146352 693396
rect 146588 693160 146620 693396
rect 182000 693480 182032 693716
rect 182268 693480 182352 693716
rect 182588 693480 182620 693716
rect 182000 693396 182620 693480
rect 182000 693160 182032 693396
rect 182268 693160 182352 693396
rect 182588 693160 182620 693396
rect 218000 693480 218032 693716
rect 218268 693480 218352 693716
rect 218588 693480 218620 693716
rect 218000 693396 218620 693480
rect 218000 693160 218032 693396
rect 218268 693160 218352 693396
rect 218588 693160 218620 693396
rect 254000 693480 254032 693716
rect 254268 693480 254352 693716
rect 254588 693480 254620 693716
rect 254000 693396 254620 693480
rect 254000 693160 254032 693396
rect 254268 693160 254352 693396
rect 254588 693160 254620 693396
rect 290000 693480 290032 693716
rect 290268 693480 290352 693716
rect 290588 693480 290620 693716
rect 290000 693396 290620 693480
rect 290000 693160 290032 693396
rect 290268 693160 290352 693396
rect 290588 693160 290620 693396
rect 326000 693480 326032 693716
rect 326268 693480 326352 693716
rect 326588 693480 326620 693716
rect 326000 693396 326620 693480
rect 326000 693160 326032 693396
rect 326268 693160 326352 693396
rect 326588 693160 326620 693396
rect 362000 693480 362032 693716
rect 362268 693480 362352 693716
rect 362588 693480 362620 693716
rect 362000 693396 362620 693480
rect 362000 693160 362032 693396
rect 362268 693160 362352 693396
rect 362588 693160 362620 693396
rect 398000 693480 398032 693716
rect 398268 693480 398352 693716
rect 398588 693480 398620 693716
rect 398000 693396 398620 693480
rect 398000 693160 398032 693396
rect 398268 693160 398352 693396
rect 398588 693160 398620 693396
rect 434000 693480 434032 693716
rect 434268 693480 434352 693716
rect 434588 693480 434620 693716
rect 434000 693396 434620 693480
rect 434000 693160 434032 693396
rect 434268 693160 434352 693396
rect 434588 693160 434620 693396
rect 470000 693480 470032 693716
rect 470268 693480 470352 693716
rect 470588 693480 470620 693716
rect 470000 693396 470620 693480
rect 470000 693160 470032 693396
rect 470268 693160 470352 693396
rect 470588 693160 470620 693396
rect 506000 693480 506032 693716
rect 506268 693480 506352 693716
rect 506588 693480 506620 693716
rect 506000 693396 506620 693480
rect 506000 693160 506032 693396
rect 506268 693160 506352 693396
rect 506588 693160 506620 693396
rect 542000 693480 542032 693716
rect 542268 693480 542352 693716
rect 542588 693480 542620 693716
rect 542000 693396 542620 693480
rect 542000 693160 542032 693396
rect 542268 693160 542352 693396
rect 542588 693160 542620 693396
rect 571500 693480 571532 693716
rect 571768 693480 571852 693716
rect 572088 693480 572120 693716
rect 571500 693396 572120 693480
rect 571500 693160 571532 693396
rect 571768 693160 571852 693396
rect 572088 693160 572120 693396
rect 9084 692240 9116 692476
rect 9352 692240 9436 692476
rect 9672 692240 9704 692476
rect 9084 692156 9704 692240
rect 9084 691920 9116 692156
rect 9352 691920 9436 692156
rect 9672 691920 9704 692156
rect 56620 692240 56652 692476
rect 56888 692240 56972 692476
rect 57208 692240 57240 692476
rect 56620 692156 57240 692240
rect 56620 691920 56652 692156
rect 56888 691920 56972 692156
rect 57208 691920 57240 692156
rect 92620 692240 92652 692476
rect 92888 692240 92972 692476
rect 93208 692240 93240 692476
rect 92620 692156 93240 692240
rect 92620 691920 92652 692156
rect 92888 691920 92972 692156
rect 93208 691920 93240 692156
rect 128620 692240 128652 692476
rect 128888 692240 128972 692476
rect 129208 692240 129240 692476
rect 128620 692156 129240 692240
rect 128620 691920 128652 692156
rect 128888 691920 128972 692156
rect 129208 691920 129240 692156
rect 164620 692240 164652 692476
rect 164888 692240 164972 692476
rect 165208 692240 165240 692476
rect 164620 692156 165240 692240
rect 164620 691920 164652 692156
rect 164888 691920 164972 692156
rect 165208 691920 165240 692156
rect 200620 692240 200652 692476
rect 200888 692240 200972 692476
rect 201208 692240 201240 692476
rect 200620 692156 201240 692240
rect 200620 691920 200652 692156
rect 200888 691920 200972 692156
rect 201208 691920 201240 692156
rect 236620 692240 236652 692476
rect 236888 692240 236972 692476
rect 237208 692240 237240 692476
rect 236620 692156 237240 692240
rect 236620 691920 236652 692156
rect 236888 691920 236972 692156
rect 237208 691920 237240 692156
rect 272620 692240 272652 692476
rect 272888 692240 272972 692476
rect 273208 692240 273240 692476
rect 272620 692156 273240 692240
rect 272620 691920 272652 692156
rect 272888 691920 272972 692156
rect 273208 691920 273240 692156
rect 308620 692240 308652 692476
rect 308888 692240 308972 692476
rect 309208 692240 309240 692476
rect 308620 692156 309240 692240
rect 308620 691920 308652 692156
rect 308888 691920 308972 692156
rect 309208 691920 309240 692156
rect 344620 692240 344652 692476
rect 344888 692240 344972 692476
rect 345208 692240 345240 692476
rect 344620 692156 345240 692240
rect 344620 691920 344652 692156
rect 344888 691920 344972 692156
rect 345208 691920 345240 692156
rect 380620 692240 380652 692476
rect 380888 692240 380972 692476
rect 381208 692240 381240 692476
rect 380620 692156 381240 692240
rect 380620 691920 380652 692156
rect 380888 691920 380972 692156
rect 381208 691920 381240 692156
rect 416620 692240 416652 692476
rect 416888 692240 416972 692476
rect 417208 692240 417240 692476
rect 416620 692156 417240 692240
rect 416620 691920 416652 692156
rect 416888 691920 416972 692156
rect 417208 691920 417240 692156
rect 452620 692240 452652 692476
rect 452888 692240 452972 692476
rect 453208 692240 453240 692476
rect 452620 692156 453240 692240
rect 452620 691920 452652 692156
rect 452888 691920 452972 692156
rect 453208 691920 453240 692156
rect 488620 692240 488652 692476
rect 488888 692240 488972 692476
rect 489208 692240 489240 692476
rect 488620 692156 489240 692240
rect 488620 691920 488652 692156
rect 488888 691920 488972 692156
rect 489208 691920 489240 692156
rect 524620 692240 524652 692476
rect 524888 692240 524972 692476
rect 525208 692240 525240 692476
rect 524620 692156 525240 692240
rect 524620 691920 524652 692156
rect 524888 691920 524972 692156
rect 525208 691920 525240 692156
rect 560620 692240 560652 692476
rect 560888 692240 560972 692476
rect 561208 692240 561240 692476
rect 560620 692156 561240 692240
rect 560620 691920 560652 692156
rect 560888 691920 560972 692156
rect 561208 691920 561240 692156
rect 570260 692240 570292 692476
rect 570528 692240 570612 692476
rect 570848 692240 570880 692476
rect 570260 692156 570880 692240
rect 570260 691920 570292 692156
rect 570528 691920 570612 692156
rect 570848 691920 570880 692156
rect 581514 691174 582134 707392
rect 588420 707948 589040 707980
rect 588420 707712 588452 707948
rect 588688 707712 588772 707948
rect 589008 707712 589040 707948
rect 588420 707628 589040 707712
rect 588420 707392 588452 707628
rect 588688 707392 588772 707628
rect 589008 707392 589040 707628
rect 7844 690938 7876 691174
rect 8112 690938 8196 691174
rect 8432 690938 8464 691174
rect 7844 690854 8464 690938
rect 7844 690618 7876 690854
rect 8112 690618 8196 690854
rect 8432 690618 8464 690854
rect 38000 690938 38032 691174
rect 38268 690938 38352 691174
rect 38588 690938 38620 691174
rect 38000 690854 38620 690938
rect 38000 690618 38032 690854
rect 38268 690618 38352 690854
rect 38588 690618 38620 690854
rect 74000 690938 74032 691174
rect 74268 690938 74352 691174
rect 74588 690938 74620 691174
rect 74000 690854 74620 690938
rect 74000 690618 74032 690854
rect 74268 690618 74352 690854
rect 74588 690618 74620 690854
rect 110000 690938 110032 691174
rect 110268 690938 110352 691174
rect 110588 690938 110620 691174
rect 110000 690854 110620 690938
rect 110000 690618 110032 690854
rect 110268 690618 110352 690854
rect 110588 690618 110620 690854
rect 146000 690938 146032 691174
rect 146268 690938 146352 691174
rect 146588 690938 146620 691174
rect 146000 690854 146620 690938
rect 146000 690618 146032 690854
rect 146268 690618 146352 690854
rect 146588 690618 146620 690854
rect 182000 690938 182032 691174
rect 182268 690938 182352 691174
rect 182588 690938 182620 691174
rect 182000 690854 182620 690938
rect 182000 690618 182032 690854
rect 182268 690618 182352 690854
rect 182588 690618 182620 690854
rect 218000 690938 218032 691174
rect 218268 690938 218352 691174
rect 218588 690938 218620 691174
rect 218000 690854 218620 690938
rect 218000 690618 218032 690854
rect 218268 690618 218352 690854
rect 218588 690618 218620 690854
rect 254000 690938 254032 691174
rect 254268 690938 254352 691174
rect 254588 690938 254620 691174
rect 254000 690854 254620 690938
rect 254000 690618 254032 690854
rect 254268 690618 254352 690854
rect 254588 690618 254620 690854
rect 290000 690938 290032 691174
rect 290268 690938 290352 691174
rect 290588 690938 290620 691174
rect 290000 690854 290620 690938
rect 290000 690618 290032 690854
rect 290268 690618 290352 690854
rect 290588 690618 290620 690854
rect 326000 690938 326032 691174
rect 326268 690938 326352 691174
rect 326588 690938 326620 691174
rect 326000 690854 326620 690938
rect 326000 690618 326032 690854
rect 326268 690618 326352 690854
rect 326588 690618 326620 690854
rect 362000 690938 362032 691174
rect 362268 690938 362352 691174
rect 362588 690938 362620 691174
rect 362000 690854 362620 690938
rect 362000 690618 362032 690854
rect 362268 690618 362352 690854
rect 362588 690618 362620 690854
rect 398000 690938 398032 691174
rect 398268 690938 398352 691174
rect 398588 690938 398620 691174
rect 398000 690854 398620 690938
rect 398000 690618 398032 690854
rect 398268 690618 398352 690854
rect 398588 690618 398620 690854
rect 434000 690938 434032 691174
rect 434268 690938 434352 691174
rect 434588 690938 434620 691174
rect 434000 690854 434620 690938
rect 434000 690618 434032 690854
rect 434268 690618 434352 690854
rect 434588 690618 434620 690854
rect 470000 690938 470032 691174
rect 470268 690938 470352 691174
rect 470588 690938 470620 691174
rect 470000 690854 470620 690938
rect 470000 690618 470032 690854
rect 470268 690618 470352 690854
rect 470588 690618 470620 690854
rect 506000 690938 506032 691174
rect 506268 690938 506352 691174
rect 506588 690938 506620 691174
rect 506000 690854 506620 690938
rect 506000 690618 506032 690854
rect 506268 690618 506352 690854
rect 506588 690618 506620 690854
rect 542000 690938 542032 691174
rect 542268 690938 542352 691174
rect 542588 690938 542620 691174
rect 542000 690854 542620 690938
rect 542000 690618 542032 690854
rect 542268 690618 542352 690854
rect 542588 690618 542620 690854
rect 571500 690938 571532 691174
rect 571768 690938 571852 691174
rect 572088 690938 572120 691174
rect 571500 690854 572120 690938
rect 571500 690618 571532 690854
rect 571768 690618 571852 690854
rect 572088 690618 572120 690854
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect 9084 687218 9116 687454
rect 9352 687218 9436 687454
rect 9672 687218 9704 687454
rect 9084 687134 9704 687218
rect 9084 686898 9116 687134
rect 9352 686898 9436 687134
rect 9672 686898 9704 687134
rect 56620 687218 56652 687454
rect 56888 687218 56972 687454
rect 57208 687218 57240 687454
rect 56620 687134 57240 687218
rect 56620 686898 56652 687134
rect 56888 686898 56972 687134
rect 57208 686898 57240 687134
rect 92620 687218 92652 687454
rect 92888 687218 92972 687454
rect 93208 687218 93240 687454
rect 92620 687134 93240 687218
rect 92620 686898 92652 687134
rect 92888 686898 92972 687134
rect 93208 686898 93240 687134
rect 128620 687218 128652 687454
rect 128888 687218 128972 687454
rect 129208 687218 129240 687454
rect 128620 687134 129240 687218
rect 128620 686898 128652 687134
rect 128888 686898 128972 687134
rect 129208 686898 129240 687134
rect 164620 687218 164652 687454
rect 164888 687218 164972 687454
rect 165208 687218 165240 687454
rect 164620 687134 165240 687218
rect 164620 686898 164652 687134
rect 164888 686898 164972 687134
rect 165208 686898 165240 687134
rect 200620 687218 200652 687454
rect 200888 687218 200972 687454
rect 201208 687218 201240 687454
rect 200620 687134 201240 687218
rect 200620 686898 200652 687134
rect 200888 686898 200972 687134
rect 201208 686898 201240 687134
rect 236620 687218 236652 687454
rect 236888 687218 236972 687454
rect 237208 687218 237240 687454
rect 236620 687134 237240 687218
rect 236620 686898 236652 687134
rect 236888 686898 236972 687134
rect 237208 686898 237240 687134
rect 272620 687218 272652 687454
rect 272888 687218 272972 687454
rect 273208 687218 273240 687454
rect 272620 687134 273240 687218
rect 272620 686898 272652 687134
rect 272888 686898 272972 687134
rect 273208 686898 273240 687134
rect 308620 687218 308652 687454
rect 308888 687218 308972 687454
rect 309208 687218 309240 687454
rect 308620 687134 309240 687218
rect 308620 686898 308652 687134
rect 308888 686898 308972 687134
rect 309208 686898 309240 687134
rect 344620 687218 344652 687454
rect 344888 687218 344972 687454
rect 345208 687218 345240 687454
rect 344620 687134 345240 687218
rect 344620 686898 344652 687134
rect 344888 686898 344972 687134
rect 345208 686898 345240 687134
rect 380620 687218 380652 687454
rect 380888 687218 380972 687454
rect 381208 687218 381240 687454
rect 380620 687134 381240 687218
rect 380620 686898 380652 687134
rect 380888 686898 380972 687134
rect 381208 686898 381240 687134
rect 416620 687218 416652 687454
rect 416888 687218 416972 687454
rect 417208 687218 417240 687454
rect 416620 687134 417240 687218
rect 416620 686898 416652 687134
rect 416888 686898 416972 687134
rect 417208 686898 417240 687134
rect 452620 687218 452652 687454
rect 452888 687218 452972 687454
rect 453208 687218 453240 687454
rect 452620 687134 453240 687218
rect 452620 686898 452652 687134
rect 452888 686898 452972 687134
rect 453208 686898 453240 687134
rect 488620 687218 488652 687454
rect 488888 687218 488972 687454
rect 489208 687218 489240 687454
rect 488620 687134 489240 687218
rect 488620 686898 488652 687134
rect 488888 686898 488972 687134
rect 489208 686898 489240 687134
rect 524620 687218 524652 687454
rect 524888 687218 524972 687454
rect 525208 687218 525240 687454
rect 524620 687134 525240 687218
rect 524620 686898 524652 687134
rect 524888 686898 524972 687134
rect 525208 686898 525240 687134
rect 560620 687218 560652 687454
rect 560888 687218 560972 687454
rect 561208 687218 561240 687454
rect 560620 687134 561240 687218
rect 560620 686898 560652 687134
rect 560888 686898 560972 687134
rect 561208 686898 561240 687134
rect 570260 687218 570292 687454
rect 570528 687218 570612 687454
rect 570848 687218 570880 687454
rect 570260 687134 570880 687218
rect 570260 686898 570292 687134
rect 570528 686898 570612 687134
rect 570848 686898 570880 687134
rect -2006 651454 -1386 686898
rect 581514 655174 582134 690618
rect 7844 654938 7876 655174
rect 8112 654938 8196 655174
rect 8432 654938 8464 655174
rect 7844 654854 8464 654938
rect 7844 654618 7876 654854
rect 8112 654618 8196 654854
rect 8432 654618 8464 654854
rect 38000 654938 38032 655174
rect 38268 654938 38352 655174
rect 38588 654938 38620 655174
rect 38000 654854 38620 654938
rect 38000 654618 38032 654854
rect 38268 654618 38352 654854
rect 38588 654618 38620 654854
rect 74000 654938 74032 655174
rect 74268 654938 74352 655174
rect 74588 654938 74620 655174
rect 74000 654854 74620 654938
rect 74000 654618 74032 654854
rect 74268 654618 74352 654854
rect 74588 654618 74620 654854
rect 110000 654938 110032 655174
rect 110268 654938 110352 655174
rect 110588 654938 110620 655174
rect 110000 654854 110620 654938
rect 110000 654618 110032 654854
rect 110268 654618 110352 654854
rect 110588 654618 110620 654854
rect 146000 654938 146032 655174
rect 146268 654938 146352 655174
rect 146588 654938 146620 655174
rect 146000 654854 146620 654938
rect 146000 654618 146032 654854
rect 146268 654618 146352 654854
rect 146588 654618 146620 654854
rect 182000 654938 182032 655174
rect 182268 654938 182352 655174
rect 182588 654938 182620 655174
rect 182000 654854 182620 654938
rect 182000 654618 182032 654854
rect 182268 654618 182352 654854
rect 182588 654618 182620 654854
rect 218000 654938 218032 655174
rect 218268 654938 218352 655174
rect 218588 654938 218620 655174
rect 218000 654854 218620 654938
rect 218000 654618 218032 654854
rect 218268 654618 218352 654854
rect 218588 654618 218620 654854
rect 254000 654938 254032 655174
rect 254268 654938 254352 655174
rect 254588 654938 254620 655174
rect 254000 654854 254620 654938
rect 254000 654618 254032 654854
rect 254268 654618 254352 654854
rect 254588 654618 254620 654854
rect 290000 654938 290032 655174
rect 290268 654938 290352 655174
rect 290588 654938 290620 655174
rect 290000 654854 290620 654938
rect 290000 654618 290032 654854
rect 290268 654618 290352 654854
rect 290588 654618 290620 654854
rect 326000 654938 326032 655174
rect 326268 654938 326352 655174
rect 326588 654938 326620 655174
rect 326000 654854 326620 654938
rect 326000 654618 326032 654854
rect 326268 654618 326352 654854
rect 326588 654618 326620 654854
rect 362000 654938 362032 655174
rect 362268 654938 362352 655174
rect 362588 654938 362620 655174
rect 362000 654854 362620 654938
rect 362000 654618 362032 654854
rect 362268 654618 362352 654854
rect 362588 654618 362620 654854
rect 398000 654938 398032 655174
rect 398268 654938 398352 655174
rect 398588 654938 398620 655174
rect 398000 654854 398620 654938
rect 398000 654618 398032 654854
rect 398268 654618 398352 654854
rect 398588 654618 398620 654854
rect 434000 654938 434032 655174
rect 434268 654938 434352 655174
rect 434588 654938 434620 655174
rect 434000 654854 434620 654938
rect 434000 654618 434032 654854
rect 434268 654618 434352 654854
rect 434588 654618 434620 654854
rect 470000 654938 470032 655174
rect 470268 654938 470352 655174
rect 470588 654938 470620 655174
rect 470000 654854 470620 654938
rect 470000 654618 470032 654854
rect 470268 654618 470352 654854
rect 470588 654618 470620 654854
rect 506000 654938 506032 655174
rect 506268 654938 506352 655174
rect 506588 654938 506620 655174
rect 506000 654854 506620 654938
rect 506000 654618 506032 654854
rect 506268 654618 506352 654854
rect 506588 654618 506620 654854
rect 542000 654938 542032 655174
rect 542268 654938 542352 655174
rect 542588 654938 542620 655174
rect 542000 654854 542620 654938
rect 542000 654618 542032 654854
rect 542268 654618 542352 654854
rect 542588 654618 542620 654854
rect 571500 654938 571532 655174
rect 571768 654938 571852 655174
rect 572088 654938 572120 655174
rect 571500 654854 572120 654938
rect 571500 654618 571532 654854
rect 571768 654618 571852 654854
rect 572088 654618 572120 654854
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect 9084 651218 9116 651454
rect 9352 651218 9436 651454
rect 9672 651218 9704 651454
rect 9084 651134 9704 651218
rect 9084 650898 9116 651134
rect 9352 650898 9436 651134
rect 9672 650898 9704 651134
rect 56620 651218 56652 651454
rect 56888 651218 56972 651454
rect 57208 651218 57240 651454
rect 56620 651134 57240 651218
rect 56620 650898 56652 651134
rect 56888 650898 56972 651134
rect 57208 650898 57240 651134
rect 92620 651218 92652 651454
rect 92888 651218 92972 651454
rect 93208 651218 93240 651454
rect 92620 651134 93240 651218
rect 92620 650898 92652 651134
rect 92888 650898 92972 651134
rect 93208 650898 93240 651134
rect 128620 651218 128652 651454
rect 128888 651218 128972 651454
rect 129208 651218 129240 651454
rect 128620 651134 129240 651218
rect 128620 650898 128652 651134
rect 128888 650898 128972 651134
rect 129208 650898 129240 651134
rect 164620 651218 164652 651454
rect 164888 651218 164972 651454
rect 165208 651218 165240 651454
rect 164620 651134 165240 651218
rect 164620 650898 164652 651134
rect 164888 650898 164972 651134
rect 165208 650898 165240 651134
rect 200620 651218 200652 651454
rect 200888 651218 200972 651454
rect 201208 651218 201240 651454
rect 200620 651134 201240 651218
rect 200620 650898 200652 651134
rect 200888 650898 200972 651134
rect 201208 650898 201240 651134
rect 236620 651218 236652 651454
rect 236888 651218 236972 651454
rect 237208 651218 237240 651454
rect 236620 651134 237240 651218
rect 236620 650898 236652 651134
rect 236888 650898 236972 651134
rect 237208 650898 237240 651134
rect 272620 651218 272652 651454
rect 272888 651218 272972 651454
rect 273208 651218 273240 651454
rect 272620 651134 273240 651218
rect 272620 650898 272652 651134
rect 272888 650898 272972 651134
rect 273208 650898 273240 651134
rect 308620 651218 308652 651454
rect 308888 651218 308972 651454
rect 309208 651218 309240 651454
rect 308620 651134 309240 651218
rect 308620 650898 308652 651134
rect 308888 650898 308972 651134
rect 309208 650898 309240 651134
rect 344620 651218 344652 651454
rect 344888 651218 344972 651454
rect 345208 651218 345240 651454
rect 344620 651134 345240 651218
rect 344620 650898 344652 651134
rect 344888 650898 344972 651134
rect 345208 650898 345240 651134
rect 380620 651218 380652 651454
rect 380888 651218 380972 651454
rect 381208 651218 381240 651454
rect 380620 651134 381240 651218
rect 380620 650898 380652 651134
rect 380888 650898 380972 651134
rect 381208 650898 381240 651134
rect 416620 651218 416652 651454
rect 416888 651218 416972 651454
rect 417208 651218 417240 651454
rect 416620 651134 417240 651218
rect 416620 650898 416652 651134
rect 416888 650898 416972 651134
rect 417208 650898 417240 651134
rect 452620 651218 452652 651454
rect 452888 651218 452972 651454
rect 453208 651218 453240 651454
rect 452620 651134 453240 651218
rect 452620 650898 452652 651134
rect 452888 650898 452972 651134
rect 453208 650898 453240 651134
rect 488620 651218 488652 651454
rect 488888 651218 488972 651454
rect 489208 651218 489240 651454
rect 488620 651134 489240 651218
rect 488620 650898 488652 651134
rect 488888 650898 488972 651134
rect 489208 650898 489240 651134
rect 524620 651218 524652 651454
rect 524888 651218 524972 651454
rect 525208 651218 525240 651454
rect 524620 651134 525240 651218
rect 524620 650898 524652 651134
rect 524888 650898 524972 651134
rect 525208 650898 525240 651134
rect 560620 651218 560652 651454
rect 560888 651218 560972 651454
rect 561208 651218 561240 651454
rect 560620 651134 561240 651218
rect 560620 650898 560652 651134
rect 560888 650898 560972 651134
rect 561208 650898 561240 651134
rect 570260 651218 570292 651454
rect 570528 651218 570612 651454
rect 570848 651218 570880 651454
rect 570260 651134 570880 651218
rect 570260 650898 570292 651134
rect 570528 650898 570612 651134
rect 570848 650898 570880 651134
rect -2006 615454 -1386 650898
rect 581514 619174 582134 654618
rect 7844 618938 7876 619174
rect 8112 618938 8196 619174
rect 8432 618938 8464 619174
rect 7844 618854 8464 618938
rect 7844 618618 7876 618854
rect 8112 618618 8196 618854
rect 8432 618618 8464 618854
rect 38000 618938 38032 619174
rect 38268 618938 38352 619174
rect 38588 618938 38620 619174
rect 38000 618854 38620 618938
rect 38000 618618 38032 618854
rect 38268 618618 38352 618854
rect 38588 618618 38620 618854
rect 74000 618938 74032 619174
rect 74268 618938 74352 619174
rect 74588 618938 74620 619174
rect 74000 618854 74620 618938
rect 74000 618618 74032 618854
rect 74268 618618 74352 618854
rect 74588 618618 74620 618854
rect 110000 618938 110032 619174
rect 110268 618938 110352 619174
rect 110588 618938 110620 619174
rect 110000 618854 110620 618938
rect 110000 618618 110032 618854
rect 110268 618618 110352 618854
rect 110588 618618 110620 618854
rect 146000 618938 146032 619174
rect 146268 618938 146352 619174
rect 146588 618938 146620 619174
rect 146000 618854 146620 618938
rect 146000 618618 146032 618854
rect 146268 618618 146352 618854
rect 146588 618618 146620 618854
rect 182000 618938 182032 619174
rect 182268 618938 182352 619174
rect 182588 618938 182620 619174
rect 182000 618854 182620 618938
rect 182000 618618 182032 618854
rect 182268 618618 182352 618854
rect 182588 618618 182620 618854
rect 218000 618938 218032 619174
rect 218268 618938 218352 619174
rect 218588 618938 218620 619174
rect 218000 618854 218620 618938
rect 218000 618618 218032 618854
rect 218268 618618 218352 618854
rect 218588 618618 218620 618854
rect 254000 618938 254032 619174
rect 254268 618938 254352 619174
rect 254588 618938 254620 619174
rect 254000 618854 254620 618938
rect 254000 618618 254032 618854
rect 254268 618618 254352 618854
rect 254588 618618 254620 618854
rect 290000 618938 290032 619174
rect 290268 618938 290352 619174
rect 290588 618938 290620 619174
rect 290000 618854 290620 618938
rect 290000 618618 290032 618854
rect 290268 618618 290352 618854
rect 290588 618618 290620 618854
rect 326000 618938 326032 619174
rect 326268 618938 326352 619174
rect 326588 618938 326620 619174
rect 326000 618854 326620 618938
rect 326000 618618 326032 618854
rect 326268 618618 326352 618854
rect 326588 618618 326620 618854
rect 362000 618938 362032 619174
rect 362268 618938 362352 619174
rect 362588 618938 362620 619174
rect 362000 618854 362620 618938
rect 362000 618618 362032 618854
rect 362268 618618 362352 618854
rect 362588 618618 362620 618854
rect 398000 618938 398032 619174
rect 398268 618938 398352 619174
rect 398588 618938 398620 619174
rect 398000 618854 398620 618938
rect 398000 618618 398032 618854
rect 398268 618618 398352 618854
rect 398588 618618 398620 618854
rect 434000 618938 434032 619174
rect 434268 618938 434352 619174
rect 434588 618938 434620 619174
rect 434000 618854 434620 618938
rect 434000 618618 434032 618854
rect 434268 618618 434352 618854
rect 434588 618618 434620 618854
rect 470000 618938 470032 619174
rect 470268 618938 470352 619174
rect 470588 618938 470620 619174
rect 470000 618854 470620 618938
rect 470000 618618 470032 618854
rect 470268 618618 470352 618854
rect 470588 618618 470620 618854
rect 506000 618938 506032 619174
rect 506268 618938 506352 619174
rect 506588 618938 506620 619174
rect 506000 618854 506620 618938
rect 506000 618618 506032 618854
rect 506268 618618 506352 618854
rect 506588 618618 506620 618854
rect 542000 618938 542032 619174
rect 542268 618938 542352 619174
rect 542588 618938 542620 619174
rect 542000 618854 542620 618938
rect 542000 618618 542032 618854
rect 542268 618618 542352 618854
rect 542588 618618 542620 618854
rect 571500 618938 571532 619174
rect 571768 618938 571852 619174
rect 572088 618938 572120 619174
rect 571500 618854 572120 618938
rect 571500 618618 571532 618854
rect 571768 618618 571852 618854
rect 572088 618618 572120 618854
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect 9084 615218 9116 615454
rect 9352 615218 9436 615454
rect 9672 615218 9704 615454
rect 9084 615134 9704 615218
rect 9084 614898 9116 615134
rect 9352 614898 9436 615134
rect 9672 614898 9704 615134
rect 56620 615218 56652 615454
rect 56888 615218 56972 615454
rect 57208 615218 57240 615454
rect 56620 615134 57240 615218
rect 56620 614898 56652 615134
rect 56888 614898 56972 615134
rect 57208 614898 57240 615134
rect 92620 615218 92652 615454
rect 92888 615218 92972 615454
rect 93208 615218 93240 615454
rect 92620 615134 93240 615218
rect 92620 614898 92652 615134
rect 92888 614898 92972 615134
rect 93208 614898 93240 615134
rect 128620 615218 128652 615454
rect 128888 615218 128972 615454
rect 129208 615218 129240 615454
rect 128620 615134 129240 615218
rect 128620 614898 128652 615134
rect 128888 614898 128972 615134
rect 129208 614898 129240 615134
rect 164620 615218 164652 615454
rect 164888 615218 164972 615454
rect 165208 615218 165240 615454
rect 164620 615134 165240 615218
rect 164620 614898 164652 615134
rect 164888 614898 164972 615134
rect 165208 614898 165240 615134
rect 200620 615218 200652 615454
rect 200888 615218 200972 615454
rect 201208 615218 201240 615454
rect 200620 615134 201240 615218
rect 200620 614898 200652 615134
rect 200888 614898 200972 615134
rect 201208 614898 201240 615134
rect 236620 615218 236652 615454
rect 236888 615218 236972 615454
rect 237208 615218 237240 615454
rect 236620 615134 237240 615218
rect 236620 614898 236652 615134
rect 236888 614898 236972 615134
rect 237208 614898 237240 615134
rect 272620 615218 272652 615454
rect 272888 615218 272972 615454
rect 273208 615218 273240 615454
rect 272620 615134 273240 615218
rect 272620 614898 272652 615134
rect 272888 614898 272972 615134
rect 273208 614898 273240 615134
rect 308620 615218 308652 615454
rect 308888 615218 308972 615454
rect 309208 615218 309240 615454
rect 308620 615134 309240 615218
rect 308620 614898 308652 615134
rect 308888 614898 308972 615134
rect 309208 614898 309240 615134
rect 344620 615218 344652 615454
rect 344888 615218 344972 615454
rect 345208 615218 345240 615454
rect 344620 615134 345240 615218
rect 344620 614898 344652 615134
rect 344888 614898 344972 615134
rect 345208 614898 345240 615134
rect 380620 615218 380652 615454
rect 380888 615218 380972 615454
rect 381208 615218 381240 615454
rect 380620 615134 381240 615218
rect 380620 614898 380652 615134
rect 380888 614898 380972 615134
rect 381208 614898 381240 615134
rect 416620 615218 416652 615454
rect 416888 615218 416972 615454
rect 417208 615218 417240 615454
rect 416620 615134 417240 615218
rect 416620 614898 416652 615134
rect 416888 614898 416972 615134
rect 417208 614898 417240 615134
rect 452620 615218 452652 615454
rect 452888 615218 452972 615454
rect 453208 615218 453240 615454
rect 452620 615134 453240 615218
rect 452620 614898 452652 615134
rect 452888 614898 452972 615134
rect 453208 614898 453240 615134
rect 488620 615218 488652 615454
rect 488888 615218 488972 615454
rect 489208 615218 489240 615454
rect 488620 615134 489240 615218
rect 488620 614898 488652 615134
rect 488888 614898 488972 615134
rect 489208 614898 489240 615134
rect 524620 615218 524652 615454
rect 524888 615218 524972 615454
rect 525208 615218 525240 615454
rect 524620 615134 525240 615218
rect 524620 614898 524652 615134
rect 524888 614898 524972 615134
rect 525208 614898 525240 615134
rect 560620 615218 560652 615454
rect 560888 615218 560972 615454
rect 561208 615218 561240 615454
rect 560620 615134 561240 615218
rect 560620 614898 560652 615134
rect 560888 614898 560972 615134
rect 561208 614898 561240 615134
rect 570260 615218 570292 615454
rect 570528 615218 570612 615454
rect 570848 615218 570880 615454
rect 570260 615134 570880 615218
rect 570260 614898 570292 615134
rect 570528 614898 570612 615134
rect 570848 614898 570880 615134
rect -2006 579454 -1386 614898
rect 581514 583174 582134 618618
rect 7844 582938 7876 583174
rect 8112 582938 8196 583174
rect 8432 582938 8464 583174
rect 7844 582854 8464 582938
rect 7844 582618 7876 582854
rect 8112 582618 8196 582854
rect 8432 582618 8464 582854
rect 38000 582938 38032 583174
rect 38268 582938 38352 583174
rect 38588 582938 38620 583174
rect 38000 582854 38620 582938
rect 38000 582618 38032 582854
rect 38268 582618 38352 582854
rect 38588 582618 38620 582854
rect 74000 582938 74032 583174
rect 74268 582938 74352 583174
rect 74588 582938 74620 583174
rect 74000 582854 74620 582938
rect 74000 582618 74032 582854
rect 74268 582618 74352 582854
rect 74588 582618 74620 582854
rect 110000 582938 110032 583174
rect 110268 582938 110352 583174
rect 110588 582938 110620 583174
rect 110000 582854 110620 582938
rect 110000 582618 110032 582854
rect 110268 582618 110352 582854
rect 110588 582618 110620 582854
rect 146000 582938 146032 583174
rect 146268 582938 146352 583174
rect 146588 582938 146620 583174
rect 146000 582854 146620 582938
rect 146000 582618 146032 582854
rect 146268 582618 146352 582854
rect 146588 582618 146620 582854
rect 182000 582938 182032 583174
rect 182268 582938 182352 583174
rect 182588 582938 182620 583174
rect 182000 582854 182620 582938
rect 182000 582618 182032 582854
rect 182268 582618 182352 582854
rect 182588 582618 182620 582854
rect 218000 582938 218032 583174
rect 218268 582938 218352 583174
rect 218588 582938 218620 583174
rect 218000 582854 218620 582938
rect 218000 582618 218032 582854
rect 218268 582618 218352 582854
rect 218588 582618 218620 582854
rect 254000 582938 254032 583174
rect 254268 582938 254352 583174
rect 254588 582938 254620 583174
rect 254000 582854 254620 582938
rect 254000 582618 254032 582854
rect 254268 582618 254352 582854
rect 254588 582618 254620 582854
rect 290000 582938 290032 583174
rect 290268 582938 290352 583174
rect 290588 582938 290620 583174
rect 290000 582854 290620 582938
rect 290000 582618 290032 582854
rect 290268 582618 290352 582854
rect 290588 582618 290620 582854
rect 326000 582938 326032 583174
rect 326268 582938 326352 583174
rect 326588 582938 326620 583174
rect 326000 582854 326620 582938
rect 326000 582618 326032 582854
rect 326268 582618 326352 582854
rect 326588 582618 326620 582854
rect 362000 582938 362032 583174
rect 362268 582938 362352 583174
rect 362588 582938 362620 583174
rect 362000 582854 362620 582938
rect 362000 582618 362032 582854
rect 362268 582618 362352 582854
rect 362588 582618 362620 582854
rect 398000 582938 398032 583174
rect 398268 582938 398352 583174
rect 398588 582938 398620 583174
rect 398000 582854 398620 582938
rect 398000 582618 398032 582854
rect 398268 582618 398352 582854
rect 398588 582618 398620 582854
rect 434000 582938 434032 583174
rect 434268 582938 434352 583174
rect 434588 582938 434620 583174
rect 434000 582854 434620 582938
rect 434000 582618 434032 582854
rect 434268 582618 434352 582854
rect 434588 582618 434620 582854
rect 470000 582938 470032 583174
rect 470268 582938 470352 583174
rect 470588 582938 470620 583174
rect 470000 582854 470620 582938
rect 470000 582618 470032 582854
rect 470268 582618 470352 582854
rect 470588 582618 470620 582854
rect 506000 582938 506032 583174
rect 506268 582938 506352 583174
rect 506588 582938 506620 583174
rect 506000 582854 506620 582938
rect 506000 582618 506032 582854
rect 506268 582618 506352 582854
rect 506588 582618 506620 582854
rect 542000 582938 542032 583174
rect 542268 582938 542352 583174
rect 542588 582938 542620 583174
rect 542000 582854 542620 582938
rect 542000 582618 542032 582854
rect 542268 582618 542352 582854
rect 542588 582618 542620 582854
rect 571500 582938 571532 583174
rect 571768 582938 571852 583174
rect 572088 582938 572120 583174
rect 571500 582854 572120 582938
rect 571500 582618 571532 582854
rect 571768 582618 571852 582854
rect 572088 582618 572120 582854
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect 9084 579218 9116 579454
rect 9352 579218 9436 579454
rect 9672 579218 9704 579454
rect 9084 579134 9704 579218
rect 9084 578898 9116 579134
rect 9352 578898 9436 579134
rect 9672 578898 9704 579134
rect 56620 579218 56652 579454
rect 56888 579218 56972 579454
rect 57208 579218 57240 579454
rect 56620 579134 57240 579218
rect 56620 578898 56652 579134
rect 56888 578898 56972 579134
rect 57208 578898 57240 579134
rect 92620 579218 92652 579454
rect 92888 579218 92972 579454
rect 93208 579218 93240 579454
rect 92620 579134 93240 579218
rect 92620 578898 92652 579134
rect 92888 578898 92972 579134
rect 93208 578898 93240 579134
rect 128620 579218 128652 579454
rect 128888 579218 128972 579454
rect 129208 579218 129240 579454
rect 128620 579134 129240 579218
rect 128620 578898 128652 579134
rect 128888 578898 128972 579134
rect 129208 578898 129240 579134
rect 164620 579218 164652 579454
rect 164888 579218 164972 579454
rect 165208 579218 165240 579454
rect 164620 579134 165240 579218
rect 164620 578898 164652 579134
rect 164888 578898 164972 579134
rect 165208 578898 165240 579134
rect 200620 579218 200652 579454
rect 200888 579218 200972 579454
rect 201208 579218 201240 579454
rect 200620 579134 201240 579218
rect 200620 578898 200652 579134
rect 200888 578898 200972 579134
rect 201208 578898 201240 579134
rect 236620 579218 236652 579454
rect 236888 579218 236972 579454
rect 237208 579218 237240 579454
rect 236620 579134 237240 579218
rect 236620 578898 236652 579134
rect 236888 578898 236972 579134
rect 237208 578898 237240 579134
rect 272620 579218 272652 579454
rect 272888 579218 272972 579454
rect 273208 579218 273240 579454
rect 272620 579134 273240 579218
rect 272620 578898 272652 579134
rect 272888 578898 272972 579134
rect 273208 578898 273240 579134
rect 308620 579218 308652 579454
rect 308888 579218 308972 579454
rect 309208 579218 309240 579454
rect 308620 579134 309240 579218
rect 308620 578898 308652 579134
rect 308888 578898 308972 579134
rect 309208 578898 309240 579134
rect 344620 579218 344652 579454
rect 344888 579218 344972 579454
rect 345208 579218 345240 579454
rect 344620 579134 345240 579218
rect 344620 578898 344652 579134
rect 344888 578898 344972 579134
rect 345208 578898 345240 579134
rect 380620 579218 380652 579454
rect 380888 579218 380972 579454
rect 381208 579218 381240 579454
rect 380620 579134 381240 579218
rect 380620 578898 380652 579134
rect 380888 578898 380972 579134
rect 381208 578898 381240 579134
rect 416620 579218 416652 579454
rect 416888 579218 416972 579454
rect 417208 579218 417240 579454
rect 416620 579134 417240 579218
rect 416620 578898 416652 579134
rect 416888 578898 416972 579134
rect 417208 578898 417240 579134
rect 452620 579218 452652 579454
rect 452888 579218 452972 579454
rect 453208 579218 453240 579454
rect 452620 579134 453240 579218
rect 452620 578898 452652 579134
rect 452888 578898 452972 579134
rect 453208 578898 453240 579134
rect 488620 579218 488652 579454
rect 488888 579218 488972 579454
rect 489208 579218 489240 579454
rect 488620 579134 489240 579218
rect 488620 578898 488652 579134
rect 488888 578898 488972 579134
rect 489208 578898 489240 579134
rect 524620 579218 524652 579454
rect 524888 579218 524972 579454
rect 525208 579218 525240 579454
rect 524620 579134 525240 579218
rect 524620 578898 524652 579134
rect 524888 578898 524972 579134
rect 525208 578898 525240 579134
rect 560620 579218 560652 579454
rect 560888 579218 560972 579454
rect 561208 579218 561240 579454
rect 560620 579134 561240 579218
rect 560620 578898 560652 579134
rect 560888 578898 560972 579134
rect 561208 578898 561240 579134
rect 570260 579218 570292 579454
rect 570528 579218 570612 579454
rect 570848 579218 570880 579454
rect 570260 579134 570880 579218
rect 570260 578898 570292 579134
rect 570528 578898 570612 579134
rect 570848 578898 570880 579134
rect -2006 543454 -1386 578898
rect 581514 547174 582134 582618
rect 7844 546938 7876 547174
rect 8112 546938 8196 547174
rect 8432 546938 8464 547174
rect 7844 546854 8464 546938
rect 7844 546618 7876 546854
rect 8112 546618 8196 546854
rect 8432 546618 8464 546854
rect 38000 546938 38032 547174
rect 38268 546938 38352 547174
rect 38588 546938 38620 547174
rect 38000 546854 38620 546938
rect 38000 546618 38032 546854
rect 38268 546618 38352 546854
rect 38588 546618 38620 546854
rect 74000 546938 74032 547174
rect 74268 546938 74352 547174
rect 74588 546938 74620 547174
rect 74000 546854 74620 546938
rect 74000 546618 74032 546854
rect 74268 546618 74352 546854
rect 74588 546618 74620 546854
rect 110000 546938 110032 547174
rect 110268 546938 110352 547174
rect 110588 546938 110620 547174
rect 110000 546854 110620 546938
rect 110000 546618 110032 546854
rect 110268 546618 110352 546854
rect 110588 546618 110620 546854
rect 146000 546938 146032 547174
rect 146268 546938 146352 547174
rect 146588 546938 146620 547174
rect 146000 546854 146620 546938
rect 146000 546618 146032 546854
rect 146268 546618 146352 546854
rect 146588 546618 146620 546854
rect 182000 546938 182032 547174
rect 182268 546938 182352 547174
rect 182588 546938 182620 547174
rect 182000 546854 182620 546938
rect 182000 546618 182032 546854
rect 182268 546618 182352 546854
rect 182588 546618 182620 546854
rect 218000 546938 218032 547174
rect 218268 546938 218352 547174
rect 218588 546938 218620 547174
rect 218000 546854 218620 546938
rect 218000 546618 218032 546854
rect 218268 546618 218352 546854
rect 218588 546618 218620 546854
rect 254000 546938 254032 547174
rect 254268 546938 254352 547174
rect 254588 546938 254620 547174
rect 254000 546854 254620 546938
rect 254000 546618 254032 546854
rect 254268 546618 254352 546854
rect 254588 546618 254620 546854
rect 290000 546938 290032 547174
rect 290268 546938 290352 547174
rect 290588 546938 290620 547174
rect 290000 546854 290620 546938
rect 290000 546618 290032 546854
rect 290268 546618 290352 546854
rect 290588 546618 290620 546854
rect 326000 546938 326032 547174
rect 326268 546938 326352 547174
rect 326588 546938 326620 547174
rect 326000 546854 326620 546938
rect 326000 546618 326032 546854
rect 326268 546618 326352 546854
rect 326588 546618 326620 546854
rect 362000 546938 362032 547174
rect 362268 546938 362352 547174
rect 362588 546938 362620 547174
rect 362000 546854 362620 546938
rect 362000 546618 362032 546854
rect 362268 546618 362352 546854
rect 362588 546618 362620 546854
rect 398000 546938 398032 547174
rect 398268 546938 398352 547174
rect 398588 546938 398620 547174
rect 398000 546854 398620 546938
rect 398000 546618 398032 546854
rect 398268 546618 398352 546854
rect 398588 546618 398620 546854
rect 434000 546938 434032 547174
rect 434268 546938 434352 547174
rect 434588 546938 434620 547174
rect 434000 546854 434620 546938
rect 434000 546618 434032 546854
rect 434268 546618 434352 546854
rect 434588 546618 434620 546854
rect 470000 546938 470032 547174
rect 470268 546938 470352 547174
rect 470588 546938 470620 547174
rect 470000 546854 470620 546938
rect 470000 546618 470032 546854
rect 470268 546618 470352 546854
rect 470588 546618 470620 546854
rect 506000 546938 506032 547174
rect 506268 546938 506352 547174
rect 506588 546938 506620 547174
rect 506000 546854 506620 546938
rect 506000 546618 506032 546854
rect 506268 546618 506352 546854
rect 506588 546618 506620 546854
rect 542000 546938 542032 547174
rect 542268 546938 542352 547174
rect 542588 546938 542620 547174
rect 542000 546854 542620 546938
rect 542000 546618 542032 546854
rect 542268 546618 542352 546854
rect 542588 546618 542620 546854
rect 571500 546938 571532 547174
rect 571768 546938 571852 547174
rect 572088 546938 572120 547174
rect 571500 546854 572120 546938
rect 571500 546618 571532 546854
rect 571768 546618 571852 546854
rect 572088 546618 572120 546854
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect 9084 543218 9116 543454
rect 9352 543218 9436 543454
rect 9672 543218 9704 543454
rect 9084 543134 9704 543218
rect 9084 542898 9116 543134
rect 9352 542898 9436 543134
rect 9672 542898 9704 543134
rect 56620 543218 56652 543454
rect 56888 543218 56972 543454
rect 57208 543218 57240 543454
rect 56620 543134 57240 543218
rect 56620 542898 56652 543134
rect 56888 542898 56972 543134
rect 57208 542898 57240 543134
rect 92620 543218 92652 543454
rect 92888 543218 92972 543454
rect 93208 543218 93240 543454
rect 92620 543134 93240 543218
rect 92620 542898 92652 543134
rect 92888 542898 92972 543134
rect 93208 542898 93240 543134
rect 128620 543218 128652 543454
rect 128888 543218 128972 543454
rect 129208 543218 129240 543454
rect 128620 543134 129240 543218
rect 128620 542898 128652 543134
rect 128888 542898 128972 543134
rect 129208 542898 129240 543134
rect 164620 543218 164652 543454
rect 164888 543218 164972 543454
rect 165208 543218 165240 543454
rect 164620 543134 165240 543218
rect 164620 542898 164652 543134
rect 164888 542898 164972 543134
rect 165208 542898 165240 543134
rect 200620 543218 200652 543454
rect 200888 543218 200972 543454
rect 201208 543218 201240 543454
rect 200620 543134 201240 543218
rect 200620 542898 200652 543134
rect 200888 542898 200972 543134
rect 201208 542898 201240 543134
rect 236620 543218 236652 543454
rect 236888 543218 236972 543454
rect 237208 543218 237240 543454
rect 236620 543134 237240 543218
rect 236620 542898 236652 543134
rect 236888 542898 236972 543134
rect 237208 542898 237240 543134
rect 272620 543218 272652 543454
rect 272888 543218 272972 543454
rect 273208 543218 273240 543454
rect 272620 543134 273240 543218
rect 272620 542898 272652 543134
rect 272888 542898 272972 543134
rect 273208 542898 273240 543134
rect 308620 543218 308652 543454
rect 308888 543218 308972 543454
rect 309208 543218 309240 543454
rect 308620 543134 309240 543218
rect 308620 542898 308652 543134
rect 308888 542898 308972 543134
rect 309208 542898 309240 543134
rect 344620 543218 344652 543454
rect 344888 543218 344972 543454
rect 345208 543218 345240 543454
rect 344620 543134 345240 543218
rect 344620 542898 344652 543134
rect 344888 542898 344972 543134
rect 345208 542898 345240 543134
rect 380620 543218 380652 543454
rect 380888 543218 380972 543454
rect 381208 543218 381240 543454
rect 380620 543134 381240 543218
rect 380620 542898 380652 543134
rect 380888 542898 380972 543134
rect 381208 542898 381240 543134
rect 416620 543218 416652 543454
rect 416888 543218 416972 543454
rect 417208 543218 417240 543454
rect 416620 543134 417240 543218
rect 416620 542898 416652 543134
rect 416888 542898 416972 543134
rect 417208 542898 417240 543134
rect 452620 543218 452652 543454
rect 452888 543218 452972 543454
rect 453208 543218 453240 543454
rect 452620 543134 453240 543218
rect 452620 542898 452652 543134
rect 452888 542898 452972 543134
rect 453208 542898 453240 543134
rect 488620 543218 488652 543454
rect 488888 543218 488972 543454
rect 489208 543218 489240 543454
rect 488620 543134 489240 543218
rect 488620 542898 488652 543134
rect 488888 542898 488972 543134
rect 489208 542898 489240 543134
rect 524620 543218 524652 543454
rect 524888 543218 524972 543454
rect 525208 543218 525240 543454
rect 524620 543134 525240 543218
rect 524620 542898 524652 543134
rect 524888 542898 524972 543134
rect 525208 542898 525240 543134
rect 560620 543218 560652 543454
rect 560888 543218 560972 543454
rect 561208 543218 561240 543454
rect 560620 543134 561240 543218
rect 560620 542898 560652 543134
rect 560888 542898 560972 543134
rect 561208 542898 561240 543134
rect 570260 543218 570292 543454
rect 570528 543218 570612 543454
rect 570848 543218 570880 543454
rect 570260 543134 570880 543218
rect 570260 542898 570292 543134
rect 570528 542898 570612 543134
rect 570848 542898 570880 543134
rect -2006 507454 -1386 542898
rect 60560 511174 60920 511206
rect 7844 510938 7876 511174
rect 8112 510938 8196 511174
rect 8432 510938 8464 511174
rect 7844 510854 8464 510938
rect 7844 510618 7876 510854
rect 8112 510618 8196 510854
rect 8432 510618 8464 510854
rect 38000 510938 38032 511174
rect 38268 510938 38352 511174
rect 38588 510938 38620 511174
rect 38000 510854 38620 510938
rect 38000 510618 38032 510854
rect 38268 510618 38352 510854
rect 38588 510618 38620 510854
rect 60560 510938 60622 511174
rect 60858 510938 60920 511174
rect 60560 510854 60920 510938
rect 60560 510618 60622 510854
rect 60858 510618 60920 510854
rect 60560 510586 60920 510618
rect 159036 511174 159396 511206
rect 185560 511174 185920 511206
rect 159036 510938 159098 511174
rect 159334 510938 159396 511174
rect 159036 510854 159396 510938
rect 159036 510618 159098 510854
rect 159334 510618 159396 510854
rect 182000 510938 182032 511174
rect 182268 510938 182352 511174
rect 182588 510938 182620 511174
rect 182000 510854 182620 510938
rect 182000 510618 182032 510854
rect 182268 510618 182352 510854
rect 182588 510618 182620 510854
rect 185560 510938 185622 511174
rect 185858 510938 185920 511174
rect 185560 510854 185920 510938
rect 185560 510618 185622 510854
rect 185858 510618 185920 510854
rect 159036 510586 159396 510618
rect 185560 510586 185920 510618
rect 284036 511174 284396 511206
rect 310560 511174 310920 511206
rect 284036 510938 284098 511174
rect 284334 510938 284396 511174
rect 284036 510854 284396 510938
rect 284036 510618 284098 510854
rect 284334 510618 284396 510854
rect 290000 510938 290032 511174
rect 290268 510938 290352 511174
rect 290588 510938 290620 511174
rect 290000 510854 290620 510938
rect 290000 510618 290032 510854
rect 290268 510618 290352 510854
rect 290588 510618 290620 510854
rect 310560 510938 310622 511174
rect 310858 510938 310920 511174
rect 310560 510854 310920 510938
rect 310560 510618 310622 510854
rect 310858 510618 310920 510854
rect 284036 510586 284396 510618
rect 310560 510586 310920 510618
rect 409036 511174 409396 511206
rect 436560 511174 436920 511206
rect 409036 510938 409098 511174
rect 409334 510938 409396 511174
rect 409036 510854 409396 510938
rect 409036 510618 409098 510854
rect 409334 510618 409396 510854
rect 434000 510938 434032 511174
rect 434268 510938 434352 511174
rect 434588 510938 434620 511174
rect 434000 510854 434620 510938
rect 434000 510618 434032 510854
rect 434268 510618 434352 510854
rect 434588 510618 434620 510854
rect 436560 510938 436622 511174
rect 436858 510938 436920 511174
rect 436560 510854 436920 510938
rect 436560 510618 436622 510854
rect 436858 510618 436920 510854
rect 409036 510586 409396 510618
rect 436560 510586 436920 510618
rect 535036 511174 535396 511206
rect 581514 511174 582134 546618
rect 535036 510938 535098 511174
rect 535334 510938 535396 511174
rect 535036 510854 535396 510938
rect 535036 510618 535098 510854
rect 535334 510618 535396 510854
rect 542000 510938 542032 511174
rect 542268 510938 542352 511174
rect 542588 510938 542620 511174
rect 542000 510854 542620 510938
rect 542000 510618 542032 510854
rect 542268 510618 542352 510854
rect 542588 510618 542620 510854
rect 571500 510938 571532 511174
rect 571768 510938 571852 511174
rect 572088 510938 572120 511174
rect 571500 510854 572120 510938
rect 571500 510618 571532 510854
rect 571768 510618 571852 510854
rect 572088 510618 572120 510854
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 535036 510586 535396 510618
rect 61280 507454 61640 507486
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect 9084 507218 9116 507454
rect 9352 507218 9436 507454
rect 9672 507218 9704 507454
rect 9084 507134 9704 507218
rect 9084 506898 9116 507134
rect 9352 506898 9436 507134
rect 9672 506898 9704 507134
rect 56620 507218 56652 507454
rect 56888 507218 56972 507454
rect 57208 507218 57240 507454
rect 56620 507134 57240 507218
rect 56620 506898 56652 507134
rect 56888 506898 56972 507134
rect 57208 506898 57240 507134
rect 61280 507218 61342 507454
rect 61578 507218 61640 507454
rect 61280 507134 61640 507218
rect 61280 506898 61342 507134
rect 61578 506898 61640 507134
rect -2006 471454 -1386 506898
rect 61280 506866 61640 506898
rect 158316 507454 158676 507486
rect 186280 507454 186640 507486
rect 158316 507218 158378 507454
rect 158614 507218 158676 507454
rect 158316 507134 158676 507218
rect 158316 506898 158378 507134
rect 158614 506898 158676 507134
rect 164620 507218 164652 507454
rect 164888 507218 164972 507454
rect 165208 507218 165240 507454
rect 164620 507134 165240 507218
rect 164620 506898 164652 507134
rect 164888 506898 164972 507134
rect 165208 506898 165240 507134
rect 186280 507218 186342 507454
rect 186578 507218 186640 507454
rect 186280 507134 186640 507218
rect 186280 506898 186342 507134
rect 186578 506898 186640 507134
rect 158316 506866 158676 506898
rect 186280 506866 186640 506898
rect 283316 507454 283676 507486
rect 311280 507454 311640 507486
rect 283316 507218 283378 507454
rect 283614 507218 283676 507454
rect 283316 507134 283676 507218
rect 283316 506898 283378 507134
rect 283614 506898 283676 507134
rect 308620 507218 308652 507454
rect 308888 507218 308972 507454
rect 309208 507218 309240 507454
rect 308620 507134 309240 507218
rect 308620 506898 308652 507134
rect 308888 506898 308972 507134
rect 309208 506898 309240 507134
rect 311280 507218 311342 507454
rect 311578 507218 311640 507454
rect 311280 507134 311640 507218
rect 311280 506898 311342 507134
rect 311578 506898 311640 507134
rect 283316 506866 283676 506898
rect 311280 506866 311640 506898
rect 408316 507454 408676 507486
rect 437280 507454 437640 507486
rect 408316 507218 408378 507454
rect 408614 507218 408676 507454
rect 408316 507134 408676 507218
rect 408316 506898 408378 507134
rect 408614 506898 408676 507134
rect 416620 507218 416652 507454
rect 416888 507218 416972 507454
rect 417208 507218 417240 507454
rect 416620 507134 417240 507218
rect 416620 506898 416652 507134
rect 416888 506898 416972 507134
rect 417208 506898 417240 507134
rect 437280 507218 437342 507454
rect 437578 507218 437640 507454
rect 437280 507134 437640 507218
rect 437280 506898 437342 507134
rect 437578 506898 437640 507134
rect 408316 506866 408676 506898
rect 437280 506866 437640 506898
rect 534316 507454 534676 507486
rect 534316 507218 534378 507454
rect 534614 507218 534676 507454
rect 534316 507134 534676 507218
rect 534316 506898 534378 507134
rect 534614 506898 534676 507134
rect 560620 507218 560652 507454
rect 560888 507218 560972 507454
rect 561208 507218 561240 507454
rect 560620 507134 561240 507218
rect 560620 506898 560652 507134
rect 560888 506898 560972 507134
rect 561208 506898 561240 507134
rect 570260 507218 570292 507454
rect 570528 507218 570612 507454
rect 570848 507218 570880 507454
rect 570260 507134 570880 507218
rect 570260 506898 570292 507134
rect 570528 506898 570612 507134
rect 570848 506898 570880 507134
rect 534316 506866 534676 506898
rect 60560 475174 60920 475206
rect 7844 474938 7876 475174
rect 8112 474938 8196 475174
rect 8432 474938 8464 475174
rect 7844 474854 8464 474938
rect 7844 474618 7876 474854
rect 8112 474618 8196 474854
rect 8432 474618 8464 474854
rect 38000 474938 38032 475174
rect 38268 474938 38352 475174
rect 38588 474938 38620 475174
rect 38000 474854 38620 474938
rect 38000 474618 38032 474854
rect 38268 474618 38352 474854
rect 38588 474618 38620 474854
rect 60560 474938 60622 475174
rect 60858 474938 60920 475174
rect 60560 474854 60920 474938
rect 60560 474618 60622 474854
rect 60858 474618 60920 474854
rect 60560 474586 60920 474618
rect 159036 475174 159396 475206
rect 185560 475174 185920 475206
rect 159036 474938 159098 475174
rect 159334 474938 159396 475174
rect 159036 474854 159396 474938
rect 159036 474618 159098 474854
rect 159334 474618 159396 474854
rect 182000 474938 182032 475174
rect 182268 474938 182352 475174
rect 182588 474938 182620 475174
rect 182000 474854 182620 474938
rect 182000 474618 182032 474854
rect 182268 474618 182352 474854
rect 182588 474618 182620 474854
rect 185560 474938 185622 475174
rect 185858 474938 185920 475174
rect 185560 474854 185920 474938
rect 185560 474618 185622 474854
rect 185858 474618 185920 474854
rect 159036 474586 159396 474618
rect 185560 474586 185920 474618
rect 284036 475174 284396 475206
rect 310560 475174 310920 475206
rect 284036 474938 284098 475174
rect 284334 474938 284396 475174
rect 284036 474854 284396 474938
rect 284036 474618 284098 474854
rect 284334 474618 284396 474854
rect 290000 474938 290032 475174
rect 290268 474938 290352 475174
rect 290588 474938 290620 475174
rect 290000 474854 290620 474938
rect 290000 474618 290032 474854
rect 290268 474618 290352 474854
rect 290588 474618 290620 474854
rect 310560 474938 310622 475174
rect 310858 474938 310920 475174
rect 310560 474854 310920 474938
rect 310560 474618 310622 474854
rect 310858 474618 310920 474854
rect 284036 474586 284396 474618
rect 310560 474586 310920 474618
rect 409036 475174 409396 475206
rect 436560 475174 436920 475206
rect 409036 474938 409098 475174
rect 409334 474938 409396 475174
rect 409036 474854 409396 474938
rect 409036 474618 409098 474854
rect 409334 474618 409396 474854
rect 434000 474938 434032 475174
rect 434268 474938 434352 475174
rect 434588 474938 434620 475174
rect 434000 474854 434620 474938
rect 434000 474618 434032 474854
rect 434268 474618 434352 474854
rect 434588 474618 434620 474854
rect 436560 474938 436622 475174
rect 436858 474938 436920 475174
rect 436560 474854 436920 474938
rect 436560 474618 436622 474854
rect 436858 474618 436920 474854
rect 409036 474586 409396 474618
rect 436560 474586 436920 474618
rect 535036 475174 535396 475206
rect 581514 475174 582134 510618
rect 535036 474938 535098 475174
rect 535334 474938 535396 475174
rect 535036 474854 535396 474938
rect 535036 474618 535098 474854
rect 535334 474618 535396 474854
rect 542000 474938 542032 475174
rect 542268 474938 542352 475174
rect 542588 474938 542620 475174
rect 542000 474854 542620 474938
rect 542000 474618 542032 474854
rect 542268 474618 542352 474854
rect 542588 474618 542620 474854
rect 571500 474938 571532 475174
rect 571768 474938 571852 475174
rect 572088 474938 572120 475174
rect 571500 474854 572120 474938
rect 571500 474618 571532 474854
rect 571768 474618 571852 474854
rect 572088 474618 572120 474854
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 535036 474586 535396 474618
rect 61280 471454 61640 471486
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect 9084 471218 9116 471454
rect 9352 471218 9436 471454
rect 9672 471218 9704 471454
rect 9084 471134 9704 471218
rect 9084 470898 9116 471134
rect 9352 470898 9436 471134
rect 9672 470898 9704 471134
rect 56620 471218 56652 471454
rect 56888 471218 56972 471454
rect 57208 471218 57240 471454
rect 56620 471134 57240 471218
rect 56620 470898 56652 471134
rect 56888 470898 56972 471134
rect 57208 470898 57240 471134
rect 61280 471218 61342 471454
rect 61578 471218 61640 471454
rect 61280 471134 61640 471218
rect 61280 470898 61342 471134
rect 61578 470898 61640 471134
rect -2006 435454 -1386 470898
rect 61280 470866 61640 470898
rect 158316 471454 158676 471486
rect 186280 471454 186640 471486
rect 158316 471218 158378 471454
rect 158614 471218 158676 471454
rect 158316 471134 158676 471218
rect 158316 470898 158378 471134
rect 158614 470898 158676 471134
rect 164620 471218 164652 471454
rect 164888 471218 164972 471454
rect 165208 471218 165240 471454
rect 164620 471134 165240 471218
rect 164620 470898 164652 471134
rect 164888 470898 164972 471134
rect 165208 470898 165240 471134
rect 186280 471218 186342 471454
rect 186578 471218 186640 471454
rect 186280 471134 186640 471218
rect 186280 470898 186342 471134
rect 186578 470898 186640 471134
rect 158316 470866 158676 470898
rect 186280 470866 186640 470898
rect 283316 471454 283676 471486
rect 311280 471454 311640 471486
rect 283316 471218 283378 471454
rect 283614 471218 283676 471454
rect 283316 471134 283676 471218
rect 283316 470898 283378 471134
rect 283614 470898 283676 471134
rect 308620 471218 308652 471454
rect 308888 471218 308972 471454
rect 309208 471218 309240 471454
rect 308620 471134 309240 471218
rect 308620 470898 308652 471134
rect 308888 470898 308972 471134
rect 309208 470898 309240 471134
rect 311280 471218 311342 471454
rect 311578 471218 311640 471454
rect 311280 471134 311640 471218
rect 311280 470898 311342 471134
rect 311578 470898 311640 471134
rect 283316 470866 283676 470898
rect 311280 470866 311640 470898
rect 408316 471454 408676 471486
rect 437280 471454 437640 471486
rect 408316 471218 408378 471454
rect 408614 471218 408676 471454
rect 408316 471134 408676 471218
rect 408316 470898 408378 471134
rect 408614 470898 408676 471134
rect 416620 471218 416652 471454
rect 416888 471218 416972 471454
rect 417208 471218 417240 471454
rect 416620 471134 417240 471218
rect 416620 470898 416652 471134
rect 416888 470898 416972 471134
rect 417208 470898 417240 471134
rect 437280 471218 437342 471454
rect 437578 471218 437640 471454
rect 437280 471134 437640 471218
rect 437280 470898 437342 471134
rect 437578 470898 437640 471134
rect 408316 470866 408676 470898
rect 437280 470866 437640 470898
rect 534316 471454 534676 471486
rect 534316 471218 534378 471454
rect 534614 471218 534676 471454
rect 534316 471134 534676 471218
rect 534316 470898 534378 471134
rect 534614 470898 534676 471134
rect 560620 471218 560652 471454
rect 560888 471218 560972 471454
rect 561208 471218 561240 471454
rect 560620 471134 561240 471218
rect 560620 470898 560652 471134
rect 560888 470898 560972 471134
rect 561208 470898 561240 471134
rect 570260 471218 570292 471454
rect 570528 471218 570612 471454
rect 570848 471218 570880 471454
rect 570260 471134 570880 471218
rect 570260 470898 570292 471134
rect 570528 470898 570612 471134
rect 570848 470898 570880 471134
rect 534316 470866 534676 470898
rect 60560 439174 60920 439206
rect 7844 438938 7876 439174
rect 8112 438938 8196 439174
rect 8432 438938 8464 439174
rect 7844 438854 8464 438938
rect 7844 438618 7876 438854
rect 8112 438618 8196 438854
rect 8432 438618 8464 438854
rect 38000 438938 38032 439174
rect 38268 438938 38352 439174
rect 38588 438938 38620 439174
rect 38000 438854 38620 438938
rect 38000 438618 38032 438854
rect 38268 438618 38352 438854
rect 38588 438618 38620 438854
rect 60560 438938 60622 439174
rect 60858 438938 60920 439174
rect 60560 438854 60920 438938
rect 60560 438618 60622 438854
rect 60858 438618 60920 438854
rect 60560 438586 60920 438618
rect 159036 439174 159396 439206
rect 185560 439174 185920 439206
rect 159036 438938 159098 439174
rect 159334 438938 159396 439174
rect 159036 438854 159396 438938
rect 159036 438618 159098 438854
rect 159334 438618 159396 438854
rect 182000 438938 182032 439174
rect 182268 438938 182352 439174
rect 182588 438938 182620 439174
rect 182000 438854 182620 438938
rect 182000 438618 182032 438854
rect 182268 438618 182352 438854
rect 182588 438618 182620 438854
rect 185560 438938 185622 439174
rect 185858 438938 185920 439174
rect 185560 438854 185920 438938
rect 185560 438618 185622 438854
rect 185858 438618 185920 438854
rect 159036 438586 159396 438618
rect 185560 438586 185920 438618
rect 284036 439174 284396 439206
rect 310560 439174 310920 439206
rect 284036 438938 284098 439174
rect 284334 438938 284396 439174
rect 284036 438854 284396 438938
rect 284036 438618 284098 438854
rect 284334 438618 284396 438854
rect 290000 438938 290032 439174
rect 290268 438938 290352 439174
rect 290588 438938 290620 439174
rect 290000 438854 290620 438938
rect 290000 438618 290032 438854
rect 290268 438618 290352 438854
rect 290588 438618 290620 438854
rect 310560 438938 310622 439174
rect 310858 438938 310920 439174
rect 310560 438854 310920 438938
rect 310560 438618 310622 438854
rect 310858 438618 310920 438854
rect 284036 438586 284396 438618
rect 310560 438586 310920 438618
rect 409036 439174 409396 439206
rect 436560 439174 436920 439206
rect 409036 438938 409098 439174
rect 409334 438938 409396 439174
rect 409036 438854 409396 438938
rect 409036 438618 409098 438854
rect 409334 438618 409396 438854
rect 434000 438938 434032 439174
rect 434268 438938 434352 439174
rect 434588 438938 434620 439174
rect 434000 438854 434620 438938
rect 434000 438618 434032 438854
rect 434268 438618 434352 438854
rect 434588 438618 434620 438854
rect 436560 438938 436622 439174
rect 436858 438938 436920 439174
rect 436560 438854 436920 438938
rect 436560 438618 436622 438854
rect 436858 438618 436920 438854
rect 409036 438586 409396 438618
rect 436560 438586 436920 438618
rect 535036 439174 535396 439206
rect 581514 439174 582134 474618
rect 535036 438938 535098 439174
rect 535334 438938 535396 439174
rect 535036 438854 535396 438938
rect 535036 438618 535098 438854
rect 535334 438618 535396 438854
rect 542000 438938 542032 439174
rect 542268 438938 542352 439174
rect 542588 438938 542620 439174
rect 542000 438854 542620 438938
rect 542000 438618 542032 438854
rect 542268 438618 542352 438854
rect 542588 438618 542620 438854
rect 571500 438938 571532 439174
rect 571768 438938 571852 439174
rect 572088 438938 572120 439174
rect 571500 438854 572120 438938
rect 571500 438618 571532 438854
rect 571768 438618 571852 438854
rect 572088 438618 572120 438854
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 535036 438586 535396 438618
rect 61280 435454 61640 435486
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect 9084 435218 9116 435454
rect 9352 435218 9436 435454
rect 9672 435218 9704 435454
rect 9084 435134 9704 435218
rect 9084 434898 9116 435134
rect 9352 434898 9436 435134
rect 9672 434898 9704 435134
rect 56620 435218 56652 435454
rect 56888 435218 56972 435454
rect 57208 435218 57240 435454
rect 56620 435134 57240 435218
rect 56620 434898 56652 435134
rect 56888 434898 56972 435134
rect 57208 434898 57240 435134
rect 61280 435218 61342 435454
rect 61578 435218 61640 435454
rect 61280 435134 61640 435218
rect 61280 434898 61342 435134
rect 61578 434898 61640 435134
rect -2006 399454 -1386 434898
rect 61280 434866 61640 434898
rect 158316 435454 158676 435486
rect 186280 435454 186640 435486
rect 158316 435218 158378 435454
rect 158614 435218 158676 435454
rect 158316 435134 158676 435218
rect 158316 434898 158378 435134
rect 158614 434898 158676 435134
rect 164620 435218 164652 435454
rect 164888 435218 164972 435454
rect 165208 435218 165240 435454
rect 164620 435134 165240 435218
rect 164620 434898 164652 435134
rect 164888 434898 164972 435134
rect 165208 434898 165240 435134
rect 186280 435218 186342 435454
rect 186578 435218 186640 435454
rect 186280 435134 186640 435218
rect 186280 434898 186342 435134
rect 186578 434898 186640 435134
rect 158316 434866 158676 434898
rect 186280 434866 186640 434898
rect 283316 435454 283676 435486
rect 311280 435454 311640 435486
rect 283316 435218 283378 435454
rect 283614 435218 283676 435454
rect 283316 435134 283676 435218
rect 283316 434898 283378 435134
rect 283614 434898 283676 435134
rect 308620 435218 308652 435454
rect 308888 435218 308972 435454
rect 309208 435218 309240 435454
rect 308620 435134 309240 435218
rect 308620 434898 308652 435134
rect 308888 434898 308972 435134
rect 309208 434898 309240 435134
rect 311280 435218 311342 435454
rect 311578 435218 311640 435454
rect 311280 435134 311640 435218
rect 311280 434898 311342 435134
rect 311578 434898 311640 435134
rect 283316 434866 283676 434898
rect 311280 434866 311640 434898
rect 408316 435454 408676 435486
rect 437280 435454 437640 435486
rect 408316 435218 408378 435454
rect 408614 435218 408676 435454
rect 408316 435134 408676 435218
rect 408316 434898 408378 435134
rect 408614 434898 408676 435134
rect 416620 435218 416652 435454
rect 416888 435218 416972 435454
rect 417208 435218 417240 435454
rect 416620 435134 417240 435218
rect 416620 434898 416652 435134
rect 416888 434898 416972 435134
rect 417208 434898 417240 435134
rect 437280 435218 437342 435454
rect 437578 435218 437640 435454
rect 437280 435134 437640 435218
rect 437280 434898 437342 435134
rect 437578 434898 437640 435134
rect 408316 434866 408676 434898
rect 437280 434866 437640 434898
rect 534316 435454 534676 435486
rect 534316 435218 534378 435454
rect 534614 435218 534676 435454
rect 534316 435134 534676 435218
rect 534316 434898 534378 435134
rect 534614 434898 534676 435134
rect 560620 435218 560652 435454
rect 560888 435218 560972 435454
rect 561208 435218 561240 435454
rect 560620 435134 561240 435218
rect 560620 434898 560652 435134
rect 560888 434898 560972 435134
rect 561208 434898 561240 435134
rect 570260 435218 570292 435454
rect 570528 435218 570612 435454
rect 570848 435218 570880 435454
rect 570260 435134 570880 435218
rect 570260 434898 570292 435134
rect 570528 434898 570612 435134
rect 570848 434898 570880 435134
rect 534316 434866 534676 434898
rect 61280 433244 61640 433300
rect 61280 433008 61342 433244
rect 61578 433008 61640 433244
rect 61280 432952 61640 433008
rect 62952 433244 63300 433300
rect 62952 433008 63008 433244
rect 63244 433008 63300 433244
rect 62952 432952 63300 433008
rect 281656 433244 282004 433300
rect 281656 433008 281712 433244
rect 281948 433008 282004 433244
rect 281656 432952 282004 433008
rect 283316 433244 283676 433300
rect 283316 433008 283378 433244
rect 283614 433008 283676 433244
rect 283316 432952 283676 433008
rect 311280 433244 311640 433300
rect 311280 433008 311342 433244
rect 311578 433008 311640 433244
rect 311280 432952 311640 433008
rect 312952 433244 313300 433300
rect 312952 433008 313008 433244
rect 313244 433008 313300 433244
rect 312952 432952 313300 433008
rect 532656 433244 533004 433300
rect 532656 433008 532712 433244
rect 532948 433008 533004 433244
rect 532656 432952 533004 433008
rect 534316 433244 534676 433300
rect 534316 433008 534378 433244
rect 534614 433008 534676 433244
rect 534316 432952 534676 433008
rect 157336 432564 157684 432620
rect 157336 432328 157392 432564
rect 157628 432328 157684 432564
rect 157336 432272 157684 432328
rect 159036 432564 159396 432620
rect 159036 432328 159098 432564
rect 159334 432328 159396 432564
rect 159036 432272 159396 432328
rect 185560 432564 185920 432620
rect 185560 432328 185622 432564
rect 185858 432328 185920 432564
rect 185560 432272 185920 432328
rect 187272 432564 187620 432620
rect 187272 432328 187328 432564
rect 187564 432328 187620 432564
rect 187272 432272 187620 432328
rect 407336 432564 407684 432620
rect 407336 432328 407392 432564
rect 407628 432328 407684 432564
rect 407336 432272 407684 432328
rect 409036 432564 409396 432620
rect 409036 432328 409098 432564
rect 409334 432328 409396 432564
rect 409036 432272 409396 432328
rect 436560 432564 436920 432620
rect 436560 432328 436622 432564
rect 436858 432328 436920 432564
rect 436560 432272 436920 432328
rect 438272 432564 438620 432620
rect 438272 432328 438328 432564
rect 438564 432328 438620 432564
rect 438272 432272 438620 432328
rect 581514 403174 582134 438618
rect 7844 402938 7876 403174
rect 8112 402938 8196 403174
rect 8432 402938 8464 403174
rect 7844 402854 8464 402938
rect 7844 402618 7876 402854
rect 8112 402618 8196 402854
rect 8432 402618 8464 402854
rect 38000 402938 38032 403174
rect 38268 402938 38352 403174
rect 38588 402938 38620 403174
rect 38000 402854 38620 402938
rect 38000 402618 38032 402854
rect 38268 402618 38352 402854
rect 38588 402618 38620 402854
rect 74000 402938 74032 403174
rect 74268 402938 74352 403174
rect 74588 402938 74620 403174
rect 74000 402854 74620 402938
rect 74000 402618 74032 402854
rect 74268 402618 74352 402854
rect 74588 402618 74620 402854
rect 110000 402938 110032 403174
rect 110268 402938 110352 403174
rect 110588 402938 110620 403174
rect 110000 402854 110620 402938
rect 110000 402618 110032 402854
rect 110268 402618 110352 402854
rect 110588 402618 110620 402854
rect 146000 402938 146032 403174
rect 146268 402938 146352 403174
rect 146588 402938 146620 403174
rect 146000 402854 146620 402938
rect 146000 402618 146032 402854
rect 146268 402618 146352 402854
rect 146588 402618 146620 402854
rect 182000 402938 182032 403174
rect 182268 402938 182352 403174
rect 182588 402938 182620 403174
rect 182000 402854 182620 402938
rect 182000 402618 182032 402854
rect 182268 402618 182352 402854
rect 182588 402618 182620 402854
rect 218000 402938 218032 403174
rect 218268 402938 218352 403174
rect 218588 402938 218620 403174
rect 218000 402854 218620 402938
rect 218000 402618 218032 402854
rect 218268 402618 218352 402854
rect 218588 402618 218620 402854
rect 254000 402938 254032 403174
rect 254268 402938 254352 403174
rect 254588 402938 254620 403174
rect 254000 402854 254620 402938
rect 254000 402618 254032 402854
rect 254268 402618 254352 402854
rect 254588 402618 254620 402854
rect 290000 402938 290032 403174
rect 290268 402938 290352 403174
rect 290588 402938 290620 403174
rect 290000 402854 290620 402938
rect 290000 402618 290032 402854
rect 290268 402618 290352 402854
rect 290588 402618 290620 402854
rect 326000 402938 326032 403174
rect 326268 402938 326352 403174
rect 326588 402938 326620 403174
rect 326000 402854 326620 402938
rect 326000 402618 326032 402854
rect 326268 402618 326352 402854
rect 326588 402618 326620 402854
rect 362000 402938 362032 403174
rect 362268 402938 362352 403174
rect 362588 402938 362620 403174
rect 362000 402854 362620 402938
rect 362000 402618 362032 402854
rect 362268 402618 362352 402854
rect 362588 402618 362620 402854
rect 398000 402938 398032 403174
rect 398268 402938 398352 403174
rect 398588 402938 398620 403174
rect 398000 402854 398620 402938
rect 398000 402618 398032 402854
rect 398268 402618 398352 402854
rect 398588 402618 398620 402854
rect 434000 402938 434032 403174
rect 434268 402938 434352 403174
rect 434588 402938 434620 403174
rect 434000 402854 434620 402938
rect 434000 402618 434032 402854
rect 434268 402618 434352 402854
rect 434588 402618 434620 402854
rect 470000 402938 470032 403174
rect 470268 402938 470352 403174
rect 470588 402938 470620 403174
rect 470000 402854 470620 402938
rect 470000 402618 470032 402854
rect 470268 402618 470352 402854
rect 470588 402618 470620 402854
rect 506000 402938 506032 403174
rect 506268 402938 506352 403174
rect 506588 402938 506620 403174
rect 506000 402854 506620 402938
rect 506000 402618 506032 402854
rect 506268 402618 506352 402854
rect 506588 402618 506620 402854
rect 542000 402938 542032 403174
rect 542268 402938 542352 403174
rect 542588 402938 542620 403174
rect 542000 402854 542620 402938
rect 542000 402618 542032 402854
rect 542268 402618 542352 402854
rect 542588 402618 542620 402854
rect 571500 402938 571532 403174
rect 571768 402938 571852 403174
rect 572088 402938 572120 403174
rect 571500 402854 572120 402938
rect 571500 402618 571532 402854
rect 571768 402618 571852 402854
rect 572088 402618 572120 402854
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect 9084 399218 9116 399454
rect 9352 399218 9436 399454
rect 9672 399218 9704 399454
rect 9084 399134 9704 399218
rect 9084 398898 9116 399134
rect 9352 398898 9436 399134
rect 9672 398898 9704 399134
rect 56620 399218 56652 399454
rect 56888 399218 56972 399454
rect 57208 399218 57240 399454
rect 56620 399134 57240 399218
rect 56620 398898 56652 399134
rect 56888 398898 56972 399134
rect 57208 398898 57240 399134
rect 92620 399218 92652 399454
rect 92888 399218 92972 399454
rect 93208 399218 93240 399454
rect 92620 399134 93240 399218
rect 92620 398898 92652 399134
rect 92888 398898 92972 399134
rect 93208 398898 93240 399134
rect 128620 399218 128652 399454
rect 128888 399218 128972 399454
rect 129208 399218 129240 399454
rect 128620 399134 129240 399218
rect 128620 398898 128652 399134
rect 128888 398898 128972 399134
rect 129208 398898 129240 399134
rect 164620 399218 164652 399454
rect 164888 399218 164972 399454
rect 165208 399218 165240 399454
rect 164620 399134 165240 399218
rect 164620 398898 164652 399134
rect 164888 398898 164972 399134
rect 165208 398898 165240 399134
rect 200620 399218 200652 399454
rect 200888 399218 200972 399454
rect 201208 399218 201240 399454
rect 200620 399134 201240 399218
rect 200620 398898 200652 399134
rect 200888 398898 200972 399134
rect 201208 398898 201240 399134
rect 236620 399218 236652 399454
rect 236888 399218 236972 399454
rect 237208 399218 237240 399454
rect 236620 399134 237240 399218
rect 236620 398898 236652 399134
rect 236888 398898 236972 399134
rect 237208 398898 237240 399134
rect 272620 399218 272652 399454
rect 272888 399218 272972 399454
rect 273208 399218 273240 399454
rect 272620 399134 273240 399218
rect 272620 398898 272652 399134
rect 272888 398898 272972 399134
rect 273208 398898 273240 399134
rect 308620 399218 308652 399454
rect 308888 399218 308972 399454
rect 309208 399218 309240 399454
rect 308620 399134 309240 399218
rect 308620 398898 308652 399134
rect 308888 398898 308972 399134
rect 309208 398898 309240 399134
rect 344620 399218 344652 399454
rect 344888 399218 344972 399454
rect 345208 399218 345240 399454
rect 344620 399134 345240 399218
rect 344620 398898 344652 399134
rect 344888 398898 344972 399134
rect 345208 398898 345240 399134
rect 380620 399218 380652 399454
rect 380888 399218 380972 399454
rect 381208 399218 381240 399454
rect 380620 399134 381240 399218
rect 380620 398898 380652 399134
rect 380888 398898 380972 399134
rect 381208 398898 381240 399134
rect 416620 399218 416652 399454
rect 416888 399218 416972 399454
rect 417208 399218 417240 399454
rect 416620 399134 417240 399218
rect 416620 398898 416652 399134
rect 416888 398898 416972 399134
rect 417208 398898 417240 399134
rect 452620 399218 452652 399454
rect 452888 399218 452972 399454
rect 453208 399218 453240 399454
rect 452620 399134 453240 399218
rect 452620 398898 452652 399134
rect 452888 398898 452972 399134
rect 453208 398898 453240 399134
rect 488620 399218 488652 399454
rect 488888 399218 488972 399454
rect 489208 399218 489240 399454
rect 488620 399134 489240 399218
rect 488620 398898 488652 399134
rect 488888 398898 488972 399134
rect 489208 398898 489240 399134
rect 524620 399218 524652 399454
rect 524888 399218 524972 399454
rect 525208 399218 525240 399454
rect 524620 399134 525240 399218
rect 524620 398898 524652 399134
rect 524888 398898 524972 399134
rect 525208 398898 525240 399134
rect 560620 399218 560652 399454
rect 560888 399218 560972 399454
rect 561208 399218 561240 399454
rect 560620 399134 561240 399218
rect 560620 398898 560652 399134
rect 560888 398898 560972 399134
rect 561208 398898 561240 399134
rect 570260 399218 570292 399454
rect 570528 399218 570612 399454
rect 570848 399218 570880 399454
rect 570260 399134 570880 399218
rect 570260 398898 570292 399134
rect 570528 398898 570612 399134
rect 570848 398898 570880 399134
rect -2006 363454 -1386 398898
rect 581514 367174 582134 402618
rect 7844 366938 7876 367174
rect 8112 366938 8196 367174
rect 8432 366938 8464 367174
rect 7844 366854 8464 366938
rect 7844 366618 7876 366854
rect 8112 366618 8196 366854
rect 8432 366618 8464 366854
rect 38000 366938 38032 367174
rect 38268 366938 38352 367174
rect 38588 366938 38620 367174
rect 38000 366854 38620 366938
rect 38000 366618 38032 366854
rect 38268 366618 38352 366854
rect 38588 366618 38620 366854
rect 74000 366938 74032 367174
rect 74268 366938 74352 367174
rect 74588 366938 74620 367174
rect 74000 366854 74620 366938
rect 74000 366618 74032 366854
rect 74268 366618 74352 366854
rect 74588 366618 74620 366854
rect 110000 366938 110032 367174
rect 110268 366938 110352 367174
rect 110588 366938 110620 367174
rect 110000 366854 110620 366938
rect 110000 366618 110032 366854
rect 110268 366618 110352 366854
rect 110588 366618 110620 366854
rect 146000 366938 146032 367174
rect 146268 366938 146352 367174
rect 146588 366938 146620 367174
rect 146000 366854 146620 366938
rect 146000 366618 146032 366854
rect 146268 366618 146352 366854
rect 146588 366618 146620 366854
rect 182000 366938 182032 367174
rect 182268 366938 182352 367174
rect 182588 366938 182620 367174
rect 182000 366854 182620 366938
rect 182000 366618 182032 366854
rect 182268 366618 182352 366854
rect 182588 366618 182620 366854
rect 218000 366938 218032 367174
rect 218268 366938 218352 367174
rect 218588 366938 218620 367174
rect 218000 366854 218620 366938
rect 218000 366618 218032 366854
rect 218268 366618 218352 366854
rect 218588 366618 218620 366854
rect 254000 366938 254032 367174
rect 254268 366938 254352 367174
rect 254588 366938 254620 367174
rect 254000 366854 254620 366938
rect 254000 366618 254032 366854
rect 254268 366618 254352 366854
rect 254588 366618 254620 366854
rect 290000 366938 290032 367174
rect 290268 366938 290352 367174
rect 290588 366938 290620 367174
rect 290000 366854 290620 366938
rect 290000 366618 290032 366854
rect 290268 366618 290352 366854
rect 290588 366618 290620 366854
rect 326000 366938 326032 367174
rect 326268 366938 326352 367174
rect 326588 366938 326620 367174
rect 326000 366854 326620 366938
rect 326000 366618 326032 366854
rect 326268 366618 326352 366854
rect 326588 366618 326620 366854
rect 362000 366938 362032 367174
rect 362268 366938 362352 367174
rect 362588 366938 362620 367174
rect 362000 366854 362620 366938
rect 362000 366618 362032 366854
rect 362268 366618 362352 366854
rect 362588 366618 362620 366854
rect 398000 366938 398032 367174
rect 398268 366938 398352 367174
rect 398588 366938 398620 367174
rect 398000 366854 398620 366938
rect 398000 366618 398032 366854
rect 398268 366618 398352 366854
rect 398588 366618 398620 366854
rect 434000 366938 434032 367174
rect 434268 366938 434352 367174
rect 434588 366938 434620 367174
rect 434000 366854 434620 366938
rect 434000 366618 434032 366854
rect 434268 366618 434352 366854
rect 434588 366618 434620 366854
rect 470000 366938 470032 367174
rect 470268 366938 470352 367174
rect 470588 366938 470620 367174
rect 470000 366854 470620 366938
rect 470000 366618 470032 366854
rect 470268 366618 470352 366854
rect 470588 366618 470620 366854
rect 506000 366938 506032 367174
rect 506268 366938 506352 367174
rect 506588 366938 506620 367174
rect 506000 366854 506620 366938
rect 506000 366618 506032 366854
rect 506268 366618 506352 366854
rect 506588 366618 506620 366854
rect 542000 366938 542032 367174
rect 542268 366938 542352 367174
rect 542588 366938 542620 367174
rect 542000 366854 542620 366938
rect 542000 366618 542032 366854
rect 542268 366618 542352 366854
rect 542588 366618 542620 366854
rect 571500 366938 571532 367174
rect 571768 366938 571852 367174
rect 572088 366938 572120 367174
rect 571500 366854 572120 366938
rect 571500 366618 571532 366854
rect 571768 366618 571852 366854
rect 572088 366618 572120 366854
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect 9084 363218 9116 363454
rect 9352 363218 9436 363454
rect 9672 363218 9704 363454
rect 9084 363134 9704 363218
rect 9084 362898 9116 363134
rect 9352 362898 9436 363134
rect 9672 362898 9704 363134
rect 56620 363218 56652 363454
rect 56888 363218 56972 363454
rect 57208 363218 57240 363454
rect 56620 363134 57240 363218
rect 56620 362898 56652 363134
rect 56888 362898 56972 363134
rect 57208 362898 57240 363134
rect 92620 363218 92652 363454
rect 92888 363218 92972 363454
rect 93208 363218 93240 363454
rect 92620 363134 93240 363218
rect 92620 362898 92652 363134
rect 92888 362898 92972 363134
rect 93208 362898 93240 363134
rect 128620 363218 128652 363454
rect 128888 363218 128972 363454
rect 129208 363218 129240 363454
rect 128620 363134 129240 363218
rect 128620 362898 128652 363134
rect 128888 362898 128972 363134
rect 129208 362898 129240 363134
rect 164620 363218 164652 363454
rect 164888 363218 164972 363454
rect 165208 363218 165240 363454
rect 164620 363134 165240 363218
rect 164620 362898 164652 363134
rect 164888 362898 164972 363134
rect 165208 362898 165240 363134
rect 200620 363218 200652 363454
rect 200888 363218 200972 363454
rect 201208 363218 201240 363454
rect 200620 363134 201240 363218
rect 200620 362898 200652 363134
rect 200888 362898 200972 363134
rect 201208 362898 201240 363134
rect 236620 363218 236652 363454
rect 236888 363218 236972 363454
rect 237208 363218 237240 363454
rect 236620 363134 237240 363218
rect 236620 362898 236652 363134
rect 236888 362898 236972 363134
rect 237208 362898 237240 363134
rect 272620 363218 272652 363454
rect 272888 363218 272972 363454
rect 273208 363218 273240 363454
rect 272620 363134 273240 363218
rect 272620 362898 272652 363134
rect 272888 362898 272972 363134
rect 273208 362898 273240 363134
rect 308620 363218 308652 363454
rect 308888 363218 308972 363454
rect 309208 363218 309240 363454
rect 308620 363134 309240 363218
rect 308620 362898 308652 363134
rect 308888 362898 308972 363134
rect 309208 362898 309240 363134
rect 344620 363218 344652 363454
rect 344888 363218 344972 363454
rect 345208 363218 345240 363454
rect 344620 363134 345240 363218
rect 344620 362898 344652 363134
rect 344888 362898 344972 363134
rect 345208 362898 345240 363134
rect 380620 363218 380652 363454
rect 380888 363218 380972 363454
rect 381208 363218 381240 363454
rect 380620 363134 381240 363218
rect 380620 362898 380652 363134
rect 380888 362898 380972 363134
rect 381208 362898 381240 363134
rect 416620 363218 416652 363454
rect 416888 363218 416972 363454
rect 417208 363218 417240 363454
rect 416620 363134 417240 363218
rect 416620 362898 416652 363134
rect 416888 362898 416972 363134
rect 417208 362898 417240 363134
rect 452620 363218 452652 363454
rect 452888 363218 452972 363454
rect 453208 363218 453240 363454
rect 452620 363134 453240 363218
rect 452620 362898 452652 363134
rect 452888 362898 452972 363134
rect 453208 362898 453240 363134
rect 488620 363218 488652 363454
rect 488888 363218 488972 363454
rect 489208 363218 489240 363454
rect 488620 363134 489240 363218
rect 488620 362898 488652 363134
rect 488888 362898 488972 363134
rect 489208 362898 489240 363134
rect 524620 363218 524652 363454
rect 524888 363218 524972 363454
rect 525208 363218 525240 363454
rect 524620 363134 525240 363218
rect 524620 362898 524652 363134
rect 524888 362898 524972 363134
rect 525208 362898 525240 363134
rect 560620 363218 560652 363454
rect 560888 363218 560972 363454
rect 561208 363218 561240 363454
rect 560620 363134 561240 363218
rect 560620 362898 560652 363134
rect 560888 362898 560972 363134
rect 561208 362898 561240 363134
rect 570260 363218 570292 363454
rect 570528 363218 570612 363454
rect 570848 363218 570880 363454
rect 570260 363134 570880 363218
rect 570260 362898 570292 363134
rect 570528 362898 570612 363134
rect 570848 362898 570880 363134
rect -2006 327454 -1386 362898
rect 581514 331174 582134 366618
rect 7844 330938 7876 331174
rect 8112 330938 8196 331174
rect 8432 330938 8464 331174
rect 7844 330854 8464 330938
rect 7844 330618 7876 330854
rect 8112 330618 8196 330854
rect 8432 330618 8464 330854
rect 38000 330938 38032 331174
rect 38268 330938 38352 331174
rect 38588 330938 38620 331174
rect 38000 330854 38620 330938
rect 38000 330618 38032 330854
rect 38268 330618 38352 330854
rect 38588 330618 38620 330854
rect 74000 330938 74032 331174
rect 74268 330938 74352 331174
rect 74588 330938 74620 331174
rect 74000 330854 74620 330938
rect 74000 330618 74032 330854
rect 74268 330618 74352 330854
rect 74588 330618 74620 330854
rect 110000 330938 110032 331174
rect 110268 330938 110352 331174
rect 110588 330938 110620 331174
rect 110000 330854 110620 330938
rect 110000 330618 110032 330854
rect 110268 330618 110352 330854
rect 110588 330618 110620 330854
rect 146000 330938 146032 331174
rect 146268 330938 146352 331174
rect 146588 330938 146620 331174
rect 146000 330854 146620 330938
rect 146000 330618 146032 330854
rect 146268 330618 146352 330854
rect 146588 330618 146620 330854
rect 182000 330938 182032 331174
rect 182268 330938 182352 331174
rect 182588 330938 182620 331174
rect 182000 330854 182620 330938
rect 182000 330618 182032 330854
rect 182268 330618 182352 330854
rect 182588 330618 182620 330854
rect 218000 330938 218032 331174
rect 218268 330938 218352 331174
rect 218588 330938 218620 331174
rect 218000 330854 218620 330938
rect 218000 330618 218032 330854
rect 218268 330618 218352 330854
rect 218588 330618 218620 330854
rect 254000 330938 254032 331174
rect 254268 330938 254352 331174
rect 254588 330938 254620 331174
rect 254000 330854 254620 330938
rect 254000 330618 254032 330854
rect 254268 330618 254352 330854
rect 254588 330618 254620 330854
rect 290000 330938 290032 331174
rect 290268 330938 290352 331174
rect 290588 330938 290620 331174
rect 290000 330854 290620 330938
rect 290000 330618 290032 330854
rect 290268 330618 290352 330854
rect 290588 330618 290620 330854
rect 326000 330938 326032 331174
rect 326268 330938 326352 331174
rect 326588 330938 326620 331174
rect 326000 330854 326620 330938
rect 326000 330618 326032 330854
rect 326268 330618 326352 330854
rect 326588 330618 326620 330854
rect 362000 330938 362032 331174
rect 362268 330938 362352 331174
rect 362588 330938 362620 331174
rect 362000 330854 362620 330938
rect 362000 330618 362032 330854
rect 362268 330618 362352 330854
rect 362588 330618 362620 330854
rect 398000 330938 398032 331174
rect 398268 330938 398352 331174
rect 398588 330938 398620 331174
rect 398000 330854 398620 330938
rect 398000 330618 398032 330854
rect 398268 330618 398352 330854
rect 398588 330618 398620 330854
rect 434000 330938 434032 331174
rect 434268 330938 434352 331174
rect 434588 330938 434620 331174
rect 434000 330854 434620 330938
rect 434000 330618 434032 330854
rect 434268 330618 434352 330854
rect 434588 330618 434620 330854
rect 470000 330938 470032 331174
rect 470268 330938 470352 331174
rect 470588 330938 470620 331174
rect 470000 330854 470620 330938
rect 470000 330618 470032 330854
rect 470268 330618 470352 330854
rect 470588 330618 470620 330854
rect 506000 330938 506032 331174
rect 506268 330938 506352 331174
rect 506588 330938 506620 331174
rect 506000 330854 506620 330938
rect 506000 330618 506032 330854
rect 506268 330618 506352 330854
rect 506588 330618 506620 330854
rect 542000 330938 542032 331174
rect 542268 330938 542352 331174
rect 542588 330938 542620 331174
rect 542000 330854 542620 330938
rect 542000 330618 542032 330854
rect 542268 330618 542352 330854
rect 542588 330618 542620 330854
rect 571500 330938 571532 331174
rect 571768 330938 571852 331174
rect 572088 330938 572120 331174
rect 571500 330854 572120 330938
rect 571500 330618 571532 330854
rect 571768 330618 571852 330854
rect 572088 330618 572120 330854
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect 9084 327218 9116 327454
rect 9352 327218 9436 327454
rect 9672 327218 9704 327454
rect 9084 327134 9704 327218
rect 9084 326898 9116 327134
rect 9352 326898 9436 327134
rect 9672 326898 9704 327134
rect 56620 327218 56652 327454
rect 56888 327218 56972 327454
rect 57208 327218 57240 327454
rect 56620 327134 57240 327218
rect 56620 326898 56652 327134
rect 56888 326898 56972 327134
rect 57208 326898 57240 327134
rect 92620 327218 92652 327454
rect 92888 327218 92972 327454
rect 93208 327218 93240 327454
rect 92620 327134 93240 327218
rect 92620 326898 92652 327134
rect 92888 326898 92972 327134
rect 93208 326898 93240 327134
rect 128620 327218 128652 327454
rect 128888 327218 128972 327454
rect 129208 327218 129240 327454
rect 128620 327134 129240 327218
rect 128620 326898 128652 327134
rect 128888 326898 128972 327134
rect 129208 326898 129240 327134
rect 164620 327218 164652 327454
rect 164888 327218 164972 327454
rect 165208 327218 165240 327454
rect 164620 327134 165240 327218
rect 164620 326898 164652 327134
rect 164888 326898 164972 327134
rect 165208 326898 165240 327134
rect 200620 327218 200652 327454
rect 200888 327218 200972 327454
rect 201208 327218 201240 327454
rect 200620 327134 201240 327218
rect 200620 326898 200652 327134
rect 200888 326898 200972 327134
rect 201208 326898 201240 327134
rect 236620 327218 236652 327454
rect 236888 327218 236972 327454
rect 237208 327218 237240 327454
rect 236620 327134 237240 327218
rect 236620 326898 236652 327134
rect 236888 326898 236972 327134
rect 237208 326898 237240 327134
rect 272620 327218 272652 327454
rect 272888 327218 272972 327454
rect 273208 327218 273240 327454
rect 272620 327134 273240 327218
rect 272620 326898 272652 327134
rect 272888 326898 272972 327134
rect 273208 326898 273240 327134
rect 308620 327218 308652 327454
rect 308888 327218 308972 327454
rect 309208 327218 309240 327454
rect 308620 327134 309240 327218
rect 308620 326898 308652 327134
rect 308888 326898 308972 327134
rect 309208 326898 309240 327134
rect 344620 327218 344652 327454
rect 344888 327218 344972 327454
rect 345208 327218 345240 327454
rect 344620 327134 345240 327218
rect 344620 326898 344652 327134
rect 344888 326898 344972 327134
rect 345208 326898 345240 327134
rect 380620 327218 380652 327454
rect 380888 327218 380972 327454
rect 381208 327218 381240 327454
rect 380620 327134 381240 327218
rect 380620 326898 380652 327134
rect 380888 326898 380972 327134
rect 381208 326898 381240 327134
rect 416620 327218 416652 327454
rect 416888 327218 416972 327454
rect 417208 327218 417240 327454
rect 416620 327134 417240 327218
rect 416620 326898 416652 327134
rect 416888 326898 416972 327134
rect 417208 326898 417240 327134
rect 452620 327218 452652 327454
rect 452888 327218 452972 327454
rect 453208 327218 453240 327454
rect 452620 327134 453240 327218
rect 452620 326898 452652 327134
rect 452888 326898 452972 327134
rect 453208 326898 453240 327134
rect 488620 327218 488652 327454
rect 488888 327218 488972 327454
rect 489208 327218 489240 327454
rect 488620 327134 489240 327218
rect 488620 326898 488652 327134
rect 488888 326898 488972 327134
rect 489208 326898 489240 327134
rect 524620 327218 524652 327454
rect 524888 327218 524972 327454
rect 525208 327218 525240 327454
rect 524620 327134 525240 327218
rect 524620 326898 524652 327134
rect 524888 326898 524972 327134
rect 525208 326898 525240 327134
rect 560620 327218 560652 327454
rect 560888 327218 560972 327454
rect 561208 327218 561240 327454
rect 560620 327134 561240 327218
rect 560620 326898 560652 327134
rect 560888 326898 560972 327134
rect 561208 326898 561240 327134
rect 570260 327218 570292 327454
rect 570528 327218 570612 327454
rect 570848 327218 570880 327454
rect 570260 327134 570880 327218
rect 570260 326898 570292 327134
rect 570528 326898 570612 327134
rect 570848 326898 570880 327134
rect -2006 291454 -1386 326898
rect 581514 295174 582134 330618
rect 7844 294938 7876 295174
rect 8112 294938 8196 295174
rect 8432 294938 8464 295174
rect 7844 294854 8464 294938
rect 7844 294618 7876 294854
rect 8112 294618 8196 294854
rect 8432 294618 8464 294854
rect 38000 294938 38032 295174
rect 38268 294938 38352 295174
rect 38588 294938 38620 295174
rect 38000 294854 38620 294938
rect 38000 294618 38032 294854
rect 38268 294618 38352 294854
rect 38588 294618 38620 294854
rect 74000 294938 74032 295174
rect 74268 294938 74352 295174
rect 74588 294938 74620 295174
rect 74000 294854 74620 294938
rect 74000 294618 74032 294854
rect 74268 294618 74352 294854
rect 74588 294618 74620 294854
rect 110000 294938 110032 295174
rect 110268 294938 110352 295174
rect 110588 294938 110620 295174
rect 110000 294854 110620 294938
rect 110000 294618 110032 294854
rect 110268 294618 110352 294854
rect 110588 294618 110620 294854
rect 146000 294938 146032 295174
rect 146268 294938 146352 295174
rect 146588 294938 146620 295174
rect 146000 294854 146620 294938
rect 146000 294618 146032 294854
rect 146268 294618 146352 294854
rect 146588 294618 146620 294854
rect 182000 294938 182032 295174
rect 182268 294938 182352 295174
rect 182588 294938 182620 295174
rect 182000 294854 182620 294938
rect 182000 294618 182032 294854
rect 182268 294618 182352 294854
rect 182588 294618 182620 294854
rect 218000 294938 218032 295174
rect 218268 294938 218352 295174
rect 218588 294938 218620 295174
rect 218000 294854 218620 294938
rect 218000 294618 218032 294854
rect 218268 294618 218352 294854
rect 218588 294618 218620 294854
rect 254000 294938 254032 295174
rect 254268 294938 254352 295174
rect 254588 294938 254620 295174
rect 254000 294854 254620 294938
rect 254000 294618 254032 294854
rect 254268 294618 254352 294854
rect 254588 294618 254620 294854
rect 290000 294938 290032 295174
rect 290268 294938 290352 295174
rect 290588 294938 290620 295174
rect 290000 294854 290620 294938
rect 290000 294618 290032 294854
rect 290268 294618 290352 294854
rect 290588 294618 290620 294854
rect 326000 294938 326032 295174
rect 326268 294938 326352 295174
rect 326588 294938 326620 295174
rect 326000 294854 326620 294938
rect 326000 294618 326032 294854
rect 326268 294618 326352 294854
rect 326588 294618 326620 294854
rect 362000 294938 362032 295174
rect 362268 294938 362352 295174
rect 362588 294938 362620 295174
rect 362000 294854 362620 294938
rect 362000 294618 362032 294854
rect 362268 294618 362352 294854
rect 362588 294618 362620 294854
rect 398000 294938 398032 295174
rect 398268 294938 398352 295174
rect 398588 294938 398620 295174
rect 398000 294854 398620 294938
rect 398000 294618 398032 294854
rect 398268 294618 398352 294854
rect 398588 294618 398620 294854
rect 434000 294938 434032 295174
rect 434268 294938 434352 295174
rect 434588 294938 434620 295174
rect 434000 294854 434620 294938
rect 434000 294618 434032 294854
rect 434268 294618 434352 294854
rect 434588 294618 434620 294854
rect 470000 294938 470032 295174
rect 470268 294938 470352 295174
rect 470588 294938 470620 295174
rect 470000 294854 470620 294938
rect 470000 294618 470032 294854
rect 470268 294618 470352 294854
rect 470588 294618 470620 294854
rect 506000 294938 506032 295174
rect 506268 294938 506352 295174
rect 506588 294938 506620 295174
rect 506000 294854 506620 294938
rect 506000 294618 506032 294854
rect 506268 294618 506352 294854
rect 506588 294618 506620 294854
rect 542000 294938 542032 295174
rect 542268 294938 542352 295174
rect 542588 294938 542620 295174
rect 542000 294854 542620 294938
rect 542000 294618 542032 294854
rect 542268 294618 542352 294854
rect 542588 294618 542620 294854
rect 571500 294938 571532 295174
rect 571768 294938 571852 295174
rect 572088 294938 572120 295174
rect 571500 294854 572120 294938
rect 571500 294618 571532 294854
rect 571768 294618 571852 294854
rect 572088 294618 572120 294854
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect 9084 291218 9116 291454
rect 9352 291218 9436 291454
rect 9672 291218 9704 291454
rect 9084 291134 9704 291218
rect 9084 290898 9116 291134
rect 9352 290898 9436 291134
rect 9672 290898 9704 291134
rect 56620 291218 56652 291454
rect 56888 291218 56972 291454
rect 57208 291218 57240 291454
rect 56620 291134 57240 291218
rect 56620 290898 56652 291134
rect 56888 290898 56972 291134
rect 57208 290898 57240 291134
rect 92620 291218 92652 291454
rect 92888 291218 92972 291454
rect 93208 291218 93240 291454
rect 92620 291134 93240 291218
rect 92620 290898 92652 291134
rect 92888 290898 92972 291134
rect 93208 290898 93240 291134
rect 128620 291218 128652 291454
rect 128888 291218 128972 291454
rect 129208 291218 129240 291454
rect 128620 291134 129240 291218
rect 128620 290898 128652 291134
rect 128888 290898 128972 291134
rect 129208 290898 129240 291134
rect 164620 291218 164652 291454
rect 164888 291218 164972 291454
rect 165208 291218 165240 291454
rect 164620 291134 165240 291218
rect 164620 290898 164652 291134
rect 164888 290898 164972 291134
rect 165208 290898 165240 291134
rect 200620 291218 200652 291454
rect 200888 291218 200972 291454
rect 201208 291218 201240 291454
rect 200620 291134 201240 291218
rect 200620 290898 200652 291134
rect 200888 290898 200972 291134
rect 201208 290898 201240 291134
rect 236620 291218 236652 291454
rect 236888 291218 236972 291454
rect 237208 291218 237240 291454
rect 236620 291134 237240 291218
rect 236620 290898 236652 291134
rect 236888 290898 236972 291134
rect 237208 290898 237240 291134
rect 272620 291218 272652 291454
rect 272888 291218 272972 291454
rect 273208 291218 273240 291454
rect 272620 291134 273240 291218
rect 272620 290898 272652 291134
rect 272888 290898 272972 291134
rect 273208 290898 273240 291134
rect 308620 291218 308652 291454
rect 308888 291218 308972 291454
rect 309208 291218 309240 291454
rect 308620 291134 309240 291218
rect 308620 290898 308652 291134
rect 308888 290898 308972 291134
rect 309208 290898 309240 291134
rect 344620 291218 344652 291454
rect 344888 291218 344972 291454
rect 345208 291218 345240 291454
rect 344620 291134 345240 291218
rect 344620 290898 344652 291134
rect 344888 290898 344972 291134
rect 345208 290898 345240 291134
rect 380620 291218 380652 291454
rect 380888 291218 380972 291454
rect 381208 291218 381240 291454
rect 380620 291134 381240 291218
rect 380620 290898 380652 291134
rect 380888 290898 380972 291134
rect 381208 290898 381240 291134
rect 416620 291218 416652 291454
rect 416888 291218 416972 291454
rect 417208 291218 417240 291454
rect 416620 291134 417240 291218
rect 416620 290898 416652 291134
rect 416888 290898 416972 291134
rect 417208 290898 417240 291134
rect 452620 291218 452652 291454
rect 452888 291218 452972 291454
rect 453208 291218 453240 291454
rect 452620 291134 453240 291218
rect 452620 290898 452652 291134
rect 452888 290898 452972 291134
rect 453208 290898 453240 291134
rect 488620 291218 488652 291454
rect 488888 291218 488972 291454
rect 489208 291218 489240 291454
rect 488620 291134 489240 291218
rect 488620 290898 488652 291134
rect 488888 290898 488972 291134
rect 489208 290898 489240 291134
rect 524620 291218 524652 291454
rect 524888 291218 524972 291454
rect 525208 291218 525240 291454
rect 524620 291134 525240 291218
rect 524620 290898 524652 291134
rect 524888 290898 524972 291134
rect 525208 290898 525240 291134
rect 560620 291218 560652 291454
rect 560888 291218 560972 291454
rect 561208 291218 561240 291454
rect 560620 291134 561240 291218
rect 560620 290898 560652 291134
rect 560888 290898 560972 291134
rect 561208 290898 561240 291134
rect 570260 291218 570292 291454
rect 570528 291218 570612 291454
rect 570848 291218 570880 291454
rect 570260 291134 570880 291218
rect 570260 290898 570292 291134
rect 570528 290898 570612 291134
rect 570848 290898 570880 291134
rect -2006 255454 -1386 290898
rect 581514 259174 582134 294618
rect 7844 258938 7876 259174
rect 8112 258938 8196 259174
rect 8432 258938 8464 259174
rect 7844 258854 8464 258938
rect 7844 258618 7876 258854
rect 8112 258618 8196 258854
rect 8432 258618 8464 258854
rect 38000 258938 38032 259174
rect 38268 258938 38352 259174
rect 38588 258938 38620 259174
rect 38000 258854 38620 258938
rect 38000 258618 38032 258854
rect 38268 258618 38352 258854
rect 38588 258618 38620 258854
rect 74000 258938 74032 259174
rect 74268 258938 74352 259174
rect 74588 258938 74620 259174
rect 74000 258854 74620 258938
rect 74000 258618 74032 258854
rect 74268 258618 74352 258854
rect 74588 258618 74620 258854
rect 110000 258938 110032 259174
rect 110268 258938 110352 259174
rect 110588 258938 110620 259174
rect 110000 258854 110620 258938
rect 110000 258618 110032 258854
rect 110268 258618 110352 258854
rect 110588 258618 110620 258854
rect 146000 258938 146032 259174
rect 146268 258938 146352 259174
rect 146588 258938 146620 259174
rect 146000 258854 146620 258938
rect 146000 258618 146032 258854
rect 146268 258618 146352 258854
rect 146588 258618 146620 258854
rect 182000 258938 182032 259174
rect 182268 258938 182352 259174
rect 182588 258938 182620 259174
rect 182000 258854 182620 258938
rect 182000 258618 182032 258854
rect 182268 258618 182352 258854
rect 182588 258618 182620 258854
rect 218000 258938 218032 259174
rect 218268 258938 218352 259174
rect 218588 258938 218620 259174
rect 218000 258854 218620 258938
rect 218000 258618 218032 258854
rect 218268 258618 218352 258854
rect 218588 258618 218620 258854
rect 254000 258938 254032 259174
rect 254268 258938 254352 259174
rect 254588 258938 254620 259174
rect 254000 258854 254620 258938
rect 254000 258618 254032 258854
rect 254268 258618 254352 258854
rect 254588 258618 254620 258854
rect 290000 258938 290032 259174
rect 290268 258938 290352 259174
rect 290588 258938 290620 259174
rect 290000 258854 290620 258938
rect 290000 258618 290032 258854
rect 290268 258618 290352 258854
rect 290588 258618 290620 258854
rect 326000 258938 326032 259174
rect 326268 258938 326352 259174
rect 326588 258938 326620 259174
rect 326000 258854 326620 258938
rect 326000 258618 326032 258854
rect 326268 258618 326352 258854
rect 326588 258618 326620 258854
rect 362000 258938 362032 259174
rect 362268 258938 362352 259174
rect 362588 258938 362620 259174
rect 362000 258854 362620 258938
rect 362000 258618 362032 258854
rect 362268 258618 362352 258854
rect 362588 258618 362620 258854
rect 398000 258938 398032 259174
rect 398268 258938 398352 259174
rect 398588 258938 398620 259174
rect 398000 258854 398620 258938
rect 398000 258618 398032 258854
rect 398268 258618 398352 258854
rect 398588 258618 398620 258854
rect 434000 258938 434032 259174
rect 434268 258938 434352 259174
rect 434588 258938 434620 259174
rect 434000 258854 434620 258938
rect 434000 258618 434032 258854
rect 434268 258618 434352 258854
rect 434588 258618 434620 258854
rect 470000 258938 470032 259174
rect 470268 258938 470352 259174
rect 470588 258938 470620 259174
rect 470000 258854 470620 258938
rect 470000 258618 470032 258854
rect 470268 258618 470352 258854
rect 470588 258618 470620 258854
rect 506000 258938 506032 259174
rect 506268 258938 506352 259174
rect 506588 258938 506620 259174
rect 506000 258854 506620 258938
rect 506000 258618 506032 258854
rect 506268 258618 506352 258854
rect 506588 258618 506620 258854
rect 542000 258938 542032 259174
rect 542268 258938 542352 259174
rect 542588 258938 542620 259174
rect 542000 258854 542620 258938
rect 542000 258618 542032 258854
rect 542268 258618 542352 258854
rect 542588 258618 542620 258854
rect 571500 258938 571532 259174
rect 571768 258938 571852 259174
rect 572088 258938 572120 259174
rect 571500 258854 572120 258938
rect 571500 258618 571532 258854
rect 571768 258618 571852 258854
rect 572088 258618 572120 258854
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect 9084 255218 9116 255454
rect 9352 255218 9436 255454
rect 9672 255218 9704 255454
rect 9084 255134 9704 255218
rect 9084 254898 9116 255134
rect 9352 254898 9436 255134
rect 9672 254898 9704 255134
rect 56620 255218 56652 255454
rect 56888 255218 56972 255454
rect 57208 255218 57240 255454
rect 56620 255134 57240 255218
rect 56620 254898 56652 255134
rect 56888 254898 56972 255134
rect 57208 254898 57240 255134
rect 92620 255218 92652 255454
rect 92888 255218 92972 255454
rect 93208 255218 93240 255454
rect 92620 255134 93240 255218
rect 92620 254898 92652 255134
rect 92888 254898 92972 255134
rect 93208 254898 93240 255134
rect 128620 255218 128652 255454
rect 128888 255218 128972 255454
rect 129208 255218 129240 255454
rect 128620 255134 129240 255218
rect 128620 254898 128652 255134
rect 128888 254898 128972 255134
rect 129208 254898 129240 255134
rect 164620 255218 164652 255454
rect 164888 255218 164972 255454
rect 165208 255218 165240 255454
rect 164620 255134 165240 255218
rect 164620 254898 164652 255134
rect 164888 254898 164972 255134
rect 165208 254898 165240 255134
rect 200620 255218 200652 255454
rect 200888 255218 200972 255454
rect 201208 255218 201240 255454
rect 200620 255134 201240 255218
rect 200620 254898 200652 255134
rect 200888 254898 200972 255134
rect 201208 254898 201240 255134
rect 236620 255218 236652 255454
rect 236888 255218 236972 255454
rect 237208 255218 237240 255454
rect 236620 255134 237240 255218
rect 236620 254898 236652 255134
rect 236888 254898 236972 255134
rect 237208 254898 237240 255134
rect 272620 255218 272652 255454
rect 272888 255218 272972 255454
rect 273208 255218 273240 255454
rect 272620 255134 273240 255218
rect 272620 254898 272652 255134
rect 272888 254898 272972 255134
rect 273208 254898 273240 255134
rect 308620 255218 308652 255454
rect 308888 255218 308972 255454
rect 309208 255218 309240 255454
rect 308620 255134 309240 255218
rect 308620 254898 308652 255134
rect 308888 254898 308972 255134
rect 309208 254898 309240 255134
rect 344620 255218 344652 255454
rect 344888 255218 344972 255454
rect 345208 255218 345240 255454
rect 344620 255134 345240 255218
rect 344620 254898 344652 255134
rect 344888 254898 344972 255134
rect 345208 254898 345240 255134
rect 380620 255218 380652 255454
rect 380888 255218 380972 255454
rect 381208 255218 381240 255454
rect 380620 255134 381240 255218
rect 380620 254898 380652 255134
rect 380888 254898 380972 255134
rect 381208 254898 381240 255134
rect 416620 255218 416652 255454
rect 416888 255218 416972 255454
rect 417208 255218 417240 255454
rect 416620 255134 417240 255218
rect 416620 254898 416652 255134
rect 416888 254898 416972 255134
rect 417208 254898 417240 255134
rect 452620 255218 452652 255454
rect 452888 255218 452972 255454
rect 453208 255218 453240 255454
rect 452620 255134 453240 255218
rect 452620 254898 452652 255134
rect 452888 254898 452972 255134
rect 453208 254898 453240 255134
rect 488620 255218 488652 255454
rect 488888 255218 488972 255454
rect 489208 255218 489240 255454
rect 488620 255134 489240 255218
rect 488620 254898 488652 255134
rect 488888 254898 488972 255134
rect 489208 254898 489240 255134
rect 524620 255218 524652 255454
rect 524888 255218 524972 255454
rect 525208 255218 525240 255454
rect 524620 255134 525240 255218
rect 524620 254898 524652 255134
rect 524888 254898 524972 255134
rect 525208 254898 525240 255134
rect 560620 255218 560652 255454
rect 560888 255218 560972 255454
rect 561208 255218 561240 255454
rect 560620 255134 561240 255218
rect 560620 254898 560652 255134
rect 560888 254898 560972 255134
rect 561208 254898 561240 255134
rect 570260 255218 570292 255454
rect 570528 255218 570612 255454
rect 570848 255218 570880 255454
rect 570260 255134 570880 255218
rect 570260 254898 570292 255134
rect 570528 254898 570612 255134
rect 570848 254898 570880 255134
rect -2006 219454 -1386 254898
rect 581514 223174 582134 258618
rect 7844 222938 7876 223174
rect 8112 222938 8196 223174
rect 8432 222938 8464 223174
rect 7844 222854 8464 222938
rect 7844 222618 7876 222854
rect 8112 222618 8196 222854
rect 8432 222618 8464 222854
rect 38000 222938 38032 223174
rect 38268 222938 38352 223174
rect 38588 222938 38620 223174
rect 38000 222854 38620 222938
rect 38000 222618 38032 222854
rect 38268 222618 38352 222854
rect 38588 222618 38620 222854
rect 74000 222938 74032 223174
rect 74268 222938 74352 223174
rect 74588 222938 74620 223174
rect 74000 222854 74620 222938
rect 74000 222618 74032 222854
rect 74268 222618 74352 222854
rect 74588 222618 74620 222854
rect 110000 222938 110032 223174
rect 110268 222938 110352 223174
rect 110588 222938 110620 223174
rect 110000 222854 110620 222938
rect 110000 222618 110032 222854
rect 110268 222618 110352 222854
rect 110588 222618 110620 222854
rect 146000 222938 146032 223174
rect 146268 222938 146352 223174
rect 146588 222938 146620 223174
rect 146000 222854 146620 222938
rect 146000 222618 146032 222854
rect 146268 222618 146352 222854
rect 146588 222618 146620 222854
rect 182000 222938 182032 223174
rect 182268 222938 182352 223174
rect 182588 222938 182620 223174
rect 182000 222854 182620 222938
rect 182000 222618 182032 222854
rect 182268 222618 182352 222854
rect 182588 222618 182620 222854
rect 218000 222938 218032 223174
rect 218268 222938 218352 223174
rect 218588 222938 218620 223174
rect 218000 222854 218620 222938
rect 218000 222618 218032 222854
rect 218268 222618 218352 222854
rect 218588 222618 218620 222854
rect 254000 222938 254032 223174
rect 254268 222938 254352 223174
rect 254588 222938 254620 223174
rect 254000 222854 254620 222938
rect 254000 222618 254032 222854
rect 254268 222618 254352 222854
rect 254588 222618 254620 222854
rect 290000 222938 290032 223174
rect 290268 222938 290352 223174
rect 290588 222938 290620 223174
rect 290000 222854 290620 222938
rect 290000 222618 290032 222854
rect 290268 222618 290352 222854
rect 290588 222618 290620 222854
rect 326000 222938 326032 223174
rect 326268 222938 326352 223174
rect 326588 222938 326620 223174
rect 326000 222854 326620 222938
rect 326000 222618 326032 222854
rect 326268 222618 326352 222854
rect 326588 222618 326620 222854
rect 362000 222938 362032 223174
rect 362268 222938 362352 223174
rect 362588 222938 362620 223174
rect 362000 222854 362620 222938
rect 362000 222618 362032 222854
rect 362268 222618 362352 222854
rect 362588 222618 362620 222854
rect 398000 222938 398032 223174
rect 398268 222938 398352 223174
rect 398588 222938 398620 223174
rect 398000 222854 398620 222938
rect 398000 222618 398032 222854
rect 398268 222618 398352 222854
rect 398588 222618 398620 222854
rect 434000 222938 434032 223174
rect 434268 222938 434352 223174
rect 434588 222938 434620 223174
rect 434000 222854 434620 222938
rect 434000 222618 434032 222854
rect 434268 222618 434352 222854
rect 434588 222618 434620 222854
rect 470000 222938 470032 223174
rect 470268 222938 470352 223174
rect 470588 222938 470620 223174
rect 470000 222854 470620 222938
rect 470000 222618 470032 222854
rect 470268 222618 470352 222854
rect 470588 222618 470620 222854
rect 506000 222938 506032 223174
rect 506268 222938 506352 223174
rect 506588 222938 506620 223174
rect 506000 222854 506620 222938
rect 506000 222618 506032 222854
rect 506268 222618 506352 222854
rect 506588 222618 506620 222854
rect 542000 222938 542032 223174
rect 542268 222938 542352 223174
rect 542588 222938 542620 223174
rect 542000 222854 542620 222938
rect 542000 222618 542032 222854
rect 542268 222618 542352 222854
rect 542588 222618 542620 222854
rect 571500 222938 571532 223174
rect 571768 222938 571852 223174
rect 572088 222938 572120 223174
rect 571500 222854 572120 222938
rect 571500 222618 571532 222854
rect 571768 222618 571852 222854
rect 572088 222618 572120 222854
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect 9084 219218 9116 219454
rect 9352 219218 9436 219454
rect 9672 219218 9704 219454
rect 9084 219134 9704 219218
rect 9084 218898 9116 219134
rect 9352 218898 9436 219134
rect 9672 218898 9704 219134
rect 56620 219218 56652 219454
rect 56888 219218 56972 219454
rect 57208 219218 57240 219454
rect 56620 219134 57240 219218
rect 56620 218898 56652 219134
rect 56888 218898 56972 219134
rect 57208 218898 57240 219134
rect 92620 219218 92652 219454
rect 92888 219218 92972 219454
rect 93208 219218 93240 219454
rect 92620 219134 93240 219218
rect 92620 218898 92652 219134
rect 92888 218898 92972 219134
rect 93208 218898 93240 219134
rect 128620 219218 128652 219454
rect 128888 219218 128972 219454
rect 129208 219218 129240 219454
rect 128620 219134 129240 219218
rect 128620 218898 128652 219134
rect 128888 218898 128972 219134
rect 129208 218898 129240 219134
rect 164620 219218 164652 219454
rect 164888 219218 164972 219454
rect 165208 219218 165240 219454
rect 164620 219134 165240 219218
rect 164620 218898 164652 219134
rect 164888 218898 164972 219134
rect 165208 218898 165240 219134
rect 200620 219218 200652 219454
rect 200888 219218 200972 219454
rect 201208 219218 201240 219454
rect 200620 219134 201240 219218
rect 200620 218898 200652 219134
rect 200888 218898 200972 219134
rect 201208 218898 201240 219134
rect 236620 219218 236652 219454
rect 236888 219218 236972 219454
rect 237208 219218 237240 219454
rect 236620 219134 237240 219218
rect 236620 218898 236652 219134
rect 236888 218898 236972 219134
rect 237208 218898 237240 219134
rect 272620 219218 272652 219454
rect 272888 219218 272972 219454
rect 273208 219218 273240 219454
rect 272620 219134 273240 219218
rect 272620 218898 272652 219134
rect 272888 218898 272972 219134
rect 273208 218898 273240 219134
rect 308620 219218 308652 219454
rect 308888 219218 308972 219454
rect 309208 219218 309240 219454
rect 308620 219134 309240 219218
rect 308620 218898 308652 219134
rect 308888 218898 308972 219134
rect 309208 218898 309240 219134
rect 344620 219218 344652 219454
rect 344888 219218 344972 219454
rect 345208 219218 345240 219454
rect 344620 219134 345240 219218
rect 344620 218898 344652 219134
rect 344888 218898 344972 219134
rect 345208 218898 345240 219134
rect 380620 219218 380652 219454
rect 380888 219218 380972 219454
rect 381208 219218 381240 219454
rect 380620 219134 381240 219218
rect 380620 218898 380652 219134
rect 380888 218898 380972 219134
rect 381208 218898 381240 219134
rect 416620 219218 416652 219454
rect 416888 219218 416972 219454
rect 417208 219218 417240 219454
rect 416620 219134 417240 219218
rect 416620 218898 416652 219134
rect 416888 218898 416972 219134
rect 417208 218898 417240 219134
rect 452620 219218 452652 219454
rect 452888 219218 452972 219454
rect 453208 219218 453240 219454
rect 452620 219134 453240 219218
rect 452620 218898 452652 219134
rect 452888 218898 452972 219134
rect 453208 218898 453240 219134
rect 488620 219218 488652 219454
rect 488888 219218 488972 219454
rect 489208 219218 489240 219454
rect 488620 219134 489240 219218
rect 488620 218898 488652 219134
rect 488888 218898 488972 219134
rect 489208 218898 489240 219134
rect 524620 219218 524652 219454
rect 524888 219218 524972 219454
rect 525208 219218 525240 219454
rect 524620 219134 525240 219218
rect 524620 218898 524652 219134
rect 524888 218898 524972 219134
rect 525208 218898 525240 219134
rect 560620 219218 560652 219454
rect 560888 219218 560972 219454
rect 561208 219218 561240 219454
rect 560620 219134 561240 219218
rect 560620 218898 560652 219134
rect 560888 218898 560972 219134
rect 561208 218898 561240 219134
rect 570260 219218 570292 219454
rect 570528 219218 570612 219454
rect 570848 219218 570880 219454
rect 570260 219134 570880 219218
rect 570260 218898 570292 219134
rect 570528 218898 570612 219134
rect 570848 218898 570880 219134
rect -2006 183454 -1386 218898
rect 60560 187174 60920 187206
rect 7844 186938 7876 187174
rect 8112 186938 8196 187174
rect 8432 186938 8464 187174
rect 7844 186854 8464 186938
rect 7844 186618 7876 186854
rect 8112 186618 8196 186854
rect 8432 186618 8464 186854
rect 38000 186938 38032 187174
rect 38268 186938 38352 187174
rect 38588 186938 38620 187174
rect 38000 186854 38620 186938
rect 38000 186618 38032 186854
rect 38268 186618 38352 186854
rect 38588 186618 38620 186854
rect 60560 186938 60622 187174
rect 60858 186938 60920 187174
rect 60560 186854 60920 186938
rect 60560 186618 60622 186854
rect 60858 186618 60920 186854
rect 60560 186586 60920 186618
rect 159036 187174 159396 187206
rect 185560 187174 185920 187206
rect 159036 186938 159098 187174
rect 159334 186938 159396 187174
rect 159036 186854 159396 186938
rect 159036 186618 159098 186854
rect 159334 186618 159396 186854
rect 182000 186938 182032 187174
rect 182268 186938 182352 187174
rect 182588 186938 182620 187174
rect 182000 186854 182620 186938
rect 182000 186618 182032 186854
rect 182268 186618 182352 186854
rect 182588 186618 182620 186854
rect 185560 186938 185622 187174
rect 185858 186938 185920 187174
rect 185560 186854 185920 186938
rect 185560 186618 185622 186854
rect 185858 186618 185920 186854
rect 159036 186586 159396 186618
rect 185560 186586 185920 186618
rect 284036 187174 284396 187206
rect 310560 187174 310920 187206
rect 284036 186938 284098 187174
rect 284334 186938 284396 187174
rect 284036 186854 284396 186938
rect 284036 186618 284098 186854
rect 284334 186618 284396 186854
rect 290000 186938 290032 187174
rect 290268 186938 290352 187174
rect 290588 186938 290620 187174
rect 290000 186854 290620 186938
rect 290000 186618 290032 186854
rect 290268 186618 290352 186854
rect 290588 186618 290620 186854
rect 310560 186938 310622 187174
rect 310858 186938 310920 187174
rect 310560 186854 310920 186938
rect 310560 186618 310622 186854
rect 310858 186618 310920 186854
rect 284036 186586 284396 186618
rect 310560 186586 310920 186618
rect 409036 187174 409396 187206
rect 436560 187174 436920 187206
rect 409036 186938 409098 187174
rect 409334 186938 409396 187174
rect 409036 186854 409396 186938
rect 409036 186618 409098 186854
rect 409334 186618 409396 186854
rect 434000 186938 434032 187174
rect 434268 186938 434352 187174
rect 434588 186938 434620 187174
rect 434000 186854 434620 186938
rect 434000 186618 434032 186854
rect 434268 186618 434352 186854
rect 434588 186618 434620 186854
rect 436560 186938 436622 187174
rect 436858 186938 436920 187174
rect 436560 186854 436920 186938
rect 436560 186618 436622 186854
rect 436858 186618 436920 186854
rect 409036 186586 409396 186618
rect 436560 186586 436920 186618
rect 535036 187174 535396 187206
rect 581514 187174 582134 222618
rect 535036 186938 535098 187174
rect 535334 186938 535396 187174
rect 535036 186854 535396 186938
rect 535036 186618 535098 186854
rect 535334 186618 535396 186854
rect 542000 186938 542032 187174
rect 542268 186938 542352 187174
rect 542588 186938 542620 187174
rect 542000 186854 542620 186938
rect 542000 186618 542032 186854
rect 542268 186618 542352 186854
rect 542588 186618 542620 186854
rect 571500 186938 571532 187174
rect 571768 186938 571852 187174
rect 572088 186938 572120 187174
rect 571500 186854 572120 186938
rect 571500 186618 571532 186854
rect 571768 186618 571852 186854
rect 572088 186618 572120 186854
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 535036 186586 535396 186618
rect 61280 183454 61640 183486
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect 9084 183218 9116 183454
rect 9352 183218 9436 183454
rect 9672 183218 9704 183454
rect 9084 183134 9704 183218
rect 9084 182898 9116 183134
rect 9352 182898 9436 183134
rect 9672 182898 9704 183134
rect 56620 183218 56652 183454
rect 56888 183218 56972 183454
rect 57208 183218 57240 183454
rect 56620 183134 57240 183218
rect 56620 182898 56652 183134
rect 56888 182898 56972 183134
rect 57208 182898 57240 183134
rect 61280 183218 61342 183454
rect 61578 183218 61640 183454
rect 61280 183134 61640 183218
rect 61280 182898 61342 183134
rect 61578 182898 61640 183134
rect -2006 147454 -1386 182898
rect 61280 182866 61640 182898
rect 158316 183454 158676 183486
rect 186280 183454 186640 183486
rect 158316 183218 158378 183454
rect 158614 183218 158676 183454
rect 158316 183134 158676 183218
rect 158316 182898 158378 183134
rect 158614 182898 158676 183134
rect 164620 183218 164652 183454
rect 164888 183218 164972 183454
rect 165208 183218 165240 183454
rect 164620 183134 165240 183218
rect 164620 182898 164652 183134
rect 164888 182898 164972 183134
rect 165208 182898 165240 183134
rect 186280 183218 186342 183454
rect 186578 183218 186640 183454
rect 186280 183134 186640 183218
rect 186280 182898 186342 183134
rect 186578 182898 186640 183134
rect 158316 182866 158676 182898
rect 186280 182866 186640 182898
rect 283316 183454 283676 183486
rect 311280 183454 311640 183486
rect 283316 183218 283378 183454
rect 283614 183218 283676 183454
rect 283316 183134 283676 183218
rect 283316 182898 283378 183134
rect 283614 182898 283676 183134
rect 308620 183218 308652 183454
rect 308888 183218 308972 183454
rect 309208 183218 309240 183454
rect 308620 183134 309240 183218
rect 308620 182898 308652 183134
rect 308888 182898 308972 183134
rect 309208 182898 309240 183134
rect 311280 183218 311342 183454
rect 311578 183218 311640 183454
rect 311280 183134 311640 183218
rect 311280 182898 311342 183134
rect 311578 182898 311640 183134
rect 283316 182866 283676 182898
rect 311280 182866 311640 182898
rect 408316 183454 408676 183486
rect 437280 183454 437640 183486
rect 408316 183218 408378 183454
rect 408614 183218 408676 183454
rect 408316 183134 408676 183218
rect 408316 182898 408378 183134
rect 408614 182898 408676 183134
rect 416620 183218 416652 183454
rect 416888 183218 416972 183454
rect 417208 183218 417240 183454
rect 416620 183134 417240 183218
rect 416620 182898 416652 183134
rect 416888 182898 416972 183134
rect 417208 182898 417240 183134
rect 437280 183218 437342 183454
rect 437578 183218 437640 183454
rect 437280 183134 437640 183218
rect 437280 182898 437342 183134
rect 437578 182898 437640 183134
rect 408316 182866 408676 182898
rect 437280 182866 437640 182898
rect 534316 183454 534676 183486
rect 534316 183218 534378 183454
rect 534614 183218 534676 183454
rect 534316 183134 534676 183218
rect 534316 182898 534378 183134
rect 534614 182898 534676 183134
rect 560620 183218 560652 183454
rect 560888 183218 560972 183454
rect 561208 183218 561240 183454
rect 560620 183134 561240 183218
rect 560620 182898 560652 183134
rect 560888 182898 560972 183134
rect 561208 182898 561240 183134
rect 570260 183218 570292 183454
rect 570528 183218 570612 183454
rect 570848 183218 570880 183454
rect 570260 183134 570880 183218
rect 570260 182898 570292 183134
rect 570528 182898 570612 183134
rect 570848 182898 570880 183134
rect 534316 182866 534676 182898
rect 60560 151174 60920 151206
rect 7844 150938 7876 151174
rect 8112 150938 8196 151174
rect 8432 150938 8464 151174
rect 7844 150854 8464 150938
rect 7844 150618 7876 150854
rect 8112 150618 8196 150854
rect 8432 150618 8464 150854
rect 38000 150938 38032 151174
rect 38268 150938 38352 151174
rect 38588 150938 38620 151174
rect 38000 150854 38620 150938
rect 38000 150618 38032 150854
rect 38268 150618 38352 150854
rect 38588 150618 38620 150854
rect 60560 150938 60622 151174
rect 60858 150938 60920 151174
rect 60560 150854 60920 150938
rect 60560 150618 60622 150854
rect 60858 150618 60920 150854
rect 60560 150586 60920 150618
rect 159036 151174 159396 151206
rect 185560 151174 185920 151206
rect 159036 150938 159098 151174
rect 159334 150938 159396 151174
rect 159036 150854 159396 150938
rect 159036 150618 159098 150854
rect 159334 150618 159396 150854
rect 182000 150938 182032 151174
rect 182268 150938 182352 151174
rect 182588 150938 182620 151174
rect 182000 150854 182620 150938
rect 182000 150618 182032 150854
rect 182268 150618 182352 150854
rect 182588 150618 182620 150854
rect 185560 150938 185622 151174
rect 185858 150938 185920 151174
rect 185560 150854 185920 150938
rect 185560 150618 185622 150854
rect 185858 150618 185920 150854
rect 159036 150586 159396 150618
rect 185560 150586 185920 150618
rect 284036 151174 284396 151206
rect 310560 151174 310920 151206
rect 284036 150938 284098 151174
rect 284334 150938 284396 151174
rect 284036 150854 284396 150938
rect 284036 150618 284098 150854
rect 284334 150618 284396 150854
rect 290000 150938 290032 151174
rect 290268 150938 290352 151174
rect 290588 150938 290620 151174
rect 290000 150854 290620 150938
rect 290000 150618 290032 150854
rect 290268 150618 290352 150854
rect 290588 150618 290620 150854
rect 310560 150938 310622 151174
rect 310858 150938 310920 151174
rect 310560 150854 310920 150938
rect 310560 150618 310622 150854
rect 310858 150618 310920 150854
rect 284036 150586 284396 150618
rect 310560 150586 310920 150618
rect 409036 151174 409396 151206
rect 436560 151174 436920 151206
rect 409036 150938 409098 151174
rect 409334 150938 409396 151174
rect 409036 150854 409396 150938
rect 409036 150618 409098 150854
rect 409334 150618 409396 150854
rect 434000 150938 434032 151174
rect 434268 150938 434352 151174
rect 434588 150938 434620 151174
rect 434000 150854 434620 150938
rect 434000 150618 434032 150854
rect 434268 150618 434352 150854
rect 434588 150618 434620 150854
rect 436560 150938 436622 151174
rect 436858 150938 436920 151174
rect 436560 150854 436920 150938
rect 436560 150618 436622 150854
rect 436858 150618 436920 150854
rect 409036 150586 409396 150618
rect 436560 150586 436920 150618
rect 535036 151174 535396 151206
rect 581514 151174 582134 186618
rect 535036 150938 535098 151174
rect 535334 150938 535396 151174
rect 535036 150854 535396 150938
rect 535036 150618 535098 150854
rect 535334 150618 535396 150854
rect 542000 150938 542032 151174
rect 542268 150938 542352 151174
rect 542588 150938 542620 151174
rect 542000 150854 542620 150938
rect 542000 150618 542032 150854
rect 542268 150618 542352 150854
rect 542588 150618 542620 150854
rect 571500 150938 571532 151174
rect 571768 150938 571852 151174
rect 572088 150938 572120 151174
rect 571500 150854 572120 150938
rect 571500 150618 571532 150854
rect 571768 150618 571852 150854
rect 572088 150618 572120 150854
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 535036 150586 535396 150618
rect 61280 147454 61640 147486
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect 9084 147218 9116 147454
rect 9352 147218 9436 147454
rect 9672 147218 9704 147454
rect 9084 147134 9704 147218
rect 9084 146898 9116 147134
rect 9352 146898 9436 147134
rect 9672 146898 9704 147134
rect 56620 147218 56652 147454
rect 56888 147218 56972 147454
rect 57208 147218 57240 147454
rect 56620 147134 57240 147218
rect 56620 146898 56652 147134
rect 56888 146898 56972 147134
rect 57208 146898 57240 147134
rect 61280 147218 61342 147454
rect 61578 147218 61640 147454
rect 61280 147134 61640 147218
rect 61280 146898 61342 147134
rect 61578 146898 61640 147134
rect -2006 111454 -1386 146898
rect 61280 146866 61640 146898
rect 158316 147454 158676 147486
rect 186280 147454 186640 147486
rect 158316 147218 158378 147454
rect 158614 147218 158676 147454
rect 158316 147134 158676 147218
rect 158316 146898 158378 147134
rect 158614 146898 158676 147134
rect 164620 147218 164652 147454
rect 164888 147218 164972 147454
rect 165208 147218 165240 147454
rect 164620 147134 165240 147218
rect 164620 146898 164652 147134
rect 164888 146898 164972 147134
rect 165208 146898 165240 147134
rect 186280 147218 186342 147454
rect 186578 147218 186640 147454
rect 186280 147134 186640 147218
rect 186280 146898 186342 147134
rect 186578 146898 186640 147134
rect 158316 146866 158676 146898
rect 186280 146866 186640 146898
rect 283316 147454 283676 147486
rect 311280 147454 311640 147486
rect 283316 147218 283378 147454
rect 283614 147218 283676 147454
rect 283316 147134 283676 147218
rect 283316 146898 283378 147134
rect 283614 146898 283676 147134
rect 308620 147218 308652 147454
rect 308888 147218 308972 147454
rect 309208 147218 309240 147454
rect 308620 147134 309240 147218
rect 308620 146898 308652 147134
rect 308888 146898 308972 147134
rect 309208 146898 309240 147134
rect 311280 147218 311342 147454
rect 311578 147218 311640 147454
rect 311280 147134 311640 147218
rect 311280 146898 311342 147134
rect 311578 146898 311640 147134
rect 283316 146866 283676 146898
rect 311280 146866 311640 146898
rect 408316 147454 408676 147486
rect 437280 147454 437640 147486
rect 408316 147218 408378 147454
rect 408614 147218 408676 147454
rect 408316 147134 408676 147218
rect 408316 146898 408378 147134
rect 408614 146898 408676 147134
rect 416620 147218 416652 147454
rect 416888 147218 416972 147454
rect 417208 147218 417240 147454
rect 416620 147134 417240 147218
rect 416620 146898 416652 147134
rect 416888 146898 416972 147134
rect 417208 146898 417240 147134
rect 437280 147218 437342 147454
rect 437578 147218 437640 147454
rect 437280 147134 437640 147218
rect 437280 146898 437342 147134
rect 437578 146898 437640 147134
rect 408316 146866 408676 146898
rect 437280 146866 437640 146898
rect 534316 147454 534676 147486
rect 534316 147218 534378 147454
rect 534614 147218 534676 147454
rect 534316 147134 534676 147218
rect 534316 146898 534378 147134
rect 534614 146898 534676 147134
rect 560620 147218 560652 147454
rect 560888 147218 560972 147454
rect 561208 147218 561240 147454
rect 560620 147134 561240 147218
rect 560620 146898 560652 147134
rect 560888 146898 560972 147134
rect 561208 146898 561240 147134
rect 570260 147218 570292 147454
rect 570528 147218 570612 147454
rect 570848 147218 570880 147454
rect 570260 147134 570880 147218
rect 570260 146898 570292 147134
rect 570528 146898 570612 147134
rect 570848 146898 570880 147134
rect 534316 146866 534676 146898
rect 61280 121244 61640 121300
rect 61280 121008 61342 121244
rect 61578 121008 61640 121244
rect 61280 120952 61640 121008
rect 62952 121244 63300 121300
rect 62952 121008 63008 121244
rect 63244 121008 63300 121244
rect 62952 120952 63300 121008
rect 281656 121244 282004 121300
rect 281656 121008 281712 121244
rect 281948 121008 282004 121244
rect 281656 120952 282004 121008
rect 283316 121244 283676 121300
rect 283316 121008 283378 121244
rect 283614 121008 283676 121244
rect 283316 120952 283676 121008
rect 311280 121244 311640 121300
rect 311280 121008 311342 121244
rect 311578 121008 311640 121244
rect 311280 120952 311640 121008
rect 312952 121244 313300 121300
rect 312952 121008 313008 121244
rect 313244 121008 313300 121244
rect 312952 120952 313300 121008
rect 532656 121244 533004 121300
rect 532656 121008 532712 121244
rect 532948 121008 533004 121244
rect 532656 120952 533004 121008
rect 534316 121244 534676 121300
rect 534316 121008 534378 121244
rect 534614 121008 534676 121244
rect 534316 120952 534676 121008
rect 157336 120564 157684 120620
rect 157336 120328 157392 120564
rect 157628 120328 157684 120564
rect 157336 120272 157684 120328
rect 159036 120564 159396 120620
rect 159036 120328 159098 120564
rect 159334 120328 159396 120564
rect 159036 120272 159396 120328
rect 185560 120564 185920 120620
rect 185560 120328 185622 120564
rect 185858 120328 185920 120564
rect 185560 120272 185920 120328
rect 187272 120564 187620 120620
rect 187272 120328 187328 120564
rect 187564 120328 187620 120564
rect 187272 120272 187620 120328
rect 407336 120564 407684 120620
rect 407336 120328 407392 120564
rect 407628 120328 407684 120564
rect 407336 120272 407684 120328
rect 409036 120564 409396 120620
rect 409036 120328 409098 120564
rect 409334 120328 409396 120564
rect 409036 120272 409396 120328
rect 436560 120564 436920 120620
rect 436560 120328 436622 120564
rect 436858 120328 436920 120564
rect 436560 120272 436920 120328
rect 438272 120564 438620 120620
rect 438272 120328 438328 120564
rect 438564 120328 438620 120564
rect 438272 120272 438620 120328
rect 581514 115174 582134 150618
rect 7844 114938 7876 115174
rect 8112 114938 8196 115174
rect 8432 114938 8464 115174
rect 7844 114854 8464 114938
rect 7844 114618 7876 114854
rect 8112 114618 8196 114854
rect 8432 114618 8464 114854
rect 38000 114938 38032 115174
rect 38268 114938 38352 115174
rect 38588 114938 38620 115174
rect 38000 114854 38620 114938
rect 38000 114618 38032 114854
rect 38268 114618 38352 114854
rect 38588 114618 38620 114854
rect 74000 114938 74032 115174
rect 74268 114938 74352 115174
rect 74588 114938 74620 115174
rect 74000 114854 74620 114938
rect 74000 114618 74032 114854
rect 74268 114618 74352 114854
rect 74588 114618 74620 114854
rect 110000 114938 110032 115174
rect 110268 114938 110352 115174
rect 110588 114938 110620 115174
rect 110000 114854 110620 114938
rect 110000 114618 110032 114854
rect 110268 114618 110352 114854
rect 110588 114618 110620 114854
rect 146000 114938 146032 115174
rect 146268 114938 146352 115174
rect 146588 114938 146620 115174
rect 146000 114854 146620 114938
rect 146000 114618 146032 114854
rect 146268 114618 146352 114854
rect 146588 114618 146620 114854
rect 182000 114938 182032 115174
rect 182268 114938 182352 115174
rect 182588 114938 182620 115174
rect 182000 114854 182620 114938
rect 182000 114618 182032 114854
rect 182268 114618 182352 114854
rect 182588 114618 182620 114854
rect 218000 114938 218032 115174
rect 218268 114938 218352 115174
rect 218588 114938 218620 115174
rect 218000 114854 218620 114938
rect 218000 114618 218032 114854
rect 218268 114618 218352 114854
rect 218588 114618 218620 114854
rect 254000 114938 254032 115174
rect 254268 114938 254352 115174
rect 254588 114938 254620 115174
rect 254000 114854 254620 114938
rect 254000 114618 254032 114854
rect 254268 114618 254352 114854
rect 254588 114618 254620 114854
rect 290000 114938 290032 115174
rect 290268 114938 290352 115174
rect 290588 114938 290620 115174
rect 290000 114854 290620 114938
rect 290000 114618 290032 114854
rect 290268 114618 290352 114854
rect 290588 114618 290620 114854
rect 326000 114938 326032 115174
rect 326268 114938 326352 115174
rect 326588 114938 326620 115174
rect 326000 114854 326620 114938
rect 326000 114618 326032 114854
rect 326268 114618 326352 114854
rect 326588 114618 326620 114854
rect 362000 114938 362032 115174
rect 362268 114938 362352 115174
rect 362588 114938 362620 115174
rect 362000 114854 362620 114938
rect 362000 114618 362032 114854
rect 362268 114618 362352 114854
rect 362588 114618 362620 114854
rect 398000 114938 398032 115174
rect 398268 114938 398352 115174
rect 398588 114938 398620 115174
rect 398000 114854 398620 114938
rect 398000 114618 398032 114854
rect 398268 114618 398352 114854
rect 398588 114618 398620 114854
rect 434000 114938 434032 115174
rect 434268 114938 434352 115174
rect 434588 114938 434620 115174
rect 434000 114854 434620 114938
rect 434000 114618 434032 114854
rect 434268 114618 434352 114854
rect 434588 114618 434620 114854
rect 470000 114938 470032 115174
rect 470268 114938 470352 115174
rect 470588 114938 470620 115174
rect 470000 114854 470620 114938
rect 470000 114618 470032 114854
rect 470268 114618 470352 114854
rect 470588 114618 470620 114854
rect 506000 114938 506032 115174
rect 506268 114938 506352 115174
rect 506588 114938 506620 115174
rect 506000 114854 506620 114938
rect 506000 114618 506032 114854
rect 506268 114618 506352 114854
rect 506588 114618 506620 114854
rect 542000 114938 542032 115174
rect 542268 114938 542352 115174
rect 542588 114938 542620 115174
rect 542000 114854 542620 114938
rect 542000 114618 542032 114854
rect 542268 114618 542352 114854
rect 542588 114618 542620 114854
rect 571500 114938 571532 115174
rect 571768 114938 571852 115174
rect 572088 114938 572120 115174
rect 571500 114854 572120 114938
rect 571500 114618 571532 114854
rect 571768 114618 571852 114854
rect 572088 114618 572120 114854
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect 9084 111218 9116 111454
rect 9352 111218 9436 111454
rect 9672 111218 9704 111454
rect 9084 111134 9704 111218
rect 9084 110898 9116 111134
rect 9352 110898 9436 111134
rect 9672 110898 9704 111134
rect 56620 111218 56652 111454
rect 56888 111218 56972 111454
rect 57208 111218 57240 111454
rect 56620 111134 57240 111218
rect 56620 110898 56652 111134
rect 56888 110898 56972 111134
rect 57208 110898 57240 111134
rect 92620 111218 92652 111454
rect 92888 111218 92972 111454
rect 93208 111218 93240 111454
rect 92620 111134 93240 111218
rect 92620 110898 92652 111134
rect 92888 110898 92972 111134
rect 93208 110898 93240 111134
rect 128620 111218 128652 111454
rect 128888 111218 128972 111454
rect 129208 111218 129240 111454
rect 128620 111134 129240 111218
rect 128620 110898 128652 111134
rect 128888 110898 128972 111134
rect 129208 110898 129240 111134
rect 164620 111218 164652 111454
rect 164888 111218 164972 111454
rect 165208 111218 165240 111454
rect 164620 111134 165240 111218
rect 164620 110898 164652 111134
rect 164888 110898 164972 111134
rect 165208 110898 165240 111134
rect 200620 111218 200652 111454
rect 200888 111218 200972 111454
rect 201208 111218 201240 111454
rect 200620 111134 201240 111218
rect 200620 110898 200652 111134
rect 200888 110898 200972 111134
rect 201208 110898 201240 111134
rect 236620 111218 236652 111454
rect 236888 111218 236972 111454
rect 237208 111218 237240 111454
rect 236620 111134 237240 111218
rect 236620 110898 236652 111134
rect 236888 110898 236972 111134
rect 237208 110898 237240 111134
rect 272620 111218 272652 111454
rect 272888 111218 272972 111454
rect 273208 111218 273240 111454
rect 272620 111134 273240 111218
rect 272620 110898 272652 111134
rect 272888 110898 272972 111134
rect 273208 110898 273240 111134
rect 308620 111218 308652 111454
rect 308888 111218 308972 111454
rect 309208 111218 309240 111454
rect 308620 111134 309240 111218
rect 308620 110898 308652 111134
rect 308888 110898 308972 111134
rect 309208 110898 309240 111134
rect 344620 111218 344652 111454
rect 344888 111218 344972 111454
rect 345208 111218 345240 111454
rect 344620 111134 345240 111218
rect 344620 110898 344652 111134
rect 344888 110898 344972 111134
rect 345208 110898 345240 111134
rect 380620 111218 380652 111454
rect 380888 111218 380972 111454
rect 381208 111218 381240 111454
rect 380620 111134 381240 111218
rect 380620 110898 380652 111134
rect 380888 110898 380972 111134
rect 381208 110898 381240 111134
rect 416620 111218 416652 111454
rect 416888 111218 416972 111454
rect 417208 111218 417240 111454
rect 416620 111134 417240 111218
rect 416620 110898 416652 111134
rect 416888 110898 416972 111134
rect 417208 110898 417240 111134
rect 452620 111218 452652 111454
rect 452888 111218 452972 111454
rect 453208 111218 453240 111454
rect 452620 111134 453240 111218
rect 452620 110898 452652 111134
rect 452888 110898 452972 111134
rect 453208 110898 453240 111134
rect 488620 111218 488652 111454
rect 488888 111218 488972 111454
rect 489208 111218 489240 111454
rect 488620 111134 489240 111218
rect 488620 110898 488652 111134
rect 488888 110898 488972 111134
rect 489208 110898 489240 111134
rect 524620 111218 524652 111454
rect 524888 111218 524972 111454
rect 525208 111218 525240 111454
rect 524620 111134 525240 111218
rect 524620 110898 524652 111134
rect 524888 110898 524972 111134
rect 525208 110898 525240 111134
rect 560620 111218 560652 111454
rect 560888 111218 560972 111454
rect 561208 111218 561240 111454
rect 560620 111134 561240 111218
rect 560620 110898 560652 111134
rect 560888 110898 560972 111134
rect 561208 110898 561240 111134
rect 570260 111218 570292 111454
rect 570528 111218 570612 111454
rect 570848 111218 570880 111454
rect 570260 111134 570880 111218
rect 570260 110898 570292 111134
rect 570528 110898 570612 111134
rect 570848 110898 570880 111134
rect -2006 75454 -1386 110898
rect 60560 79174 60920 79206
rect 7844 78938 7876 79174
rect 8112 78938 8196 79174
rect 8432 78938 8464 79174
rect 7844 78854 8464 78938
rect 7844 78618 7876 78854
rect 8112 78618 8196 78854
rect 8432 78618 8464 78854
rect 38000 78938 38032 79174
rect 38268 78938 38352 79174
rect 38588 78938 38620 79174
rect 38000 78854 38620 78938
rect 38000 78618 38032 78854
rect 38268 78618 38352 78854
rect 38588 78618 38620 78854
rect 60560 78938 60622 79174
rect 60858 78938 60920 79174
rect 60560 78854 60920 78938
rect 60560 78618 60622 78854
rect 60858 78618 60920 78854
rect 60560 78586 60920 78618
rect 159036 79174 159396 79206
rect 185560 79174 185920 79206
rect 159036 78938 159098 79174
rect 159334 78938 159396 79174
rect 159036 78854 159396 78938
rect 159036 78618 159098 78854
rect 159334 78618 159396 78854
rect 182000 78938 182032 79174
rect 182268 78938 182352 79174
rect 182588 78938 182620 79174
rect 182000 78854 182620 78938
rect 182000 78618 182032 78854
rect 182268 78618 182352 78854
rect 182588 78618 182620 78854
rect 185560 78938 185622 79174
rect 185858 78938 185920 79174
rect 185560 78854 185920 78938
rect 185560 78618 185622 78854
rect 185858 78618 185920 78854
rect 159036 78586 159396 78618
rect 185560 78586 185920 78618
rect 284036 79174 284396 79206
rect 310560 79174 310920 79206
rect 284036 78938 284098 79174
rect 284334 78938 284396 79174
rect 284036 78854 284396 78938
rect 284036 78618 284098 78854
rect 284334 78618 284396 78854
rect 290000 78938 290032 79174
rect 290268 78938 290352 79174
rect 290588 78938 290620 79174
rect 290000 78854 290620 78938
rect 290000 78618 290032 78854
rect 290268 78618 290352 78854
rect 290588 78618 290620 78854
rect 310560 78938 310622 79174
rect 310858 78938 310920 79174
rect 310560 78854 310920 78938
rect 310560 78618 310622 78854
rect 310858 78618 310920 78854
rect 284036 78586 284396 78618
rect 310560 78586 310920 78618
rect 409036 79174 409396 79206
rect 436560 79174 436920 79206
rect 409036 78938 409098 79174
rect 409334 78938 409396 79174
rect 409036 78854 409396 78938
rect 409036 78618 409098 78854
rect 409334 78618 409396 78854
rect 434000 78938 434032 79174
rect 434268 78938 434352 79174
rect 434588 78938 434620 79174
rect 434000 78854 434620 78938
rect 434000 78618 434032 78854
rect 434268 78618 434352 78854
rect 434588 78618 434620 78854
rect 436560 78938 436622 79174
rect 436858 78938 436920 79174
rect 436560 78854 436920 78938
rect 436560 78618 436622 78854
rect 436858 78618 436920 78854
rect 409036 78586 409396 78618
rect 436560 78586 436920 78618
rect 535036 79174 535396 79206
rect 581514 79174 582134 114618
rect 535036 78938 535098 79174
rect 535334 78938 535396 79174
rect 535036 78854 535396 78938
rect 535036 78618 535098 78854
rect 535334 78618 535396 78854
rect 542000 78938 542032 79174
rect 542268 78938 542352 79174
rect 542588 78938 542620 79174
rect 542000 78854 542620 78938
rect 542000 78618 542032 78854
rect 542268 78618 542352 78854
rect 542588 78618 542620 78854
rect 571500 78938 571532 79174
rect 571768 78938 571852 79174
rect 572088 78938 572120 79174
rect 571500 78854 572120 78938
rect 571500 78618 571532 78854
rect 571768 78618 571852 78854
rect 572088 78618 572120 78854
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 535036 78586 535396 78618
rect 61280 75454 61640 75486
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect 9084 75218 9116 75454
rect 9352 75218 9436 75454
rect 9672 75218 9704 75454
rect 9084 75134 9704 75218
rect 9084 74898 9116 75134
rect 9352 74898 9436 75134
rect 9672 74898 9704 75134
rect 56620 75218 56652 75454
rect 56888 75218 56972 75454
rect 57208 75218 57240 75454
rect 56620 75134 57240 75218
rect 56620 74898 56652 75134
rect 56888 74898 56972 75134
rect 57208 74898 57240 75134
rect 61280 75218 61342 75454
rect 61578 75218 61640 75454
rect 61280 75134 61640 75218
rect 61280 74898 61342 75134
rect 61578 74898 61640 75134
rect -2006 39454 -1386 74898
rect 61280 74866 61640 74898
rect 158316 75454 158676 75486
rect 186280 75454 186640 75486
rect 158316 75218 158378 75454
rect 158614 75218 158676 75454
rect 158316 75134 158676 75218
rect 158316 74898 158378 75134
rect 158614 74898 158676 75134
rect 164620 75218 164652 75454
rect 164888 75218 164972 75454
rect 165208 75218 165240 75454
rect 164620 75134 165240 75218
rect 164620 74898 164652 75134
rect 164888 74898 164972 75134
rect 165208 74898 165240 75134
rect 186280 75218 186342 75454
rect 186578 75218 186640 75454
rect 186280 75134 186640 75218
rect 186280 74898 186342 75134
rect 186578 74898 186640 75134
rect 158316 74866 158676 74898
rect 186280 74866 186640 74898
rect 283316 75454 283676 75486
rect 311280 75454 311640 75486
rect 283316 75218 283378 75454
rect 283614 75218 283676 75454
rect 283316 75134 283676 75218
rect 283316 74898 283378 75134
rect 283614 74898 283676 75134
rect 308620 75218 308652 75454
rect 308888 75218 308972 75454
rect 309208 75218 309240 75454
rect 308620 75134 309240 75218
rect 308620 74898 308652 75134
rect 308888 74898 308972 75134
rect 309208 74898 309240 75134
rect 311280 75218 311342 75454
rect 311578 75218 311640 75454
rect 311280 75134 311640 75218
rect 311280 74898 311342 75134
rect 311578 74898 311640 75134
rect 283316 74866 283676 74898
rect 311280 74866 311640 74898
rect 408316 75454 408676 75486
rect 437280 75454 437640 75486
rect 408316 75218 408378 75454
rect 408614 75218 408676 75454
rect 408316 75134 408676 75218
rect 408316 74898 408378 75134
rect 408614 74898 408676 75134
rect 416620 75218 416652 75454
rect 416888 75218 416972 75454
rect 417208 75218 417240 75454
rect 416620 75134 417240 75218
rect 416620 74898 416652 75134
rect 416888 74898 416972 75134
rect 417208 74898 417240 75134
rect 437280 75218 437342 75454
rect 437578 75218 437640 75454
rect 437280 75134 437640 75218
rect 437280 74898 437342 75134
rect 437578 74898 437640 75134
rect 408316 74866 408676 74898
rect 437280 74866 437640 74898
rect 534316 75454 534676 75486
rect 534316 75218 534378 75454
rect 534614 75218 534676 75454
rect 534316 75134 534676 75218
rect 534316 74898 534378 75134
rect 534614 74898 534676 75134
rect 560620 75218 560652 75454
rect 560888 75218 560972 75454
rect 561208 75218 561240 75454
rect 560620 75134 561240 75218
rect 560620 74898 560652 75134
rect 560888 74898 560972 75134
rect 561208 74898 561240 75134
rect 570260 75218 570292 75454
rect 570528 75218 570612 75454
rect 570848 75218 570880 75454
rect 570260 75134 570880 75218
rect 570260 74898 570292 75134
rect 570528 74898 570612 75134
rect 570848 74898 570880 75134
rect 534316 74866 534676 74898
rect 60560 43174 60920 43206
rect 7844 42938 7876 43174
rect 8112 42938 8196 43174
rect 8432 42938 8464 43174
rect 7844 42854 8464 42938
rect 7844 42618 7876 42854
rect 8112 42618 8196 42854
rect 8432 42618 8464 42854
rect 38000 42938 38032 43174
rect 38268 42938 38352 43174
rect 38588 42938 38620 43174
rect 38000 42854 38620 42938
rect 38000 42618 38032 42854
rect 38268 42618 38352 42854
rect 38588 42618 38620 42854
rect 60560 42938 60622 43174
rect 60858 42938 60920 43174
rect 60560 42854 60920 42938
rect 60560 42618 60622 42854
rect 60858 42618 60920 42854
rect 60560 42586 60920 42618
rect 159036 43174 159396 43206
rect 185560 43174 185920 43206
rect 159036 42938 159098 43174
rect 159334 42938 159396 43174
rect 159036 42854 159396 42938
rect 159036 42618 159098 42854
rect 159334 42618 159396 42854
rect 182000 42938 182032 43174
rect 182268 42938 182352 43174
rect 182588 42938 182620 43174
rect 182000 42854 182620 42938
rect 182000 42618 182032 42854
rect 182268 42618 182352 42854
rect 182588 42618 182620 42854
rect 185560 42938 185622 43174
rect 185858 42938 185920 43174
rect 185560 42854 185920 42938
rect 185560 42618 185622 42854
rect 185858 42618 185920 42854
rect 159036 42586 159396 42618
rect 185560 42586 185920 42618
rect 284036 43174 284396 43206
rect 310560 43174 310920 43206
rect 284036 42938 284098 43174
rect 284334 42938 284396 43174
rect 284036 42854 284396 42938
rect 284036 42618 284098 42854
rect 284334 42618 284396 42854
rect 290000 42938 290032 43174
rect 290268 42938 290352 43174
rect 290588 42938 290620 43174
rect 290000 42854 290620 42938
rect 290000 42618 290032 42854
rect 290268 42618 290352 42854
rect 290588 42618 290620 42854
rect 310560 42938 310622 43174
rect 310858 42938 310920 43174
rect 310560 42854 310920 42938
rect 310560 42618 310622 42854
rect 310858 42618 310920 42854
rect 284036 42586 284396 42618
rect 310560 42586 310920 42618
rect 409036 43174 409396 43206
rect 436560 43174 436920 43206
rect 409036 42938 409098 43174
rect 409334 42938 409396 43174
rect 409036 42854 409396 42938
rect 409036 42618 409098 42854
rect 409334 42618 409396 42854
rect 434000 42938 434032 43174
rect 434268 42938 434352 43174
rect 434588 42938 434620 43174
rect 434000 42854 434620 42938
rect 434000 42618 434032 42854
rect 434268 42618 434352 42854
rect 434588 42618 434620 42854
rect 436560 42938 436622 43174
rect 436858 42938 436920 43174
rect 436560 42854 436920 42938
rect 436560 42618 436622 42854
rect 436858 42618 436920 42854
rect 409036 42586 409396 42618
rect 436560 42586 436920 42618
rect 535036 43174 535396 43206
rect 581514 43174 582134 78618
rect 535036 42938 535098 43174
rect 535334 42938 535396 43174
rect 535036 42854 535396 42938
rect 535036 42618 535098 42854
rect 535334 42618 535396 42854
rect 542000 42938 542032 43174
rect 542268 42938 542352 43174
rect 542588 42938 542620 43174
rect 542000 42854 542620 42938
rect 542000 42618 542032 42854
rect 542268 42618 542352 42854
rect 542588 42618 542620 42854
rect 571500 42938 571532 43174
rect 571768 42938 571852 43174
rect 572088 42938 572120 43174
rect 571500 42854 572120 42938
rect 571500 42618 571532 42854
rect 571768 42618 571852 42854
rect 572088 42618 572120 42854
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 535036 42586 535396 42618
rect 61280 39454 61640 39486
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect 9084 39218 9116 39454
rect 9352 39218 9436 39454
rect 9672 39218 9704 39454
rect 9084 39134 9704 39218
rect 9084 38898 9116 39134
rect 9352 38898 9436 39134
rect 9672 38898 9704 39134
rect 56620 39218 56652 39454
rect 56888 39218 56972 39454
rect 57208 39218 57240 39454
rect 56620 39134 57240 39218
rect 56620 38898 56652 39134
rect 56888 38898 56972 39134
rect 57208 38898 57240 39134
rect 61280 39218 61342 39454
rect 61578 39218 61640 39454
rect 61280 39134 61640 39218
rect 61280 38898 61342 39134
rect 61578 38898 61640 39134
rect -2006 3454 -1386 38898
rect 61280 38866 61640 38898
rect 158316 39454 158676 39486
rect 186280 39454 186640 39486
rect 158316 39218 158378 39454
rect 158614 39218 158676 39454
rect 158316 39134 158676 39218
rect 158316 38898 158378 39134
rect 158614 38898 158676 39134
rect 164620 39218 164652 39454
rect 164888 39218 164972 39454
rect 165208 39218 165240 39454
rect 164620 39134 165240 39218
rect 164620 38898 164652 39134
rect 164888 38898 164972 39134
rect 165208 38898 165240 39134
rect 186280 39218 186342 39454
rect 186578 39218 186640 39454
rect 186280 39134 186640 39218
rect 186280 38898 186342 39134
rect 186578 38898 186640 39134
rect 158316 38866 158676 38898
rect 186280 38866 186640 38898
rect 283316 39454 283676 39486
rect 311280 39454 311640 39486
rect 283316 39218 283378 39454
rect 283614 39218 283676 39454
rect 283316 39134 283676 39218
rect 283316 38898 283378 39134
rect 283614 38898 283676 39134
rect 308620 39218 308652 39454
rect 308888 39218 308972 39454
rect 309208 39218 309240 39454
rect 308620 39134 309240 39218
rect 308620 38898 308652 39134
rect 308888 38898 308972 39134
rect 309208 38898 309240 39134
rect 311280 39218 311342 39454
rect 311578 39218 311640 39454
rect 311280 39134 311640 39218
rect 311280 38898 311342 39134
rect 311578 38898 311640 39134
rect 283316 38866 283676 38898
rect 311280 38866 311640 38898
rect 408316 39454 408676 39486
rect 437280 39454 437640 39486
rect 408316 39218 408378 39454
rect 408614 39218 408676 39454
rect 408316 39134 408676 39218
rect 408316 38898 408378 39134
rect 408614 38898 408676 39134
rect 416620 39218 416652 39454
rect 416888 39218 416972 39454
rect 417208 39218 417240 39454
rect 416620 39134 417240 39218
rect 416620 38898 416652 39134
rect 416888 38898 416972 39134
rect 417208 38898 417240 39134
rect 437280 39218 437342 39454
rect 437578 39218 437640 39454
rect 437280 39134 437640 39218
rect 437280 38898 437342 39134
rect 437578 38898 437640 39134
rect 408316 38866 408676 38898
rect 437280 38866 437640 38898
rect 534316 39454 534676 39486
rect 534316 39218 534378 39454
rect 534614 39218 534676 39454
rect 534316 39134 534676 39218
rect 534316 38898 534378 39134
rect 534614 38898 534676 39134
rect 560620 39218 560652 39454
rect 560888 39218 560972 39454
rect 561208 39218 561240 39454
rect 560620 39134 561240 39218
rect 560620 38898 560652 39134
rect 560888 38898 560972 39134
rect 561208 38898 561240 39134
rect 570260 39218 570292 39454
rect 570528 39218 570612 39454
rect 570848 39218 570880 39454
rect 570260 39134 570880 39218
rect 570260 38898 570292 39134
rect 570528 38898 570612 39134
rect 570848 38898 570880 39134
rect 534316 38866 534676 38898
rect 61280 21244 61640 21300
rect 61280 21008 61342 21244
rect 61578 21008 61640 21244
rect 61280 20952 61640 21008
rect 62952 21244 63300 21300
rect 62952 21008 63008 21244
rect 63244 21008 63300 21244
rect 62952 20952 63300 21008
rect 187952 21244 188300 21300
rect 187952 21008 188008 21244
rect 188244 21008 188300 21244
rect 187952 20952 188300 21008
rect 311280 21244 311640 21300
rect 311280 21008 311342 21244
rect 311578 21008 311640 21244
rect 311280 20952 311640 21008
rect 312952 21244 313300 21300
rect 312952 21008 313008 21244
rect 313244 21008 313300 21244
rect 312952 20952 313300 21008
rect 438952 21244 439300 21300
rect 438952 21008 439008 21244
rect 439244 21008 439300 21244
rect 438952 20952 439300 21008
rect 62272 20564 62620 20620
rect 62272 20328 62328 20564
rect 62564 20328 62620 20564
rect 62272 20272 62620 20328
rect 185560 20564 185920 20620
rect 185560 20328 185622 20564
rect 185858 20328 185920 20564
rect 185560 20272 185920 20328
rect 187272 20564 187620 20620
rect 187272 20328 187328 20564
rect 187564 20328 187620 20564
rect 187272 20272 187620 20328
rect 312272 20564 312620 20620
rect 312272 20328 312328 20564
rect 312564 20328 312620 20564
rect 312272 20272 312620 20328
rect 436560 20564 436920 20620
rect 436560 20328 436622 20564
rect 436858 20328 436920 20564
rect 436560 20272 436920 20328
rect 438272 20564 438620 20620
rect 438272 20328 438328 20564
rect 438564 20328 438620 20564
rect 438272 20272 438620 20328
rect 62272 19834 62620 19858
rect 62272 19598 62328 19834
rect 62564 19598 62620 19834
rect 312272 19834 312620 19858
rect 62272 19574 62620 19598
rect 187952 19578 188300 19640
rect 187952 19342 188008 19578
rect 188244 19342 188300 19578
rect 312272 19598 312328 19834
rect 312564 19598 312620 19834
rect 312272 19574 312620 19598
rect 438952 19578 439300 19640
rect 187952 19280 188300 19342
rect 438952 19342 439008 19578
rect 439244 19342 439300 19578
rect 438952 19280 439300 19342
rect 9084 9444 9116 9680
rect 9352 9444 9436 9680
rect 9672 9444 9704 9680
rect 9084 9360 9704 9444
rect 9084 9124 9116 9360
rect 9352 9124 9436 9360
rect 9672 9124 9704 9360
rect 56620 9444 56652 9680
rect 56888 9444 56972 9680
rect 57208 9444 57240 9680
rect 56620 9360 57240 9444
rect 56620 9124 56652 9360
rect 56888 9124 56972 9360
rect 57208 9124 57240 9360
rect 92620 9444 92652 9680
rect 92888 9444 92972 9680
rect 93208 9444 93240 9680
rect 92620 9360 93240 9444
rect 92620 9124 92652 9360
rect 92888 9124 92972 9360
rect 93208 9124 93240 9360
rect 128620 9444 128652 9680
rect 128888 9444 128972 9680
rect 129208 9444 129240 9680
rect 128620 9360 129240 9444
rect 128620 9124 128652 9360
rect 128888 9124 128972 9360
rect 129208 9124 129240 9360
rect 164620 9444 164652 9680
rect 164888 9444 164972 9680
rect 165208 9444 165240 9680
rect 164620 9360 165240 9444
rect 164620 9124 164652 9360
rect 164888 9124 164972 9360
rect 165208 9124 165240 9360
rect 200620 9444 200652 9680
rect 200888 9444 200972 9680
rect 201208 9444 201240 9680
rect 200620 9360 201240 9444
rect 200620 9124 200652 9360
rect 200888 9124 200972 9360
rect 201208 9124 201240 9360
rect 236620 9444 236652 9680
rect 236888 9444 236972 9680
rect 237208 9444 237240 9680
rect 236620 9360 237240 9444
rect 236620 9124 236652 9360
rect 236888 9124 236972 9360
rect 237208 9124 237240 9360
rect 272620 9444 272652 9680
rect 272888 9444 272972 9680
rect 273208 9444 273240 9680
rect 272620 9360 273240 9444
rect 272620 9124 272652 9360
rect 272888 9124 272972 9360
rect 273208 9124 273240 9360
rect 308620 9444 308652 9680
rect 308888 9444 308972 9680
rect 309208 9444 309240 9680
rect 308620 9360 309240 9444
rect 308620 9124 308652 9360
rect 308888 9124 308972 9360
rect 309208 9124 309240 9360
rect 344620 9444 344652 9680
rect 344888 9444 344972 9680
rect 345208 9444 345240 9680
rect 344620 9360 345240 9444
rect 344620 9124 344652 9360
rect 344888 9124 344972 9360
rect 345208 9124 345240 9360
rect 380620 9444 380652 9680
rect 380888 9444 380972 9680
rect 381208 9444 381240 9680
rect 380620 9360 381240 9444
rect 380620 9124 380652 9360
rect 380888 9124 380972 9360
rect 381208 9124 381240 9360
rect 416620 9444 416652 9680
rect 416888 9444 416972 9680
rect 417208 9444 417240 9680
rect 416620 9360 417240 9444
rect 416620 9124 416652 9360
rect 416888 9124 416972 9360
rect 417208 9124 417240 9360
rect 452620 9444 452652 9680
rect 452888 9444 452972 9680
rect 453208 9444 453240 9680
rect 452620 9360 453240 9444
rect 452620 9124 452652 9360
rect 452888 9124 452972 9360
rect 453208 9124 453240 9360
rect 488620 9444 488652 9680
rect 488888 9444 488972 9680
rect 489208 9444 489240 9680
rect 488620 9360 489240 9444
rect 488620 9124 488652 9360
rect 488888 9124 488972 9360
rect 489208 9124 489240 9360
rect 524620 9444 524652 9680
rect 524888 9444 524972 9680
rect 525208 9444 525240 9680
rect 524620 9360 525240 9444
rect 524620 9124 524652 9360
rect 524888 9124 524972 9360
rect 525208 9124 525240 9360
rect 560620 9444 560652 9680
rect 560888 9444 560972 9680
rect 561208 9444 561240 9680
rect 560620 9360 561240 9444
rect 560620 9124 560652 9360
rect 560888 9124 560972 9360
rect 561208 9124 561240 9360
rect 570260 9444 570292 9680
rect 570528 9444 570612 9680
rect 570848 9444 570880 9680
rect 570260 9360 570880 9444
rect 570260 9124 570292 9360
rect 570528 9124 570612 9360
rect 570848 9124 570880 9360
rect 7844 8204 7876 8440
rect 8112 8204 8196 8440
rect 8432 8204 8464 8440
rect 7844 8120 8464 8204
rect 7844 7884 7876 8120
rect 8112 7884 8196 8120
rect 8432 7884 8464 8120
rect 38000 8204 38032 8440
rect 38268 8204 38352 8440
rect 38588 8204 38620 8440
rect 38000 8120 38620 8204
rect 38000 7884 38032 8120
rect 38268 7884 38352 8120
rect 38588 7884 38620 8120
rect 74000 8204 74032 8440
rect 74268 8204 74352 8440
rect 74588 8204 74620 8440
rect 74000 8120 74620 8204
rect 74000 7884 74032 8120
rect 74268 7884 74352 8120
rect 74588 7884 74620 8120
rect 110000 8204 110032 8440
rect 110268 8204 110352 8440
rect 110588 8204 110620 8440
rect 110000 8120 110620 8204
rect 110000 7884 110032 8120
rect 110268 7884 110352 8120
rect 110588 7884 110620 8120
rect 146000 8204 146032 8440
rect 146268 8204 146352 8440
rect 146588 8204 146620 8440
rect 146000 8120 146620 8204
rect 146000 7884 146032 8120
rect 146268 7884 146352 8120
rect 146588 7884 146620 8120
rect 182000 8204 182032 8440
rect 182268 8204 182352 8440
rect 182588 8204 182620 8440
rect 182000 8120 182620 8204
rect 182000 7884 182032 8120
rect 182268 7884 182352 8120
rect 182588 7884 182620 8120
rect 218000 8204 218032 8440
rect 218268 8204 218352 8440
rect 218588 8204 218620 8440
rect 218000 8120 218620 8204
rect 218000 7884 218032 8120
rect 218268 7884 218352 8120
rect 218588 7884 218620 8120
rect 254000 8204 254032 8440
rect 254268 8204 254352 8440
rect 254588 8204 254620 8440
rect 254000 8120 254620 8204
rect 254000 7884 254032 8120
rect 254268 7884 254352 8120
rect 254588 7884 254620 8120
rect 290000 8204 290032 8440
rect 290268 8204 290352 8440
rect 290588 8204 290620 8440
rect 290000 8120 290620 8204
rect 290000 7884 290032 8120
rect 290268 7884 290352 8120
rect 290588 7884 290620 8120
rect 326000 8204 326032 8440
rect 326268 8204 326352 8440
rect 326588 8204 326620 8440
rect 326000 8120 326620 8204
rect 326000 7884 326032 8120
rect 326268 7884 326352 8120
rect 326588 7884 326620 8120
rect 362000 8204 362032 8440
rect 362268 8204 362352 8440
rect 362588 8204 362620 8440
rect 362000 8120 362620 8204
rect 362000 7884 362032 8120
rect 362268 7884 362352 8120
rect 362588 7884 362620 8120
rect 398000 8204 398032 8440
rect 398268 8204 398352 8440
rect 398588 8204 398620 8440
rect 398000 8120 398620 8204
rect 398000 7884 398032 8120
rect 398268 7884 398352 8120
rect 398588 7884 398620 8120
rect 434000 8204 434032 8440
rect 434268 8204 434352 8440
rect 434588 8204 434620 8440
rect 434000 8120 434620 8204
rect 434000 7884 434032 8120
rect 434268 7884 434352 8120
rect 434588 7884 434620 8120
rect 470000 8204 470032 8440
rect 470268 8204 470352 8440
rect 470588 8204 470620 8440
rect 470000 8120 470620 8204
rect 470000 7884 470032 8120
rect 470268 7884 470352 8120
rect 470588 7884 470620 8120
rect 506000 8204 506032 8440
rect 506268 8204 506352 8440
rect 506588 8204 506620 8440
rect 506000 8120 506620 8204
rect 506000 7884 506032 8120
rect 506268 7884 506352 8120
rect 506588 7884 506620 8120
rect 542000 8204 542032 8440
rect 542268 8204 542352 8440
rect 542588 8204 542620 8440
rect 542000 8120 542620 8204
rect 542000 7884 542032 8120
rect 542268 7884 542352 8120
rect 542588 7884 542620 8120
rect 571500 8204 571532 8440
rect 571768 8204 571852 8440
rect 572088 8204 572120 8440
rect 571500 8120 572120 8204
rect 571500 7884 571532 8120
rect 571768 7884 571852 8120
rect 572088 7884 572120 8120
rect 581514 7174 582134 42618
rect 7844 6938 7876 7174
rect 8112 6938 8196 7174
rect 8432 6938 8464 7174
rect 7844 6854 8464 6938
rect 7844 6618 7876 6854
rect 8112 6618 8196 6854
rect 8432 6618 8464 6854
rect 571500 6938 571532 7174
rect 571768 6938 571852 7174
rect 572088 6938 572120 7174
rect 571500 6854 572120 6938
rect 571500 6618 571532 6854
rect 571768 6618 571852 6854
rect 572088 6618 572120 6854
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect -5116 -3692 -5084 -3456
rect -4848 -3692 -4764 -3456
rect -4528 -3692 -4496 -3456
rect -5116 -3776 -4496 -3692
rect -5116 -4012 -5084 -3776
rect -4848 -4012 -4764 -3776
rect -4528 -4012 -4496 -3776
rect -5116 -4044 -4496 -4012
rect 581514 -3456 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 588420 691174 589040 707392
rect 588420 690938 588452 691174
rect 588688 690938 588772 691174
rect 589008 690938 589040 691174
rect 588420 690854 589040 690938
rect 588420 690618 588452 690854
rect 588688 690618 588772 690854
rect 589008 690618 589040 690854
rect 588420 655174 589040 690618
rect 588420 654938 588452 655174
rect 588688 654938 588772 655174
rect 589008 654938 589040 655174
rect 588420 654854 589040 654938
rect 588420 654618 588452 654854
rect 588688 654618 588772 654854
rect 589008 654618 589040 654854
rect 588420 619174 589040 654618
rect 588420 618938 588452 619174
rect 588688 618938 588772 619174
rect 589008 618938 589040 619174
rect 588420 618854 589040 618938
rect 588420 618618 588452 618854
rect 588688 618618 588772 618854
rect 589008 618618 589040 618854
rect 588420 583174 589040 618618
rect 588420 582938 588452 583174
rect 588688 582938 588772 583174
rect 589008 582938 589040 583174
rect 588420 582854 589040 582938
rect 588420 582618 588452 582854
rect 588688 582618 588772 582854
rect 589008 582618 589040 582854
rect 588420 547174 589040 582618
rect 588420 546938 588452 547174
rect 588688 546938 588772 547174
rect 589008 546938 589040 547174
rect 588420 546854 589040 546938
rect 588420 546618 588452 546854
rect 588688 546618 588772 546854
rect 589008 546618 589040 546854
rect 588420 511174 589040 546618
rect 588420 510938 588452 511174
rect 588688 510938 588772 511174
rect 589008 510938 589040 511174
rect 588420 510854 589040 510938
rect 588420 510618 588452 510854
rect 588688 510618 588772 510854
rect 589008 510618 589040 510854
rect 588420 475174 589040 510618
rect 588420 474938 588452 475174
rect 588688 474938 588772 475174
rect 589008 474938 589040 475174
rect 588420 474854 589040 474938
rect 588420 474618 588452 474854
rect 588688 474618 588772 474854
rect 589008 474618 589040 474854
rect 588420 439174 589040 474618
rect 588420 438938 588452 439174
rect 588688 438938 588772 439174
rect 589008 438938 589040 439174
rect 588420 438854 589040 438938
rect 588420 438618 588452 438854
rect 588688 438618 588772 438854
rect 589008 438618 589040 438854
rect 588420 403174 589040 438618
rect 588420 402938 588452 403174
rect 588688 402938 588772 403174
rect 589008 402938 589040 403174
rect 588420 402854 589040 402938
rect 588420 402618 588452 402854
rect 588688 402618 588772 402854
rect 589008 402618 589040 402854
rect 588420 367174 589040 402618
rect 588420 366938 588452 367174
rect 588688 366938 588772 367174
rect 589008 366938 589040 367174
rect 588420 366854 589040 366938
rect 588420 366618 588452 366854
rect 588688 366618 588772 366854
rect 589008 366618 589040 366854
rect 588420 331174 589040 366618
rect 588420 330938 588452 331174
rect 588688 330938 588772 331174
rect 589008 330938 589040 331174
rect 588420 330854 589040 330938
rect 588420 330618 588452 330854
rect 588688 330618 588772 330854
rect 589008 330618 589040 330854
rect 588420 295174 589040 330618
rect 588420 294938 588452 295174
rect 588688 294938 588772 295174
rect 589008 294938 589040 295174
rect 588420 294854 589040 294938
rect 588420 294618 588452 294854
rect 588688 294618 588772 294854
rect 589008 294618 589040 294854
rect 588420 259174 589040 294618
rect 588420 258938 588452 259174
rect 588688 258938 588772 259174
rect 589008 258938 589040 259174
rect 588420 258854 589040 258938
rect 588420 258618 588452 258854
rect 588688 258618 588772 258854
rect 589008 258618 589040 258854
rect 588420 223174 589040 258618
rect 588420 222938 588452 223174
rect 588688 222938 588772 223174
rect 589008 222938 589040 223174
rect 588420 222854 589040 222938
rect 588420 222618 588452 222854
rect 588688 222618 588772 222854
rect 589008 222618 589040 222854
rect 588420 187174 589040 222618
rect 588420 186938 588452 187174
rect 588688 186938 588772 187174
rect 589008 186938 589040 187174
rect 588420 186854 589040 186938
rect 588420 186618 588452 186854
rect 588688 186618 588772 186854
rect 589008 186618 589040 186854
rect 588420 151174 589040 186618
rect 588420 150938 588452 151174
rect 588688 150938 588772 151174
rect 589008 150938 589040 151174
rect 588420 150854 589040 150938
rect 588420 150618 588452 150854
rect 588688 150618 588772 150854
rect 589008 150618 589040 150854
rect 588420 115174 589040 150618
rect 588420 114938 588452 115174
rect 588688 114938 588772 115174
rect 589008 114938 589040 115174
rect 588420 114854 589040 114938
rect 588420 114618 588452 114854
rect 588688 114618 588772 114854
rect 589008 114618 589040 114854
rect 588420 79174 589040 114618
rect 588420 78938 588452 79174
rect 588688 78938 588772 79174
rect 589008 78938 589040 79174
rect 588420 78854 589040 78938
rect 588420 78618 588452 78854
rect 588688 78618 588772 78854
rect 589008 78618 589040 78854
rect 588420 43174 589040 78618
rect 588420 42938 588452 43174
rect 588688 42938 588772 43174
rect 589008 42938 589040 43174
rect 588420 42854 589040 42938
rect 588420 42618 588452 42854
rect 588688 42618 588772 42854
rect 589008 42618 589040 42854
rect 588420 7174 589040 42618
rect 588420 6938 588452 7174
rect 588688 6938 588772 7174
rect 589008 6938 589040 7174
rect 588420 6854 589040 6938
rect 588420 6618 588452 6854
rect 588688 6618 588772 6854
rect 589008 6618 589040 6854
rect 581514 -3692 581546 -3456
rect 581782 -3692 581866 -3456
rect 582102 -3692 582134 -3456
rect 581514 -3776 582134 -3692
rect 581514 -4012 581546 -3776
rect 581782 -4012 581866 -3776
rect 582102 -4012 582134 -3776
rect -8226 -6802 -8194 -6566
rect -7958 -6802 -7874 -6566
rect -7638 -6802 -7606 -6566
rect -8226 -6886 -7606 -6802
rect -8226 -7122 -8194 -6886
rect -7958 -7122 -7874 -6886
rect -7638 -7122 -7606 -6886
rect -8226 -7154 -7606 -7122
rect -11336 -9912 -11304 -9676
rect -11068 -9912 -10984 -9676
rect -10748 -9912 -10716 -9676
rect -11336 -9996 -10716 -9912
rect -11336 -10232 -11304 -9996
rect -11068 -10232 -10984 -9996
rect -10748 -10232 -10716 -9996
rect -11336 -10264 -10716 -10232
rect -14446 -13022 -14414 -12786
rect -14178 -13022 -14094 -12786
rect -13858 -13022 -13826 -12786
rect -14446 -13106 -13826 -13022
rect -14446 -13342 -14414 -13106
rect -14178 -13342 -14094 -13106
rect -13858 -13342 -13826 -13106
rect -14446 -13374 -13826 -13342
rect -17556 -16132 -17524 -15896
rect -17288 -16132 -17204 -15896
rect -16968 -16132 -16936 -15896
rect -17556 -16216 -16936 -16132
rect -17556 -16452 -17524 -16216
rect -17288 -16452 -17204 -16216
rect -16968 -16452 -16936 -16216
rect -17556 -16484 -16936 -16452
rect -20666 -19242 -20634 -19006
rect -20398 -19242 -20314 -19006
rect -20078 -19242 -20046 -19006
rect -20666 -19326 -20046 -19242
rect -20666 -19562 -20634 -19326
rect -20398 -19562 -20314 -19326
rect -20078 -19562 -20046 -19326
rect -20666 -19594 -20046 -19562
rect -23776 -22352 -23744 -22116
rect -23508 -22352 -23424 -22116
rect -23188 -22352 -23156 -22116
rect -23776 -22436 -23156 -22352
rect -23776 -22672 -23744 -22436
rect -23508 -22672 -23424 -22436
rect -23188 -22672 -23156 -22436
rect -23776 -22704 -23156 -22672
rect 581514 -22704 582134 -4012
rect 588420 -3456 589040 6618
rect 588420 -3692 588452 -3456
rect 588688 -3692 588772 -3456
rect 589008 -3692 589040 -3456
rect 588420 -3776 589040 -3692
rect 588420 -4012 588452 -3776
rect 588688 -4012 588772 -3776
rect 589008 -4012 589040 -3776
rect 588420 -4044 589040 -4012
rect 591530 694894 592150 710502
rect 591530 694658 591562 694894
rect 591798 694658 591882 694894
rect 592118 694658 592150 694894
rect 591530 694574 592150 694658
rect 591530 694338 591562 694574
rect 591798 694338 591882 694574
rect 592118 694338 592150 694574
rect 591530 658894 592150 694338
rect 591530 658658 591562 658894
rect 591798 658658 591882 658894
rect 592118 658658 592150 658894
rect 591530 658574 592150 658658
rect 591530 658338 591562 658574
rect 591798 658338 591882 658574
rect 592118 658338 592150 658574
rect 591530 622894 592150 658338
rect 591530 622658 591562 622894
rect 591798 622658 591882 622894
rect 592118 622658 592150 622894
rect 591530 622574 592150 622658
rect 591530 622338 591562 622574
rect 591798 622338 591882 622574
rect 592118 622338 592150 622574
rect 591530 586894 592150 622338
rect 591530 586658 591562 586894
rect 591798 586658 591882 586894
rect 592118 586658 592150 586894
rect 591530 586574 592150 586658
rect 591530 586338 591562 586574
rect 591798 586338 591882 586574
rect 592118 586338 592150 586574
rect 591530 550894 592150 586338
rect 591530 550658 591562 550894
rect 591798 550658 591882 550894
rect 592118 550658 592150 550894
rect 591530 550574 592150 550658
rect 591530 550338 591562 550574
rect 591798 550338 591882 550574
rect 592118 550338 592150 550574
rect 591530 514894 592150 550338
rect 591530 514658 591562 514894
rect 591798 514658 591882 514894
rect 592118 514658 592150 514894
rect 591530 514574 592150 514658
rect 591530 514338 591562 514574
rect 591798 514338 591882 514574
rect 592118 514338 592150 514574
rect 591530 478894 592150 514338
rect 591530 478658 591562 478894
rect 591798 478658 591882 478894
rect 592118 478658 592150 478894
rect 591530 478574 592150 478658
rect 591530 478338 591562 478574
rect 591798 478338 591882 478574
rect 592118 478338 592150 478574
rect 591530 442894 592150 478338
rect 591530 442658 591562 442894
rect 591798 442658 591882 442894
rect 592118 442658 592150 442894
rect 591530 442574 592150 442658
rect 591530 442338 591562 442574
rect 591798 442338 591882 442574
rect 592118 442338 592150 442574
rect 591530 406894 592150 442338
rect 591530 406658 591562 406894
rect 591798 406658 591882 406894
rect 592118 406658 592150 406894
rect 591530 406574 592150 406658
rect 591530 406338 591562 406574
rect 591798 406338 591882 406574
rect 592118 406338 592150 406574
rect 591530 370894 592150 406338
rect 591530 370658 591562 370894
rect 591798 370658 591882 370894
rect 592118 370658 592150 370894
rect 591530 370574 592150 370658
rect 591530 370338 591562 370574
rect 591798 370338 591882 370574
rect 592118 370338 592150 370574
rect 591530 334894 592150 370338
rect 591530 334658 591562 334894
rect 591798 334658 591882 334894
rect 592118 334658 592150 334894
rect 591530 334574 592150 334658
rect 591530 334338 591562 334574
rect 591798 334338 591882 334574
rect 592118 334338 592150 334574
rect 591530 298894 592150 334338
rect 591530 298658 591562 298894
rect 591798 298658 591882 298894
rect 592118 298658 592150 298894
rect 591530 298574 592150 298658
rect 591530 298338 591562 298574
rect 591798 298338 591882 298574
rect 592118 298338 592150 298574
rect 591530 262894 592150 298338
rect 591530 262658 591562 262894
rect 591798 262658 591882 262894
rect 592118 262658 592150 262894
rect 591530 262574 592150 262658
rect 591530 262338 591562 262574
rect 591798 262338 591882 262574
rect 592118 262338 592150 262574
rect 591530 226894 592150 262338
rect 591530 226658 591562 226894
rect 591798 226658 591882 226894
rect 592118 226658 592150 226894
rect 591530 226574 592150 226658
rect 591530 226338 591562 226574
rect 591798 226338 591882 226574
rect 592118 226338 592150 226574
rect 591530 190894 592150 226338
rect 591530 190658 591562 190894
rect 591798 190658 591882 190894
rect 592118 190658 592150 190894
rect 591530 190574 592150 190658
rect 591530 190338 591562 190574
rect 591798 190338 591882 190574
rect 592118 190338 592150 190574
rect 591530 154894 592150 190338
rect 591530 154658 591562 154894
rect 591798 154658 591882 154894
rect 592118 154658 592150 154894
rect 591530 154574 592150 154658
rect 591530 154338 591562 154574
rect 591798 154338 591882 154574
rect 592118 154338 592150 154574
rect 591530 118894 592150 154338
rect 591530 118658 591562 118894
rect 591798 118658 591882 118894
rect 592118 118658 592150 118894
rect 591530 118574 592150 118658
rect 591530 118338 591562 118574
rect 591798 118338 591882 118574
rect 592118 118338 592150 118574
rect 591530 82894 592150 118338
rect 591530 82658 591562 82894
rect 591798 82658 591882 82894
rect 592118 82658 592150 82894
rect 591530 82574 592150 82658
rect 591530 82338 591562 82574
rect 591798 82338 591882 82574
rect 592118 82338 592150 82574
rect 591530 46894 592150 82338
rect 591530 46658 591562 46894
rect 591798 46658 591882 46894
rect 592118 46658 592150 46894
rect 591530 46574 592150 46658
rect 591530 46338 591562 46574
rect 591798 46338 591882 46574
rect 592118 46338 592150 46574
rect 591530 10894 592150 46338
rect 591530 10658 591562 10894
rect 591798 10658 591882 10894
rect 592118 10658 592150 10894
rect 591530 10574 592150 10658
rect 591530 10338 591562 10574
rect 591798 10338 591882 10574
rect 592118 10338 592150 10574
rect 591530 -6566 592150 10338
rect 591530 -6802 591562 -6566
rect 591798 -6802 591882 -6566
rect 592118 -6802 592150 -6566
rect 591530 -6886 592150 -6802
rect 591530 -7122 591562 -6886
rect 591798 -7122 591882 -6886
rect 592118 -7122 592150 -6886
rect 591530 -7154 592150 -7122
rect 594640 698614 595260 713612
rect 594640 698378 594672 698614
rect 594908 698378 594992 698614
rect 595228 698378 595260 698614
rect 594640 698294 595260 698378
rect 594640 698058 594672 698294
rect 594908 698058 594992 698294
rect 595228 698058 595260 698294
rect 594640 662614 595260 698058
rect 594640 662378 594672 662614
rect 594908 662378 594992 662614
rect 595228 662378 595260 662614
rect 594640 662294 595260 662378
rect 594640 662058 594672 662294
rect 594908 662058 594992 662294
rect 595228 662058 595260 662294
rect 594640 626614 595260 662058
rect 594640 626378 594672 626614
rect 594908 626378 594992 626614
rect 595228 626378 595260 626614
rect 594640 626294 595260 626378
rect 594640 626058 594672 626294
rect 594908 626058 594992 626294
rect 595228 626058 595260 626294
rect 594640 590614 595260 626058
rect 594640 590378 594672 590614
rect 594908 590378 594992 590614
rect 595228 590378 595260 590614
rect 594640 590294 595260 590378
rect 594640 590058 594672 590294
rect 594908 590058 594992 590294
rect 595228 590058 595260 590294
rect 594640 554614 595260 590058
rect 594640 554378 594672 554614
rect 594908 554378 594992 554614
rect 595228 554378 595260 554614
rect 594640 554294 595260 554378
rect 594640 554058 594672 554294
rect 594908 554058 594992 554294
rect 595228 554058 595260 554294
rect 594640 518614 595260 554058
rect 594640 518378 594672 518614
rect 594908 518378 594992 518614
rect 595228 518378 595260 518614
rect 594640 518294 595260 518378
rect 594640 518058 594672 518294
rect 594908 518058 594992 518294
rect 595228 518058 595260 518294
rect 594640 482614 595260 518058
rect 594640 482378 594672 482614
rect 594908 482378 594992 482614
rect 595228 482378 595260 482614
rect 594640 482294 595260 482378
rect 594640 482058 594672 482294
rect 594908 482058 594992 482294
rect 595228 482058 595260 482294
rect 594640 446614 595260 482058
rect 594640 446378 594672 446614
rect 594908 446378 594992 446614
rect 595228 446378 595260 446614
rect 594640 446294 595260 446378
rect 594640 446058 594672 446294
rect 594908 446058 594992 446294
rect 595228 446058 595260 446294
rect 594640 410614 595260 446058
rect 594640 410378 594672 410614
rect 594908 410378 594992 410614
rect 595228 410378 595260 410614
rect 594640 410294 595260 410378
rect 594640 410058 594672 410294
rect 594908 410058 594992 410294
rect 595228 410058 595260 410294
rect 594640 374614 595260 410058
rect 594640 374378 594672 374614
rect 594908 374378 594992 374614
rect 595228 374378 595260 374614
rect 594640 374294 595260 374378
rect 594640 374058 594672 374294
rect 594908 374058 594992 374294
rect 595228 374058 595260 374294
rect 594640 338614 595260 374058
rect 594640 338378 594672 338614
rect 594908 338378 594992 338614
rect 595228 338378 595260 338614
rect 594640 338294 595260 338378
rect 594640 338058 594672 338294
rect 594908 338058 594992 338294
rect 595228 338058 595260 338294
rect 594640 302614 595260 338058
rect 594640 302378 594672 302614
rect 594908 302378 594992 302614
rect 595228 302378 595260 302614
rect 594640 302294 595260 302378
rect 594640 302058 594672 302294
rect 594908 302058 594992 302294
rect 595228 302058 595260 302294
rect 594640 266614 595260 302058
rect 594640 266378 594672 266614
rect 594908 266378 594992 266614
rect 595228 266378 595260 266614
rect 594640 266294 595260 266378
rect 594640 266058 594672 266294
rect 594908 266058 594992 266294
rect 595228 266058 595260 266294
rect 594640 230614 595260 266058
rect 594640 230378 594672 230614
rect 594908 230378 594992 230614
rect 595228 230378 595260 230614
rect 594640 230294 595260 230378
rect 594640 230058 594672 230294
rect 594908 230058 594992 230294
rect 595228 230058 595260 230294
rect 594640 194614 595260 230058
rect 594640 194378 594672 194614
rect 594908 194378 594992 194614
rect 595228 194378 595260 194614
rect 594640 194294 595260 194378
rect 594640 194058 594672 194294
rect 594908 194058 594992 194294
rect 595228 194058 595260 194294
rect 594640 158614 595260 194058
rect 594640 158378 594672 158614
rect 594908 158378 594992 158614
rect 595228 158378 595260 158614
rect 594640 158294 595260 158378
rect 594640 158058 594672 158294
rect 594908 158058 594992 158294
rect 595228 158058 595260 158294
rect 594640 122614 595260 158058
rect 594640 122378 594672 122614
rect 594908 122378 594992 122614
rect 595228 122378 595260 122614
rect 594640 122294 595260 122378
rect 594640 122058 594672 122294
rect 594908 122058 594992 122294
rect 595228 122058 595260 122294
rect 594640 86614 595260 122058
rect 594640 86378 594672 86614
rect 594908 86378 594992 86614
rect 595228 86378 595260 86614
rect 594640 86294 595260 86378
rect 594640 86058 594672 86294
rect 594908 86058 594992 86294
rect 595228 86058 595260 86294
rect 594640 50614 595260 86058
rect 594640 50378 594672 50614
rect 594908 50378 594992 50614
rect 595228 50378 595260 50614
rect 594640 50294 595260 50378
rect 594640 50058 594672 50294
rect 594908 50058 594992 50294
rect 595228 50058 595260 50294
rect 594640 14614 595260 50058
rect 594640 14378 594672 14614
rect 594908 14378 594992 14614
rect 595228 14378 595260 14614
rect 594640 14294 595260 14378
rect 594640 14058 594672 14294
rect 594908 14058 594992 14294
rect 595228 14058 595260 14294
rect 594640 -9676 595260 14058
rect 594640 -9912 594672 -9676
rect 594908 -9912 594992 -9676
rect 595228 -9912 595260 -9676
rect 594640 -9996 595260 -9912
rect 594640 -10232 594672 -9996
rect 594908 -10232 594992 -9996
rect 595228 -10232 595260 -9996
rect 594640 -10264 595260 -10232
rect 597750 666334 598370 716722
rect 597750 666098 597782 666334
rect 598018 666098 598102 666334
rect 598338 666098 598370 666334
rect 597750 666014 598370 666098
rect 597750 665778 597782 666014
rect 598018 665778 598102 666014
rect 598338 665778 598370 666014
rect 597750 630334 598370 665778
rect 597750 630098 597782 630334
rect 598018 630098 598102 630334
rect 598338 630098 598370 630334
rect 597750 630014 598370 630098
rect 597750 629778 597782 630014
rect 598018 629778 598102 630014
rect 598338 629778 598370 630014
rect 597750 594334 598370 629778
rect 597750 594098 597782 594334
rect 598018 594098 598102 594334
rect 598338 594098 598370 594334
rect 597750 594014 598370 594098
rect 597750 593778 597782 594014
rect 598018 593778 598102 594014
rect 598338 593778 598370 594014
rect 597750 558334 598370 593778
rect 597750 558098 597782 558334
rect 598018 558098 598102 558334
rect 598338 558098 598370 558334
rect 597750 558014 598370 558098
rect 597750 557778 597782 558014
rect 598018 557778 598102 558014
rect 598338 557778 598370 558014
rect 597750 522334 598370 557778
rect 597750 522098 597782 522334
rect 598018 522098 598102 522334
rect 598338 522098 598370 522334
rect 597750 522014 598370 522098
rect 597750 521778 597782 522014
rect 598018 521778 598102 522014
rect 598338 521778 598370 522014
rect 597750 486334 598370 521778
rect 597750 486098 597782 486334
rect 598018 486098 598102 486334
rect 598338 486098 598370 486334
rect 597750 486014 598370 486098
rect 597750 485778 597782 486014
rect 598018 485778 598102 486014
rect 598338 485778 598370 486014
rect 597750 450334 598370 485778
rect 597750 450098 597782 450334
rect 598018 450098 598102 450334
rect 598338 450098 598370 450334
rect 597750 450014 598370 450098
rect 597750 449778 597782 450014
rect 598018 449778 598102 450014
rect 598338 449778 598370 450014
rect 597750 414334 598370 449778
rect 597750 414098 597782 414334
rect 598018 414098 598102 414334
rect 598338 414098 598370 414334
rect 597750 414014 598370 414098
rect 597750 413778 597782 414014
rect 598018 413778 598102 414014
rect 598338 413778 598370 414014
rect 597750 378334 598370 413778
rect 597750 378098 597782 378334
rect 598018 378098 598102 378334
rect 598338 378098 598370 378334
rect 597750 378014 598370 378098
rect 597750 377778 597782 378014
rect 598018 377778 598102 378014
rect 598338 377778 598370 378014
rect 597750 342334 598370 377778
rect 597750 342098 597782 342334
rect 598018 342098 598102 342334
rect 598338 342098 598370 342334
rect 597750 342014 598370 342098
rect 597750 341778 597782 342014
rect 598018 341778 598102 342014
rect 598338 341778 598370 342014
rect 597750 306334 598370 341778
rect 597750 306098 597782 306334
rect 598018 306098 598102 306334
rect 598338 306098 598370 306334
rect 597750 306014 598370 306098
rect 597750 305778 597782 306014
rect 598018 305778 598102 306014
rect 598338 305778 598370 306014
rect 597750 270334 598370 305778
rect 597750 270098 597782 270334
rect 598018 270098 598102 270334
rect 598338 270098 598370 270334
rect 597750 270014 598370 270098
rect 597750 269778 597782 270014
rect 598018 269778 598102 270014
rect 598338 269778 598370 270014
rect 597750 234334 598370 269778
rect 597750 234098 597782 234334
rect 598018 234098 598102 234334
rect 598338 234098 598370 234334
rect 597750 234014 598370 234098
rect 597750 233778 597782 234014
rect 598018 233778 598102 234014
rect 598338 233778 598370 234014
rect 597750 198334 598370 233778
rect 597750 198098 597782 198334
rect 598018 198098 598102 198334
rect 598338 198098 598370 198334
rect 597750 198014 598370 198098
rect 597750 197778 597782 198014
rect 598018 197778 598102 198014
rect 598338 197778 598370 198014
rect 597750 162334 598370 197778
rect 597750 162098 597782 162334
rect 598018 162098 598102 162334
rect 598338 162098 598370 162334
rect 597750 162014 598370 162098
rect 597750 161778 597782 162014
rect 598018 161778 598102 162014
rect 598338 161778 598370 162014
rect 597750 126334 598370 161778
rect 597750 126098 597782 126334
rect 598018 126098 598102 126334
rect 598338 126098 598370 126334
rect 597750 126014 598370 126098
rect 597750 125778 597782 126014
rect 598018 125778 598102 126014
rect 598338 125778 598370 126014
rect 597750 90334 598370 125778
rect 597750 90098 597782 90334
rect 598018 90098 598102 90334
rect 598338 90098 598370 90334
rect 597750 90014 598370 90098
rect 597750 89778 597782 90014
rect 598018 89778 598102 90014
rect 598338 89778 598370 90014
rect 597750 54334 598370 89778
rect 597750 54098 597782 54334
rect 598018 54098 598102 54334
rect 598338 54098 598370 54334
rect 597750 54014 598370 54098
rect 597750 53778 597782 54014
rect 598018 53778 598102 54014
rect 598338 53778 598370 54014
rect 597750 18334 598370 53778
rect 597750 18098 597782 18334
rect 598018 18098 598102 18334
rect 598338 18098 598370 18334
rect 597750 18014 598370 18098
rect 597750 17778 597782 18014
rect 598018 17778 598102 18014
rect 598338 17778 598370 18014
rect 597750 -12786 598370 17778
rect 597750 -13022 597782 -12786
rect 598018 -13022 598102 -12786
rect 598338 -13022 598370 -12786
rect 597750 -13106 598370 -13022
rect 597750 -13342 597782 -13106
rect 598018 -13342 598102 -13106
rect 598338 -13342 598370 -13106
rect 597750 -13374 598370 -13342
rect 600860 670054 601480 719832
rect 600860 669818 600892 670054
rect 601128 669818 601212 670054
rect 601448 669818 601480 670054
rect 600860 669734 601480 669818
rect 600860 669498 600892 669734
rect 601128 669498 601212 669734
rect 601448 669498 601480 669734
rect 600860 634054 601480 669498
rect 600860 633818 600892 634054
rect 601128 633818 601212 634054
rect 601448 633818 601480 634054
rect 600860 633734 601480 633818
rect 600860 633498 600892 633734
rect 601128 633498 601212 633734
rect 601448 633498 601480 633734
rect 600860 598054 601480 633498
rect 600860 597818 600892 598054
rect 601128 597818 601212 598054
rect 601448 597818 601480 598054
rect 600860 597734 601480 597818
rect 600860 597498 600892 597734
rect 601128 597498 601212 597734
rect 601448 597498 601480 597734
rect 600860 562054 601480 597498
rect 600860 561818 600892 562054
rect 601128 561818 601212 562054
rect 601448 561818 601480 562054
rect 600860 561734 601480 561818
rect 600860 561498 600892 561734
rect 601128 561498 601212 561734
rect 601448 561498 601480 561734
rect 600860 526054 601480 561498
rect 600860 525818 600892 526054
rect 601128 525818 601212 526054
rect 601448 525818 601480 526054
rect 600860 525734 601480 525818
rect 600860 525498 600892 525734
rect 601128 525498 601212 525734
rect 601448 525498 601480 525734
rect 600860 490054 601480 525498
rect 600860 489818 600892 490054
rect 601128 489818 601212 490054
rect 601448 489818 601480 490054
rect 600860 489734 601480 489818
rect 600860 489498 600892 489734
rect 601128 489498 601212 489734
rect 601448 489498 601480 489734
rect 600860 454054 601480 489498
rect 600860 453818 600892 454054
rect 601128 453818 601212 454054
rect 601448 453818 601480 454054
rect 600860 453734 601480 453818
rect 600860 453498 600892 453734
rect 601128 453498 601212 453734
rect 601448 453498 601480 453734
rect 600860 418054 601480 453498
rect 600860 417818 600892 418054
rect 601128 417818 601212 418054
rect 601448 417818 601480 418054
rect 600860 417734 601480 417818
rect 600860 417498 600892 417734
rect 601128 417498 601212 417734
rect 601448 417498 601480 417734
rect 600860 382054 601480 417498
rect 600860 381818 600892 382054
rect 601128 381818 601212 382054
rect 601448 381818 601480 382054
rect 600860 381734 601480 381818
rect 600860 381498 600892 381734
rect 601128 381498 601212 381734
rect 601448 381498 601480 381734
rect 600860 346054 601480 381498
rect 600860 345818 600892 346054
rect 601128 345818 601212 346054
rect 601448 345818 601480 346054
rect 600860 345734 601480 345818
rect 600860 345498 600892 345734
rect 601128 345498 601212 345734
rect 601448 345498 601480 345734
rect 600860 310054 601480 345498
rect 600860 309818 600892 310054
rect 601128 309818 601212 310054
rect 601448 309818 601480 310054
rect 600860 309734 601480 309818
rect 600860 309498 600892 309734
rect 601128 309498 601212 309734
rect 601448 309498 601480 309734
rect 600860 274054 601480 309498
rect 600860 273818 600892 274054
rect 601128 273818 601212 274054
rect 601448 273818 601480 274054
rect 600860 273734 601480 273818
rect 600860 273498 600892 273734
rect 601128 273498 601212 273734
rect 601448 273498 601480 273734
rect 600860 238054 601480 273498
rect 600860 237818 600892 238054
rect 601128 237818 601212 238054
rect 601448 237818 601480 238054
rect 600860 237734 601480 237818
rect 600860 237498 600892 237734
rect 601128 237498 601212 237734
rect 601448 237498 601480 237734
rect 600860 202054 601480 237498
rect 600860 201818 600892 202054
rect 601128 201818 601212 202054
rect 601448 201818 601480 202054
rect 600860 201734 601480 201818
rect 600860 201498 600892 201734
rect 601128 201498 601212 201734
rect 601448 201498 601480 201734
rect 600860 166054 601480 201498
rect 600860 165818 600892 166054
rect 601128 165818 601212 166054
rect 601448 165818 601480 166054
rect 600860 165734 601480 165818
rect 600860 165498 600892 165734
rect 601128 165498 601212 165734
rect 601448 165498 601480 165734
rect 600860 130054 601480 165498
rect 600860 129818 600892 130054
rect 601128 129818 601212 130054
rect 601448 129818 601480 130054
rect 600860 129734 601480 129818
rect 600860 129498 600892 129734
rect 601128 129498 601212 129734
rect 601448 129498 601480 129734
rect 600860 94054 601480 129498
rect 600860 93818 600892 94054
rect 601128 93818 601212 94054
rect 601448 93818 601480 94054
rect 600860 93734 601480 93818
rect 600860 93498 600892 93734
rect 601128 93498 601212 93734
rect 601448 93498 601480 93734
rect 600860 58054 601480 93498
rect 600860 57818 600892 58054
rect 601128 57818 601212 58054
rect 601448 57818 601480 58054
rect 600860 57734 601480 57818
rect 600860 57498 600892 57734
rect 601128 57498 601212 57734
rect 601448 57498 601480 57734
rect 600860 -15896 601480 57498
rect 600860 -16132 600892 -15896
rect 601128 -16132 601212 -15896
rect 601448 -16132 601480 -15896
rect 600860 -16216 601480 -16132
rect 600860 -16452 600892 -16216
rect 601128 -16452 601212 -16216
rect 601448 -16452 601480 -16216
rect 600860 -16484 601480 -16452
rect 603970 673774 604590 722942
rect 603970 673538 604002 673774
rect 604238 673538 604322 673774
rect 604558 673538 604590 673774
rect 603970 673454 604590 673538
rect 603970 673218 604002 673454
rect 604238 673218 604322 673454
rect 604558 673218 604590 673454
rect 603970 637774 604590 673218
rect 603970 637538 604002 637774
rect 604238 637538 604322 637774
rect 604558 637538 604590 637774
rect 603970 637454 604590 637538
rect 603970 637218 604002 637454
rect 604238 637218 604322 637454
rect 604558 637218 604590 637454
rect 603970 601774 604590 637218
rect 603970 601538 604002 601774
rect 604238 601538 604322 601774
rect 604558 601538 604590 601774
rect 603970 601454 604590 601538
rect 603970 601218 604002 601454
rect 604238 601218 604322 601454
rect 604558 601218 604590 601454
rect 603970 565774 604590 601218
rect 603970 565538 604002 565774
rect 604238 565538 604322 565774
rect 604558 565538 604590 565774
rect 603970 565454 604590 565538
rect 603970 565218 604002 565454
rect 604238 565218 604322 565454
rect 604558 565218 604590 565454
rect 603970 529774 604590 565218
rect 603970 529538 604002 529774
rect 604238 529538 604322 529774
rect 604558 529538 604590 529774
rect 603970 529454 604590 529538
rect 603970 529218 604002 529454
rect 604238 529218 604322 529454
rect 604558 529218 604590 529454
rect 603970 493774 604590 529218
rect 603970 493538 604002 493774
rect 604238 493538 604322 493774
rect 604558 493538 604590 493774
rect 603970 493454 604590 493538
rect 603970 493218 604002 493454
rect 604238 493218 604322 493454
rect 604558 493218 604590 493454
rect 603970 457774 604590 493218
rect 603970 457538 604002 457774
rect 604238 457538 604322 457774
rect 604558 457538 604590 457774
rect 603970 457454 604590 457538
rect 603970 457218 604002 457454
rect 604238 457218 604322 457454
rect 604558 457218 604590 457454
rect 603970 421774 604590 457218
rect 603970 421538 604002 421774
rect 604238 421538 604322 421774
rect 604558 421538 604590 421774
rect 603970 421454 604590 421538
rect 603970 421218 604002 421454
rect 604238 421218 604322 421454
rect 604558 421218 604590 421454
rect 603970 385774 604590 421218
rect 603970 385538 604002 385774
rect 604238 385538 604322 385774
rect 604558 385538 604590 385774
rect 603970 385454 604590 385538
rect 603970 385218 604002 385454
rect 604238 385218 604322 385454
rect 604558 385218 604590 385454
rect 603970 349774 604590 385218
rect 603970 349538 604002 349774
rect 604238 349538 604322 349774
rect 604558 349538 604590 349774
rect 603970 349454 604590 349538
rect 603970 349218 604002 349454
rect 604238 349218 604322 349454
rect 604558 349218 604590 349454
rect 603970 313774 604590 349218
rect 603970 313538 604002 313774
rect 604238 313538 604322 313774
rect 604558 313538 604590 313774
rect 603970 313454 604590 313538
rect 603970 313218 604002 313454
rect 604238 313218 604322 313454
rect 604558 313218 604590 313454
rect 603970 277774 604590 313218
rect 603970 277538 604002 277774
rect 604238 277538 604322 277774
rect 604558 277538 604590 277774
rect 603970 277454 604590 277538
rect 603970 277218 604002 277454
rect 604238 277218 604322 277454
rect 604558 277218 604590 277454
rect 603970 241774 604590 277218
rect 603970 241538 604002 241774
rect 604238 241538 604322 241774
rect 604558 241538 604590 241774
rect 603970 241454 604590 241538
rect 603970 241218 604002 241454
rect 604238 241218 604322 241454
rect 604558 241218 604590 241454
rect 603970 205774 604590 241218
rect 603970 205538 604002 205774
rect 604238 205538 604322 205774
rect 604558 205538 604590 205774
rect 603970 205454 604590 205538
rect 603970 205218 604002 205454
rect 604238 205218 604322 205454
rect 604558 205218 604590 205454
rect 603970 169774 604590 205218
rect 603970 169538 604002 169774
rect 604238 169538 604322 169774
rect 604558 169538 604590 169774
rect 603970 169454 604590 169538
rect 603970 169218 604002 169454
rect 604238 169218 604322 169454
rect 604558 169218 604590 169454
rect 603970 133774 604590 169218
rect 603970 133538 604002 133774
rect 604238 133538 604322 133774
rect 604558 133538 604590 133774
rect 603970 133454 604590 133538
rect 603970 133218 604002 133454
rect 604238 133218 604322 133454
rect 604558 133218 604590 133454
rect 603970 97774 604590 133218
rect 603970 97538 604002 97774
rect 604238 97538 604322 97774
rect 604558 97538 604590 97774
rect 603970 97454 604590 97538
rect 603970 97218 604002 97454
rect 604238 97218 604322 97454
rect 604558 97218 604590 97454
rect 603970 61774 604590 97218
rect 603970 61538 604002 61774
rect 604238 61538 604322 61774
rect 604558 61538 604590 61774
rect 603970 61454 604590 61538
rect 603970 61218 604002 61454
rect 604238 61218 604322 61454
rect 604558 61218 604590 61454
rect 603970 25774 604590 61218
rect 603970 25538 604002 25774
rect 604238 25538 604322 25774
rect 604558 25538 604590 25774
rect 603970 25454 604590 25538
rect 603970 25218 604002 25454
rect 604238 25218 604322 25454
rect 604558 25218 604590 25454
rect 603970 -19006 604590 25218
rect 603970 -19242 604002 -19006
rect 604238 -19242 604322 -19006
rect 604558 -19242 604590 -19006
rect 603970 -19326 604590 -19242
rect 603970 -19562 604002 -19326
rect 604238 -19562 604322 -19326
rect 604558 -19562 604590 -19326
rect 603970 -19594 604590 -19562
rect 607080 677494 607700 726052
rect 607080 677258 607112 677494
rect 607348 677258 607432 677494
rect 607668 677258 607700 677494
rect 607080 677174 607700 677258
rect 607080 676938 607112 677174
rect 607348 676938 607432 677174
rect 607668 676938 607700 677174
rect 607080 641494 607700 676938
rect 607080 641258 607112 641494
rect 607348 641258 607432 641494
rect 607668 641258 607700 641494
rect 607080 641174 607700 641258
rect 607080 640938 607112 641174
rect 607348 640938 607432 641174
rect 607668 640938 607700 641174
rect 607080 605494 607700 640938
rect 607080 605258 607112 605494
rect 607348 605258 607432 605494
rect 607668 605258 607700 605494
rect 607080 605174 607700 605258
rect 607080 604938 607112 605174
rect 607348 604938 607432 605174
rect 607668 604938 607700 605174
rect 607080 569494 607700 604938
rect 607080 569258 607112 569494
rect 607348 569258 607432 569494
rect 607668 569258 607700 569494
rect 607080 569174 607700 569258
rect 607080 568938 607112 569174
rect 607348 568938 607432 569174
rect 607668 568938 607700 569174
rect 607080 533494 607700 568938
rect 607080 533258 607112 533494
rect 607348 533258 607432 533494
rect 607668 533258 607700 533494
rect 607080 533174 607700 533258
rect 607080 532938 607112 533174
rect 607348 532938 607432 533174
rect 607668 532938 607700 533174
rect 607080 497494 607700 532938
rect 607080 497258 607112 497494
rect 607348 497258 607432 497494
rect 607668 497258 607700 497494
rect 607080 497174 607700 497258
rect 607080 496938 607112 497174
rect 607348 496938 607432 497174
rect 607668 496938 607700 497174
rect 607080 461494 607700 496938
rect 607080 461258 607112 461494
rect 607348 461258 607432 461494
rect 607668 461258 607700 461494
rect 607080 461174 607700 461258
rect 607080 460938 607112 461174
rect 607348 460938 607432 461174
rect 607668 460938 607700 461174
rect 607080 425494 607700 460938
rect 607080 425258 607112 425494
rect 607348 425258 607432 425494
rect 607668 425258 607700 425494
rect 607080 425174 607700 425258
rect 607080 424938 607112 425174
rect 607348 424938 607432 425174
rect 607668 424938 607700 425174
rect 607080 389494 607700 424938
rect 607080 389258 607112 389494
rect 607348 389258 607432 389494
rect 607668 389258 607700 389494
rect 607080 389174 607700 389258
rect 607080 388938 607112 389174
rect 607348 388938 607432 389174
rect 607668 388938 607700 389174
rect 607080 353494 607700 388938
rect 607080 353258 607112 353494
rect 607348 353258 607432 353494
rect 607668 353258 607700 353494
rect 607080 353174 607700 353258
rect 607080 352938 607112 353174
rect 607348 352938 607432 353174
rect 607668 352938 607700 353174
rect 607080 317494 607700 352938
rect 607080 317258 607112 317494
rect 607348 317258 607432 317494
rect 607668 317258 607700 317494
rect 607080 317174 607700 317258
rect 607080 316938 607112 317174
rect 607348 316938 607432 317174
rect 607668 316938 607700 317174
rect 607080 281494 607700 316938
rect 607080 281258 607112 281494
rect 607348 281258 607432 281494
rect 607668 281258 607700 281494
rect 607080 281174 607700 281258
rect 607080 280938 607112 281174
rect 607348 280938 607432 281174
rect 607668 280938 607700 281174
rect 607080 245494 607700 280938
rect 607080 245258 607112 245494
rect 607348 245258 607432 245494
rect 607668 245258 607700 245494
rect 607080 245174 607700 245258
rect 607080 244938 607112 245174
rect 607348 244938 607432 245174
rect 607668 244938 607700 245174
rect 607080 209494 607700 244938
rect 607080 209258 607112 209494
rect 607348 209258 607432 209494
rect 607668 209258 607700 209494
rect 607080 209174 607700 209258
rect 607080 208938 607112 209174
rect 607348 208938 607432 209174
rect 607668 208938 607700 209174
rect 607080 173494 607700 208938
rect 607080 173258 607112 173494
rect 607348 173258 607432 173494
rect 607668 173258 607700 173494
rect 607080 173174 607700 173258
rect 607080 172938 607112 173174
rect 607348 172938 607432 173174
rect 607668 172938 607700 173174
rect 607080 137494 607700 172938
rect 607080 137258 607112 137494
rect 607348 137258 607432 137494
rect 607668 137258 607700 137494
rect 607080 137174 607700 137258
rect 607080 136938 607112 137174
rect 607348 136938 607432 137174
rect 607668 136938 607700 137174
rect 607080 101494 607700 136938
rect 607080 101258 607112 101494
rect 607348 101258 607432 101494
rect 607668 101258 607700 101494
rect 607080 101174 607700 101258
rect 607080 100938 607112 101174
rect 607348 100938 607432 101174
rect 607668 100938 607700 101174
rect 607080 65494 607700 100938
rect 607080 65258 607112 65494
rect 607348 65258 607432 65494
rect 607668 65258 607700 65494
rect 607080 65174 607700 65258
rect 607080 64938 607112 65174
rect 607348 64938 607432 65174
rect 607668 64938 607700 65174
rect 607080 29494 607700 64938
rect 607080 29258 607112 29494
rect 607348 29258 607432 29494
rect 607668 29258 607700 29494
rect 607080 29174 607700 29258
rect 607080 28938 607112 29174
rect 607348 28938 607432 29174
rect 607668 28938 607700 29174
rect 607080 -22116 607700 28938
rect 607080 -22352 607112 -22116
rect 607348 -22352 607432 -22116
rect 607668 -22352 607700 -22116
rect 607080 -22436 607700 -22352
rect 607080 -22672 607112 -22436
rect 607348 -22672 607432 -22436
rect 607668 -22672 607700 -22436
rect 607080 -22704 607700 -22672
<< via4 >>
rect -23744 726372 -23508 726608
rect -23424 726372 -23188 726608
rect -23744 726052 -23508 726288
rect -23424 726052 -23188 726288
rect -23744 677258 -23508 677494
rect -23424 677258 -23188 677494
rect -23744 676938 -23508 677174
rect -23424 676938 -23188 677174
rect -23744 641258 -23508 641494
rect -23424 641258 -23188 641494
rect -23744 640938 -23508 641174
rect -23424 640938 -23188 641174
rect -23744 605258 -23508 605494
rect -23424 605258 -23188 605494
rect -23744 604938 -23508 605174
rect -23424 604938 -23188 605174
rect -23744 569258 -23508 569494
rect -23424 569258 -23188 569494
rect -23744 568938 -23508 569174
rect -23424 568938 -23188 569174
rect -23744 533258 -23508 533494
rect -23424 533258 -23188 533494
rect -23744 532938 -23508 533174
rect -23424 532938 -23188 533174
rect -23744 497258 -23508 497494
rect -23424 497258 -23188 497494
rect -23744 496938 -23508 497174
rect -23424 496938 -23188 497174
rect -23744 461258 -23508 461494
rect -23424 461258 -23188 461494
rect -23744 460938 -23508 461174
rect -23424 460938 -23188 461174
rect -23744 425258 -23508 425494
rect -23424 425258 -23188 425494
rect -23744 424938 -23508 425174
rect -23424 424938 -23188 425174
rect -23744 389258 -23508 389494
rect -23424 389258 -23188 389494
rect -23744 388938 -23508 389174
rect -23424 388938 -23188 389174
rect -23744 353258 -23508 353494
rect -23424 353258 -23188 353494
rect -23744 352938 -23508 353174
rect -23424 352938 -23188 353174
rect -23744 317258 -23508 317494
rect -23424 317258 -23188 317494
rect -23744 316938 -23508 317174
rect -23424 316938 -23188 317174
rect -23744 281258 -23508 281494
rect -23424 281258 -23188 281494
rect -23744 280938 -23508 281174
rect -23424 280938 -23188 281174
rect -23744 245258 -23508 245494
rect -23424 245258 -23188 245494
rect -23744 244938 -23508 245174
rect -23424 244938 -23188 245174
rect -23744 209258 -23508 209494
rect -23424 209258 -23188 209494
rect -23744 208938 -23508 209174
rect -23424 208938 -23188 209174
rect -23744 173258 -23508 173494
rect -23424 173258 -23188 173494
rect -23744 172938 -23508 173174
rect -23424 172938 -23188 173174
rect -23744 137258 -23508 137494
rect -23424 137258 -23188 137494
rect -23744 136938 -23508 137174
rect -23424 136938 -23188 137174
rect -23744 101258 -23508 101494
rect -23424 101258 -23188 101494
rect -23744 100938 -23508 101174
rect -23424 100938 -23188 101174
rect -23744 65258 -23508 65494
rect -23424 65258 -23188 65494
rect -23744 64938 -23508 65174
rect -23424 64938 -23188 65174
rect -23744 29258 -23508 29494
rect -23424 29258 -23188 29494
rect -23744 28938 -23508 29174
rect -23424 28938 -23188 29174
rect -20634 723262 -20398 723498
rect -20314 723262 -20078 723498
rect -20634 722942 -20398 723178
rect -20314 722942 -20078 723178
rect -20634 673538 -20398 673774
rect -20314 673538 -20078 673774
rect -20634 673218 -20398 673454
rect -20314 673218 -20078 673454
rect -20634 637538 -20398 637774
rect -20314 637538 -20078 637774
rect -20634 637218 -20398 637454
rect -20314 637218 -20078 637454
rect -20634 601538 -20398 601774
rect -20314 601538 -20078 601774
rect -20634 601218 -20398 601454
rect -20314 601218 -20078 601454
rect -20634 565538 -20398 565774
rect -20314 565538 -20078 565774
rect -20634 565218 -20398 565454
rect -20314 565218 -20078 565454
rect -20634 529538 -20398 529774
rect -20314 529538 -20078 529774
rect -20634 529218 -20398 529454
rect -20314 529218 -20078 529454
rect -20634 493538 -20398 493774
rect -20314 493538 -20078 493774
rect -20634 493218 -20398 493454
rect -20314 493218 -20078 493454
rect -20634 457538 -20398 457774
rect -20314 457538 -20078 457774
rect -20634 457218 -20398 457454
rect -20314 457218 -20078 457454
rect -20634 421538 -20398 421774
rect -20314 421538 -20078 421774
rect -20634 421218 -20398 421454
rect -20314 421218 -20078 421454
rect -20634 385538 -20398 385774
rect -20314 385538 -20078 385774
rect -20634 385218 -20398 385454
rect -20314 385218 -20078 385454
rect -20634 349538 -20398 349774
rect -20314 349538 -20078 349774
rect -20634 349218 -20398 349454
rect -20314 349218 -20078 349454
rect -20634 313538 -20398 313774
rect -20314 313538 -20078 313774
rect -20634 313218 -20398 313454
rect -20314 313218 -20078 313454
rect -20634 277538 -20398 277774
rect -20314 277538 -20078 277774
rect -20634 277218 -20398 277454
rect -20314 277218 -20078 277454
rect -20634 241538 -20398 241774
rect -20314 241538 -20078 241774
rect -20634 241218 -20398 241454
rect -20314 241218 -20078 241454
rect -20634 205538 -20398 205774
rect -20314 205538 -20078 205774
rect -20634 205218 -20398 205454
rect -20314 205218 -20078 205454
rect -20634 169538 -20398 169774
rect -20314 169538 -20078 169774
rect -20634 169218 -20398 169454
rect -20314 169218 -20078 169454
rect -20634 133538 -20398 133774
rect -20314 133538 -20078 133774
rect -20634 133218 -20398 133454
rect -20314 133218 -20078 133454
rect -20634 97538 -20398 97774
rect -20314 97538 -20078 97774
rect -20634 97218 -20398 97454
rect -20314 97218 -20078 97454
rect -20634 61538 -20398 61774
rect -20314 61538 -20078 61774
rect -20634 61218 -20398 61454
rect -20314 61218 -20078 61454
rect -20634 25538 -20398 25774
rect -20314 25538 -20078 25774
rect -20634 25218 -20398 25454
rect -20314 25218 -20078 25454
rect -17524 720152 -17288 720388
rect -17204 720152 -16968 720388
rect -17524 719832 -17288 720068
rect -17204 719832 -16968 720068
rect -17524 669818 -17288 670054
rect -17204 669818 -16968 670054
rect -17524 669498 -17288 669734
rect -17204 669498 -16968 669734
rect -17524 633818 -17288 634054
rect -17204 633818 -16968 634054
rect -17524 633498 -17288 633734
rect -17204 633498 -16968 633734
rect -17524 597818 -17288 598054
rect -17204 597818 -16968 598054
rect -17524 597498 -17288 597734
rect -17204 597498 -16968 597734
rect -17524 561818 -17288 562054
rect -17204 561818 -16968 562054
rect -17524 561498 -17288 561734
rect -17204 561498 -16968 561734
rect -17524 525818 -17288 526054
rect -17204 525818 -16968 526054
rect -17524 525498 -17288 525734
rect -17204 525498 -16968 525734
rect -17524 489818 -17288 490054
rect -17204 489818 -16968 490054
rect -17524 489498 -17288 489734
rect -17204 489498 -16968 489734
rect -17524 453818 -17288 454054
rect -17204 453818 -16968 454054
rect -17524 453498 -17288 453734
rect -17204 453498 -16968 453734
rect -17524 417818 -17288 418054
rect -17204 417818 -16968 418054
rect -17524 417498 -17288 417734
rect -17204 417498 -16968 417734
rect -17524 381818 -17288 382054
rect -17204 381818 -16968 382054
rect -17524 381498 -17288 381734
rect -17204 381498 -16968 381734
rect -17524 345818 -17288 346054
rect -17204 345818 -16968 346054
rect -17524 345498 -17288 345734
rect -17204 345498 -16968 345734
rect -17524 309818 -17288 310054
rect -17204 309818 -16968 310054
rect -17524 309498 -17288 309734
rect -17204 309498 -16968 309734
rect -17524 273818 -17288 274054
rect -17204 273818 -16968 274054
rect -17524 273498 -17288 273734
rect -17204 273498 -16968 273734
rect -17524 237818 -17288 238054
rect -17204 237818 -16968 238054
rect -17524 237498 -17288 237734
rect -17204 237498 -16968 237734
rect -17524 201818 -17288 202054
rect -17204 201818 -16968 202054
rect -17524 201498 -17288 201734
rect -17204 201498 -16968 201734
rect -17524 165818 -17288 166054
rect -17204 165818 -16968 166054
rect -17524 165498 -17288 165734
rect -17204 165498 -16968 165734
rect -17524 129818 -17288 130054
rect -17204 129818 -16968 130054
rect -17524 129498 -17288 129734
rect -17204 129498 -16968 129734
rect -17524 93818 -17288 94054
rect -17204 93818 -16968 94054
rect -17524 93498 -17288 93734
rect -17204 93498 -16968 93734
rect -17524 57818 -17288 58054
rect -17204 57818 -16968 58054
rect -17524 57498 -17288 57734
rect -17204 57498 -16968 57734
rect -14414 717042 -14178 717278
rect -14094 717042 -13858 717278
rect -14414 716722 -14178 716958
rect -14094 716722 -13858 716958
rect -14414 666098 -14178 666334
rect -14094 666098 -13858 666334
rect -14414 665778 -14178 666014
rect -14094 665778 -13858 666014
rect -14414 630098 -14178 630334
rect -14094 630098 -13858 630334
rect -14414 629778 -14178 630014
rect -14094 629778 -13858 630014
rect -14414 594098 -14178 594334
rect -14094 594098 -13858 594334
rect -14414 593778 -14178 594014
rect -14094 593778 -13858 594014
rect -14414 558098 -14178 558334
rect -14094 558098 -13858 558334
rect -14414 557778 -14178 558014
rect -14094 557778 -13858 558014
rect -14414 522098 -14178 522334
rect -14094 522098 -13858 522334
rect -14414 521778 -14178 522014
rect -14094 521778 -13858 522014
rect -14414 486098 -14178 486334
rect -14094 486098 -13858 486334
rect -14414 485778 -14178 486014
rect -14094 485778 -13858 486014
rect -14414 450098 -14178 450334
rect -14094 450098 -13858 450334
rect -14414 449778 -14178 450014
rect -14094 449778 -13858 450014
rect -14414 414098 -14178 414334
rect -14094 414098 -13858 414334
rect -14414 413778 -14178 414014
rect -14094 413778 -13858 414014
rect -14414 378098 -14178 378334
rect -14094 378098 -13858 378334
rect -14414 377778 -14178 378014
rect -14094 377778 -13858 378014
rect -14414 342098 -14178 342334
rect -14094 342098 -13858 342334
rect -14414 341778 -14178 342014
rect -14094 341778 -13858 342014
rect -14414 306098 -14178 306334
rect -14094 306098 -13858 306334
rect -14414 305778 -14178 306014
rect -14094 305778 -13858 306014
rect -14414 270098 -14178 270334
rect -14094 270098 -13858 270334
rect -14414 269778 -14178 270014
rect -14094 269778 -13858 270014
rect -14414 234098 -14178 234334
rect -14094 234098 -13858 234334
rect -14414 233778 -14178 234014
rect -14094 233778 -13858 234014
rect -14414 198098 -14178 198334
rect -14094 198098 -13858 198334
rect -14414 197778 -14178 198014
rect -14094 197778 -13858 198014
rect -14414 162098 -14178 162334
rect -14094 162098 -13858 162334
rect -14414 161778 -14178 162014
rect -14094 161778 -13858 162014
rect -14414 126098 -14178 126334
rect -14094 126098 -13858 126334
rect -14414 125778 -14178 126014
rect -14094 125778 -13858 126014
rect -14414 90098 -14178 90334
rect -14094 90098 -13858 90334
rect -14414 89778 -14178 90014
rect -14094 89778 -13858 90014
rect -14414 54098 -14178 54334
rect -14094 54098 -13858 54334
rect -14414 53778 -14178 54014
rect -14094 53778 -13858 54014
rect -14414 18098 -14178 18334
rect -14094 18098 -13858 18334
rect -14414 17778 -14178 18014
rect -14094 17778 -13858 18014
rect -11304 713932 -11068 714168
rect -10984 713932 -10748 714168
rect -11304 713612 -11068 713848
rect -10984 713612 -10748 713848
rect -11304 698378 -11068 698614
rect -10984 698378 -10748 698614
rect -11304 698058 -11068 698294
rect -10984 698058 -10748 698294
rect -11304 662378 -11068 662614
rect -10984 662378 -10748 662614
rect -11304 662058 -11068 662294
rect -10984 662058 -10748 662294
rect -11304 626378 -11068 626614
rect -10984 626378 -10748 626614
rect -11304 626058 -11068 626294
rect -10984 626058 -10748 626294
rect -11304 590378 -11068 590614
rect -10984 590378 -10748 590614
rect -11304 590058 -11068 590294
rect -10984 590058 -10748 590294
rect -11304 554378 -11068 554614
rect -10984 554378 -10748 554614
rect -11304 554058 -11068 554294
rect -10984 554058 -10748 554294
rect -11304 518378 -11068 518614
rect -10984 518378 -10748 518614
rect -11304 518058 -11068 518294
rect -10984 518058 -10748 518294
rect -11304 482378 -11068 482614
rect -10984 482378 -10748 482614
rect -11304 482058 -11068 482294
rect -10984 482058 -10748 482294
rect -11304 446378 -11068 446614
rect -10984 446378 -10748 446614
rect -11304 446058 -11068 446294
rect -10984 446058 -10748 446294
rect -11304 410378 -11068 410614
rect -10984 410378 -10748 410614
rect -11304 410058 -11068 410294
rect -10984 410058 -10748 410294
rect -11304 374378 -11068 374614
rect -10984 374378 -10748 374614
rect -11304 374058 -11068 374294
rect -10984 374058 -10748 374294
rect -11304 338378 -11068 338614
rect -10984 338378 -10748 338614
rect -11304 338058 -11068 338294
rect -10984 338058 -10748 338294
rect -11304 302378 -11068 302614
rect -10984 302378 -10748 302614
rect -11304 302058 -11068 302294
rect -10984 302058 -10748 302294
rect -11304 266378 -11068 266614
rect -10984 266378 -10748 266614
rect -11304 266058 -11068 266294
rect -10984 266058 -10748 266294
rect -11304 230378 -11068 230614
rect -10984 230378 -10748 230614
rect -11304 230058 -11068 230294
rect -10984 230058 -10748 230294
rect -11304 194378 -11068 194614
rect -10984 194378 -10748 194614
rect -11304 194058 -11068 194294
rect -10984 194058 -10748 194294
rect -11304 158378 -11068 158614
rect -10984 158378 -10748 158614
rect -11304 158058 -11068 158294
rect -10984 158058 -10748 158294
rect -11304 122378 -11068 122614
rect -10984 122378 -10748 122614
rect -11304 122058 -11068 122294
rect -10984 122058 -10748 122294
rect -11304 86378 -11068 86614
rect -10984 86378 -10748 86614
rect -11304 86058 -11068 86294
rect -10984 86058 -10748 86294
rect -11304 50378 -11068 50614
rect -10984 50378 -10748 50614
rect -11304 50058 -11068 50294
rect -10984 50058 -10748 50294
rect -11304 14378 -11068 14614
rect -10984 14378 -10748 14614
rect -11304 14058 -11068 14294
rect -10984 14058 -10748 14294
rect -8194 710822 -7958 711058
rect -7874 710822 -7638 711058
rect -8194 710502 -7958 710738
rect -7874 710502 -7638 710738
rect -8194 694658 -7958 694894
rect -7874 694658 -7638 694894
rect -8194 694338 -7958 694574
rect -7874 694338 -7638 694574
rect -8194 658658 -7958 658894
rect -7874 658658 -7638 658894
rect -8194 658338 -7958 658574
rect -7874 658338 -7638 658574
rect -8194 622658 -7958 622894
rect -7874 622658 -7638 622894
rect -8194 622338 -7958 622574
rect -7874 622338 -7638 622574
rect -8194 586658 -7958 586894
rect -7874 586658 -7638 586894
rect -8194 586338 -7958 586574
rect -7874 586338 -7638 586574
rect -8194 550658 -7958 550894
rect -7874 550658 -7638 550894
rect -8194 550338 -7958 550574
rect -7874 550338 -7638 550574
rect -8194 514658 -7958 514894
rect -7874 514658 -7638 514894
rect -8194 514338 -7958 514574
rect -7874 514338 -7638 514574
rect -8194 478658 -7958 478894
rect -7874 478658 -7638 478894
rect -8194 478338 -7958 478574
rect -7874 478338 -7638 478574
rect -8194 442658 -7958 442894
rect -7874 442658 -7638 442894
rect -8194 442338 -7958 442574
rect -7874 442338 -7638 442574
rect -8194 406658 -7958 406894
rect -7874 406658 -7638 406894
rect -8194 406338 -7958 406574
rect -7874 406338 -7638 406574
rect -8194 370658 -7958 370894
rect -7874 370658 -7638 370894
rect -8194 370338 -7958 370574
rect -7874 370338 -7638 370574
rect -8194 334658 -7958 334894
rect -7874 334658 -7638 334894
rect -8194 334338 -7958 334574
rect -7874 334338 -7638 334574
rect -8194 298658 -7958 298894
rect -7874 298658 -7638 298894
rect -8194 298338 -7958 298574
rect -7874 298338 -7638 298574
rect -8194 262658 -7958 262894
rect -7874 262658 -7638 262894
rect -8194 262338 -7958 262574
rect -7874 262338 -7638 262574
rect -8194 226658 -7958 226894
rect -7874 226658 -7638 226894
rect -8194 226338 -7958 226574
rect -7874 226338 -7638 226574
rect -8194 190658 -7958 190894
rect -7874 190658 -7638 190894
rect -8194 190338 -7958 190574
rect -7874 190338 -7638 190574
rect -8194 154658 -7958 154894
rect -7874 154658 -7638 154894
rect -8194 154338 -7958 154574
rect -7874 154338 -7638 154574
rect -8194 118658 -7958 118894
rect -7874 118658 -7638 118894
rect -8194 118338 -7958 118574
rect -7874 118338 -7638 118574
rect -8194 82658 -7958 82894
rect -7874 82658 -7638 82894
rect -8194 82338 -7958 82574
rect -7874 82338 -7638 82574
rect -8194 46658 -7958 46894
rect -7874 46658 -7638 46894
rect -8194 46338 -7958 46574
rect -7874 46338 -7638 46574
rect -8194 10658 -7958 10894
rect -7874 10658 -7638 10894
rect -8194 10338 -7958 10574
rect -7874 10338 -7638 10574
rect -5084 707712 -4848 707948
rect -4764 707712 -4528 707948
rect -5084 707392 -4848 707628
rect -4764 707392 -4528 707628
rect 607112 726372 607348 726608
rect 607432 726372 607668 726608
rect 607112 726052 607348 726288
rect 607432 726052 607668 726288
rect 604002 723262 604238 723498
rect 604322 723262 604558 723498
rect 604002 722942 604238 723178
rect 604322 722942 604558 723178
rect 600892 720152 601128 720388
rect 601212 720152 601448 720388
rect 600892 719832 601128 720068
rect 601212 719832 601448 720068
rect 597782 717042 598018 717278
rect 598102 717042 598338 717278
rect 597782 716722 598018 716958
rect 598102 716722 598338 716958
rect 594672 713932 594908 714168
rect 594992 713932 595228 714168
rect 594672 713612 594908 713848
rect 594992 713612 595228 713848
rect 591562 710822 591798 711058
rect 591882 710822 592118 711058
rect 591562 710502 591798 710738
rect 591882 710502 592118 710738
rect 581546 707712 581782 707948
rect 581866 707712 582102 707948
rect 581546 707392 581782 707628
rect 581866 707392 582102 707628
rect -5084 690938 -4848 691174
rect -4764 690938 -4528 691174
rect -5084 690618 -4848 690854
rect -4764 690618 -4528 690854
rect -5084 654938 -4848 655174
rect -4764 654938 -4528 655174
rect -5084 654618 -4848 654854
rect -4764 654618 -4528 654854
rect -5084 618938 -4848 619174
rect -4764 618938 -4528 619174
rect -5084 618618 -4848 618854
rect -4764 618618 -4528 618854
rect -5084 582938 -4848 583174
rect -4764 582938 -4528 583174
rect -5084 582618 -4848 582854
rect -4764 582618 -4528 582854
rect -5084 546938 -4848 547174
rect -4764 546938 -4528 547174
rect -5084 546618 -4848 546854
rect -4764 546618 -4528 546854
rect -5084 510938 -4848 511174
rect -4764 510938 -4528 511174
rect -5084 510618 -4848 510854
rect -4764 510618 -4528 510854
rect -5084 474938 -4848 475174
rect -4764 474938 -4528 475174
rect -5084 474618 -4848 474854
rect -4764 474618 -4528 474854
rect -5084 438938 -4848 439174
rect -4764 438938 -4528 439174
rect -5084 438618 -4848 438854
rect -4764 438618 -4528 438854
rect -5084 402938 -4848 403174
rect -4764 402938 -4528 403174
rect -5084 402618 -4848 402854
rect -4764 402618 -4528 402854
rect -5084 366938 -4848 367174
rect -4764 366938 -4528 367174
rect -5084 366618 -4848 366854
rect -4764 366618 -4528 366854
rect -5084 330938 -4848 331174
rect -4764 330938 -4528 331174
rect -5084 330618 -4848 330854
rect -4764 330618 -4528 330854
rect -5084 294938 -4848 295174
rect -4764 294938 -4528 295174
rect -5084 294618 -4848 294854
rect -4764 294618 -4528 294854
rect -5084 258938 -4848 259174
rect -4764 258938 -4528 259174
rect -5084 258618 -4848 258854
rect -4764 258618 -4528 258854
rect -5084 222938 -4848 223174
rect -4764 222938 -4528 223174
rect -5084 222618 -4848 222854
rect -4764 222618 -4528 222854
rect -5084 186938 -4848 187174
rect -4764 186938 -4528 187174
rect -5084 186618 -4848 186854
rect -4764 186618 -4528 186854
rect -5084 150938 -4848 151174
rect -4764 150938 -4528 151174
rect -5084 150618 -4848 150854
rect -4764 150618 -4528 150854
rect -5084 114938 -4848 115174
rect -4764 114938 -4528 115174
rect -5084 114618 -4848 114854
rect -4764 114618 -4528 114854
rect -5084 78938 -4848 79174
rect -4764 78938 -4528 79174
rect -5084 78618 -4848 78854
rect -4764 78618 -4528 78854
rect -5084 42938 -4848 43174
rect -4764 42938 -4528 43174
rect -5084 42618 -4848 42854
rect -4764 42618 -4528 42854
rect -5084 6938 -4848 7174
rect -4764 6938 -4528 7174
rect -5084 6618 -4848 6854
rect -4764 6618 -4528 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect 7876 693480 8112 693716
rect 8196 693480 8432 693716
rect 7876 693160 8112 693396
rect 8196 693160 8432 693396
rect 38032 693480 38268 693716
rect 38352 693480 38588 693716
rect 38032 693160 38268 693396
rect 38352 693160 38588 693396
rect 74032 693480 74268 693716
rect 74352 693480 74588 693716
rect 74032 693160 74268 693396
rect 74352 693160 74588 693396
rect 110032 693480 110268 693716
rect 110352 693480 110588 693716
rect 110032 693160 110268 693396
rect 110352 693160 110588 693396
rect 146032 693480 146268 693716
rect 146352 693480 146588 693716
rect 146032 693160 146268 693396
rect 146352 693160 146588 693396
rect 182032 693480 182268 693716
rect 182352 693480 182588 693716
rect 182032 693160 182268 693396
rect 182352 693160 182588 693396
rect 218032 693480 218268 693716
rect 218352 693480 218588 693716
rect 218032 693160 218268 693396
rect 218352 693160 218588 693396
rect 254032 693480 254268 693716
rect 254352 693480 254588 693716
rect 254032 693160 254268 693396
rect 254352 693160 254588 693396
rect 290032 693480 290268 693716
rect 290352 693480 290588 693716
rect 290032 693160 290268 693396
rect 290352 693160 290588 693396
rect 326032 693480 326268 693716
rect 326352 693480 326588 693716
rect 326032 693160 326268 693396
rect 326352 693160 326588 693396
rect 362032 693480 362268 693716
rect 362352 693480 362588 693716
rect 362032 693160 362268 693396
rect 362352 693160 362588 693396
rect 398032 693480 398268 693716
rect 398352 693480 398588 693716
rect 398032 693160 398268 693396
rect 398352 693160 398588 693396
rect 434032 693480 434268 693716
rect 434352 693480 434588 693716
rect 434032 693160 434268 693396
rect 434352 693160 434588 693396
rect 470032 693480 470268 693716
rect 470352 693480 470588 693716
rect 470032 693160 470268 693396
rect 470352 693160 470588 693396
rect 506032 693480 506268 693716
rect 506352 693480 506588 693716
rect 506032 693160 506268 693396
rect 506352 693160 506588 693396
rect 542032 693480 542268 693716
rect 542352 693480 542588 693716
rect 542032 693160 542268 693396
rect 542352 693160 542588 693396
rect 571532 693480 571768 693716
rect 571852 693480 572088 693716
rect 571532 693160 571768 693396
rect 571852 693160 572088 693396
rect 9116 692240 9352 692476
rect 9436 692240 9672 692476
rect 9116 691920 9352 692156
rect 9436 691920 9672 692156
rect 56652 692240 56888 692476
rect 56972 692240 57208 692476
rect 56652 691920 56888 692156
rect 56972 691920 57208 692156
rect 92652 692240 92888 692476
rect 92972 692240 93208 692476
rect 92652 691920 92888 692156
rect 92972 691920 93208 692156
rect 128652 692240 128888 692476
rect 128972 692240 129208 692476
rect 128652 691920 128888 692156
rect 128972 691920 129208 692156
rect 164652 692240 164888 692476
rect 164972 692240 165208 692476
rect 164652 691920 164888 692156
rect 164972 691920 165208 692156
rect 200652 692240 200888 692476
rect 200972 692240 201208 692476
rect 200652 691920 200888 692156
rect 200972 691920 201208 692156
rect 236652 692240 236888 692476
rect 236972 692240 237208 692476
rect 236652 691920 236888 692156
rect 236972 691920 237208 692156
rect 272652 692240 272888 692476
rect 272972 692240 273208 692476
rect 272652 691920 272888 692156
rect 272972 691920 273208 692156
rect 308652 692240 308888 692476
rect 308972 692240 309208 692476
rect 308652 691920 308888 692156
rect 308972 691920 309208 692156
rect 344652 692240 344888 692476
rect 344972 692240 345208 692476
rect 344652 691920 344888 692156
rect 344972 691920 345208 692156
rect 380652 692240 380888 692476
rect 380972 692240 381208 692476
rect 380652 691920 380888 692156
rect 380972 691920 381208 692156
rect 416652 692240 416888 692476
rect 416972 692240 417208 692476
rect 416652 691920 416888 692156
rect 416972 691920 417208 692156
rect 452652 692240 452888 692476
rect 452972 692240 453208 692476
rect 452652 691920 452888 692156
rect 452972 691920 453208 692156
rect 488652 692240 488888 692476
rect 488972 692240 489208 692476
rect 488652 691920 488888 692156
rect 488972 691920 489208 692156
rect 524652 692240 524888 692476
rect 524972 692240 525208 692476
rect 524652 691920 524888 692156
rect 524972 691920 525208 692156
rect 560652 692240 560888 692476
rect 560972 692240 561208 692476
rect 560652 691920 560888 692156
rect 560972 691920 561208 692156
rect 570292 692240 570528 692476
rect 570612 692240 570848 692476
rect 570292 691920 570528 692156
rect 570612 691920 570848 692156
rect 588452 707712 588688 707948
rect 588772 707712 589008 707948
rect 588452 707392 588688 707628
rect 588772 707392 589008 707628
rect 7876 690938 8112 691174
rect 8196 690938 8432 691174
rect 7876 690618 8112 690854
rect 8196 690618 8432 690854
rect 38032 690938 38268 691174
rect 38352 690938 38588 691174
rect 38032 690618 38268 690854
rect 38352 690618 38588 690854
rect 74032 690938 74268 691174
rect 74352 690938 74588 691174
rect 74032 690618 74268 690854
rect 74352 690618 74588 690854
rect 110032 690938 110268 691174
rect 110352 690938 110588 691174
rect 110032 690618 110268 690854
rect 110352 690618 110588 690854
rect 146032 690938 146268 691174
rect 146352 690938 146588 691174
rect 146032 690618 146268 690854
rect 146352 690618 146588 690854
rect 182032 690938 182268 691174
rect 182352 690938 182588 691174
rect 182032 690618 182268 690854
rect 182352 690618 182588 690854
rect 218032 690938 218268 691174
rect 218352 690938 218588 691174
rect 218032 690618 218268 690854
rect 218352 690618 218588 690854
rect 254032 690938 254268 691174
rect 254352 690938 254588 691174
rect 254032 690618 254268 690854
rect 254352 690618 254588 690854
rect 290032 690938 290268 691174
rect 290352 690938 290588 691174
rect 290032 690618 290268 690854
rect 290352 690618 290588 690854
rect 326032 690938 326268 691174
rect 326352 690938 326588 691174
rect 326032 690618 326268 690854
rect 326352 690618 326588 690854
rect 362032 690938 362268 691174
rect 362352 690938 362588 691174
rect 362032 690618 362268 690854
rect 362352 690618 362588 690854
rect 398032 690938 398268 691174
rect 398352 690938 398588 691174
rect 398032 690618 398268 690854
rect 398352 690618 398588 690854
rect 434032 690938 434268 691174
rect 434352 690938 434588 691174
rect 434032 690618 434268 690854
rect 434352 690618 434588 690854
rect 470032 690938 470268 691174
rect 470352 690938 470588 691174
rect 470032 690618 470268 690854
rect 470352 690618 470588 690854
rect 506032 690938 506268 691174
rect 506352 690938 506588 691174
rect 506032 690618 506268 690854
rect 506352 690618 506588 690854
rect 542032 690938 542268 691174
rect 542352 690938 542588 691174
rect 542032 690618 542268 690854
rect 542352 690618 542588 690854
rect 571532 690938 571768 691174
rect 571852 690938 572088 691174
rect 571532 690618 571768 690854
rect 571852 690618 572088 690854
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect 9116 687218 9352 687454
rect 9436 687218 9672 687454
rect 9116 686898 9352 687134
rect 9436 686898 9672 687134
rect 56652 687218 56888 687454
rect 56972 687218 57208 687454
rect 56652 686898 56888 687134
rect 56972 686898 57208 687134
rect 92652 687218 92888 687454
rect 92972 687218 93208 687454
rect 92652 686898 92888 687134
rect 92972 686898 93208 687134
rect 128652 687218 128888 687454
rect 128972 687218 129208 687454
rect 128652 686898 128888 687134
rect 128972 686898 129208 687134
rect 164652 687218 164888 687454
rect 164972 687218 165208 687454
rect 164652 686898 164888 687134
rect 164972 686898 165208 687134
rect 200652 687218 200888 687454
rect 200972 687218 201208 687454
rect 200652 686898 200888 687134
rect 200972 686898 201208 687134
rect 236652 687218 236888 687454
rect 236972 687218 237208 687454
rect 236652 686898 236888 687134
rect 236972 686898 237208 687134
rect 272652 687218 272888 687454
rect 272972 687218 273208 687454
rect 272652 686898 272888 687134
rect 272972 686898 273208 687134
rect 308652 687218 308888 687454
rect 308972 687218 309208 687454
rect 308652 686898 308888 687134
rect 308972 686898 309208 687134
rect 344652 687218 344888 687454
rect 344972 687218 345208 687454
rect 344652 686898 344888 687134
rect 344972 686898 345208 687134
rect 380652 687218 380888 687454
rect 380972 687218 381208 687454
rect 380652 686898 380888 687134
rect 380972 686898 381208 687134
rect 416652 687218 416888 687454
rect 416972 687218 417208 687454
rect 416652 686898 416888 687134
rect 416972 686898 417208 687134
rect 452652 687218 452888 687454
rect 452972 687218 453208 687454
rect 452652 686898 452888 687134
rect 452972 686898 453208 687134
rect 488652 687218 488888 687454
rect 488972 687218 489208 687454
rect 488652 686898 488888 687134
rect 488972 686898 489208 687134
rect 524652 687218 524888 687454
rect 524972 687218 525208 687454
rect 524652 686898 524888 687134
rect 524972 686898 525208 687134
rect 560652 687218 560888 687454
rect 560972 687218 561208 687454
rect 560652 686898 560888 687134
rect 560972 686898 561208 687134
rect 570292 687218 570528 687454
rect 570612 687218 570848 687454
rect 570292 686898 570528 687134
rect 570612 686898 570848 687134
rect 7876 654938 8112 655174
rect 8196 654938 8432 655174
rect 7876 654618 8112 654854
rect 8196 654618 8432 654854
rect 38032 654938 38268 655174
rect 38352 654938 38588 655174
rect 38032 654618 38268 654854
rect 38352 654618 38588 654854
rect 74032 654938 74268 655174
rect 74352 654938 74588 655174
rect 74032 654618 74268 654854
rect 74352 654618 74588 654854
rect 110032 654938 110268 655174
rect 110352 654938 110588 655174
rect 110032 654618 110268 654854
rect 110352 654618 110588 654854
rect 146032 654938 146268 655174
rect 146352 654938 146588 655174
rect 146032 654618 146268 654854
rect 146352 654618 146588 654854
rect 182032 654938 182268 655174
rect 182352 654938 182588 655174
rect 182032 654618 182268 654854
rect 182352 654618 182588 654854
rect 218032 654938 218268 655174
rect 218352 654938 218588 655174
rect 218032 654618 218268 654854
rect 218352 654618 218588 654854
rect 254032 654938 254268 655174
rect 254352 654938 254588 655174
rect 254032 654618 254268 654854
rect 254352 654618 254588 654854
rect 290032 654938 290268 655174
rect 290352 654938 290588 655174
rect 290032 654618 290268 654854
rect 290352 654618 290588 654854
rect 326032 654938 326268 655174
rect 326352 654938 326588 655174
rect 326032 654618 326268 654854
rect 326352 654618 326588 654854
rect 362032 654938 362268 655174
rect 362352 654938 362588 655174
rect 362032 654618 362268 654854
rect 362352 654618 362588 654854
rect 398032 654938 398268 655174
rect 398352 654938 398588 655174
rect 398032 654618 398268 654854
rect 398352 654618 398588 654854
rect 434032 654938 434268 655174
rect 434352 654938 434588 655174
rect 434032 654618 434268 654854
rect 434352 654618 434588 654854
rect 470032 654938 470268 655174
rect 470352 654938 470588 655174
rect 470032 654618 470268 654854
rect 470352 654618 470588 654854
rect 506032 654938 506268 655174
rect 506352 654938 506588 655174
rect 506032 654618 506268 654854
rect 506352 654618 506588 654854
rect 542032 654938 542268 655174
rect 542352 654938 542588 655174
rect 542032 654618 542268 654854
rect 542352 654618 542588 654854
rect 571532 654938 571768 655174
rect 571852 654938 572088 655174
rect 571532 654618 571768 654854
rect 571852 654618 572088 654854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect 9116 651218 9352 651454
rect 9436 651218 9672 651454
rect 9116 650898 9352 651134
rect 9436 650898 9672 651134
rect 56652 651218 56888 651454
rect 56972 651218 57208 651454
rect 56652 650898 56888 651134
rect 56972 650898 57208 651134
rect 92652 651218 92888 651454
rect 92972 651218 93208 651454
rect 92652 650898 92888 651134
rect 92972 650898 93208 651134
rect 128652 651218 128888 651454
rect 128972 651218 129208 651454
rect 128652 650898 128888 651134
rect 128972 650898 129208 651134
rect 164652 651218 164888 651454
rect 164972 651218 165208 651454
rect 164652 650898 164888 651134
rect 164972 650898 165208 651134
rect 200652 651218 200888 651454
rect 200972 651218 201208 651454
rect 200652 650898 200888 651134
rect 200972 650898 201208 651134
rect 236652 651218 236888 651454
rect 236972 651218 237208 651454
rect 236652 650898 236888 651134
rect 236972 650898 237208 651134
rect 272652 651218 272888 651454
rect 272972 651218 273208 651454
rect 272652 650898 272888 651134
rect 272972 650898 273208 651134
rect 308652 651218 308888 651454
rect 308972 651218 309208 651454
rect 308652 650898 308888 651134
rect 308972 650898 309208 651134
rect 344652 651218 344888 651454
rect 344972 651218 345208 651454
rect 344652 650898 344888 651134
rect 344972 650898 345208 651134
rect 380652 651218 380888 651454
rect 380972 651218 381208 651454
rect 380652 650898 380888 651134
rect 380972 650898 381208 651134
rect 416652 651218 416888 651454
rect 416972 651218 417208 651454
rect 416652 650898 416888 651134
rect 416972 650898 417208 651134
rect 452652 651218 452888 651454
rect 452972 651218 453208 651454
rect 452652 650898 452888 651134
rect 452972 650898 453208 651134
rect 488652 651218 488888 651454
rect 488972 651218 489208 651454
rect 488652 650898 488888 651134
rect 488972 650898 489208 651134
rect 524652 651218 524888 651454
rect 524972 651218 525208 651454
rect 524652 650898 524888 651134
rect 524972 650898 525208 651134
rect 560652 651218 560888 651454
rect 560972 651218 561208 651454
rect 560652 650898 560888 651134
rect 560972 650898 561208 651134
rect 570292 651218 570528 651454
rect 570612 651218 570848 651454
rect 570292 650898 570528 651134
rect 570612 650898 570848 651134
rect 7876 618938 8112 619174
rect 8196 618938 8432 619174
rect 7876 618618 8112 618854
rect 8196 618618 8432 618854
rect 38032 618938 38268 619174
rect 38352 618938 38588 619174
rect 38032 618618 38268 618854
rect 38352 618618 38588 618854
rect 74032 618938 74268 619174
rect 74352 618938 74588 619174
rect 74032 618618 74268 618854
rect 74352 618618 74588 618854
rect 110032 618938 110268 619174
rect 110352 618938 110588 619174
rect 110032 618618 110268 618854
rect 110352 618618 110588 618854
rect 146032 618938 146268 619174
rect 146352 618938 146588 619174
rect 146032 618618 146268 618854
rect 146352 618618 146588 618854
rect 182032 618938 182268 619174
rect 182352 618938 182588 619174
rect 182032 618618 182268 618854
rect 182352 618618 182588 618854
rect 218032 618938 218268 619174
rect 218352 618938 218588 619174
rect 218032 618618 218268 618854
rect 218352 618618 218588 618854
rect 254032 618938 254268 619174
rect 254352 618938 254588 619174
rect 254032 618618 254268 618854
rect 254352 618618 254588 618854
rect 290032 618938 290268 619174
rect 290352 618938 290588 619174
rect 290032 618618 290268 618854
rect 290352 618618 290588 618854
rect 326032 618938 326268 619174
rect 326352 618938 326588 619174
rect 326032 618618 326268 618854
rect 326352 618618 326588 618854
rect 362032 618938 362268 619174
rect 362352 618938 362588 619174
rect 362032 618618 362268 618854
rect 362352 618618 362588 618854
rect 398032 618938 398268 619174
rect 398352 618938 398588 619174
rect 398032 618618 398268 618854
rect 398352 618618 398588 618854
rect 434032 618938 434268 619174
rect 434352 618938 434588 619174
rect 434032 618618 434268 618854
rect 434352 618618 434588 618854
rect 470032 618938 470268 619174
rect 470352 618938 470588 619174
rect 470032 618618 470268 618854
rect 470352 618618 470588 618854
rect 506032 618938 506268 619174
rect 506352 618938 506588 619174
rect 506032 618618 506268 618854
rect 506352 618618 506588 618854
rect 542032 618938 542268 619174
rect 542352 618938 542588 619174
rect 542032 618618 542268 618854
rect 542352 618618 542588 618854
rect 571532 618938 571768 619174
rect 571852 618938 572088 619174
rect 571532 618618 571768 618854
rect 571852 618618 572088 618854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect 9116 615218 9352 615454
rect 9436 615218 9672 615454
rect 9116 614898 9352 615134
rect 9436 614898 9672 615134
rect 56652 615218 56888 615454
rect 56972 615218 57208 615454
rect 56652 614898 56888 615134
rect 56972 614898 57208 615134
rect 92652 615218 92888 615454
rect 92972 615218 93208 615454
rect 92652 614898 92888 615134
rect 92972 614898 93208 615134
rect 128652 615218 128888 615454
rect 128972 615218 129208 615454
rect 128652 614898 128888 615134
rect 128972 614898 129208 615134
rect 164652 615218 164888 615454
rect 164972 615218 165208 615454
rect 164652 614898 164888 615134
rect 164972 614898 165208 615134
rect 200652 615218 200888 615454
rect 200972 615218 201208 615454
rect 200652 614898 200888 615134
rect 200972 614898 201208 615134
rect 236652 615218 236888 615454
rect 236972 615218 237208 615454
rect 236652 614898 236888 615134
rect 236972 614898 237208 615134
rect 272652 615218 272888 615454
rect 272972 615218 273208 615454
rect 272652 614898 272888 615134
rect 272972 614898 273208 615134
rect 308652 615218 308888 615454
rect 308972 615218 309208 615454
rect 308652 614898 308888 615134
rect 308972 614898 309208 615134
rect 344652 615218 344888 615454
rect 344972 615218 345208 615454
rect 344652 614898 344888 615134
rect 344972 614898 345208 615134
rect 380652 615218 380888 615454
rect 380972 615218 381208 615454
rect 380652 614898 380888 615134
rect 380972 614898 381208 615134
rect 416652 615218 416888 615454
rect 416972 615218 417208 615454
rect 416652 614898 416888 615134
rect 416972 614898 417208 615134
rect 452652 615218 452888 615454
rect 452972 615218 453208 615454
rect 452652 614898 452888 615134
rect 452972 614898 453208 615134
rect 488652 615218 488888 615454
rect 488972 615218 489208 615454
rect 488652 614898 488888 615134
rect 488972 614898 489208 615134
rect 524652 615218 524888 615454
rect 524972 615218 525208 615454
rect 524652 614898 524888 615134
rect 524972 614898 525208 615134
rect 560652 615218 560888 615454
rect 560972 615218 561208 615454
rect 560652 614898 560888 615134
rect 560972 614898 561208 615134
rect 570292 615218 570528 615454
rect 570612 615218 570848 615454
rect 570292 614898 570528 615134
rect 570612 614898 570848 615134
rect 7876 582938 8112 583174
rect 8196 582938 8432 583174
rect 7876 582618 8112 582854
rect 8196 582618 8432 582854
rect 38032 582938 38268 583174
rect 38352 582938 38588 583174
rect 38032 582618 38268 582854
rect 38352 582618 38588 582854
rect 74032 582938 74268 583174
rect 74352 582938 74588 583174
rect 74032 582618 74268 582854
rect 74352 582618 74588 582854
rect 110032 582938 110268 583174
rect 110352 582938 110588 583174
rect 110032 582618 110268 582854
rect 110352 582618 110588 582854
rect 146032 582938 146268 583174
rect 146352 582938 146588 583174
rect 146032 582618 146268 582854
rect 146352 582618 146588 582854
rect 182032 582938 182268 583174
rect 182352 582938 182588 583174
rect 182032 582618 182268 582854
rect 182352 582618 182588 582854
rect 218032 582938 218268 583174
rect 218352 582938 218588 583174
rect 218032 582618 218268 582854
rect 218352 582618 218588 582854
rect 254032 582938 254268 583174
rect 254352 582938 254588 583174
rect 254032 582618 254268 582854
rect 254352 582618 254588 582854
rect 290032 582938 290268 583174
rect 290352 582938 290588 583174
rect 290032 582618 290268 582854
rect 290352 582618 290588 582854
rect 326032 582938 326268 583174
rect 326352 582938 326588 583174
rect 326032 582618 326268 582854
rect 326352 582618 326588 582854
rect 362032 582938 362268 583174
rect 362352 582938 362588 583174
rect 362032 582618 362268 582854
rect 362352 582618 362588 582854
rect 398032 582938 398268 583174
rect 398352 582938 398588 583174
rect 398032 582618 398268 582854
rect 398352 582618 398588 582854
rect 434032 582938 434268 583174
rect 434352 582938 434588 583174
rect 434032 582618 434268 582854
rect 434352 582618 434588 582854
rect 470032 582938 470268 583174
rect 470352 582938 470588 583174
rect 470032 582618 470268 582854
rect 470352 582618 470588 582854
rect 506032 582938 506268 583174
rect 506352 582938 506588 583174
rect 506032 582618 506268 582854
rect 506352 582618 506588 582854
rect 542032 582938 542268 583174
rect 542352 582938 542588 583174
rect 542032 582618 542268 582854
rect 542352 582618 542588 582854
rect 571532 582938 571768 583174
rect 571852 582938 572088 583174
rect 571532 582618 571768 582854
rect 571852 582618 572088 582854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect 9116 579218 9352 579454
rect 9436 579218 9672 579454
rect 9116 578898 9352 579134
rect 9436 578898 9672 579134
rect 56652 579218 56888 579454
rect 56972 579218 57208 579454
rect 56652 578898 56888 579134
rect 56972 578898 57208 579134
rect 92652 579218 92888 579454
rect 92972 579218 93208 579454
rect 92652 578898 92888 579134
rect 92972 578898 93208 579134
rect 128652 579218 128888 579454
rect 128972 579218 129208 579454
rect 128652 578898 128888 579134
rect 128972 578898 129208 579134
rect 164652 579218 164888 579454
rect 164972 579218 165208 579454
rect 164652 578898 164888 579134
rect 164972 578898 165208 579134
rect 200652 579218 200888 579454
rect 200972 579218 201208 579454
rect 200652 578898 200888 579134
rect 200972 578898 201208 579134
rect 236652 579218 236888 579454
rect 236972 579218 237208 579454
rect 236652 578898 236888 579134
rect 236972 578898 237208 579134
rect 272652 579218 272888 579454
rect 272972 579218 273208 579454
rect 272652 578898 272888 579134
rect 272972 578898 273208 579134
rect 308652 579218 308888 579454
rect 308972 579218 309208 579454
rect 308652 578898 308888 579134
rect 308972 578898 309208 579134
rect 344652 579218 344888 579454
rect 344972 579218 345208 579454
rect 344652 578898 344888 579134
rect 344972 578898 345208 579134
rect 380652 579218 380888 579454
rect 380972 579218 381208 579454
rect 380652 578898 380888 579134
rect 380972 578898 381208 579134
rect 416652 579218 416888 579454
rect 416972 579218 417208 579454
rect 416652 578898 416888 579134
rect 416972 578898 417208 579134
rect 452652 579218 452888 579454
rect 452972 579218 453208 579454
rect 452652 578898 452888 579134
rect 452972 578898 453208 579134
rect 488652 579218 488888 579454
rect 488972 579218 489208 579454
rect 488652 578898 488888 579134
rect 488972 578898 489208 579134
rect 524652 579218 524888 579454
rect 524972 579218 525208 579454
rect 524652 578898 524888 579134
rect 524972 578898 525208 579134
rect 560652 579218 560888 579454
rect 560972 579218 561208 579454
rect 560652 578898 560888 579134
rect 560972 578898 561208 579134
rect 570292 579218 570528 579454
rect 570612 579218 570848 579454
rect 570292 578898 570528 579134
rect 570612 578898 570848 579134
rect 7876 546938 8112 547174
rect 8196 546938 8432 547174
rect 7876 546618 8112 546854
rect 8196 546618 8432 546854
rect 38032 546938 38268 547174
rect 38352 546938 38588 547174
rect 38032 546618 38268 546854
rect 38352 546618 38588 546854
rect 74032 546938 74268 547174
rect 74352 546938 74588 547174
rect 74032 546618 74268 546854
rect 74352 546618 74588 546854
rect 110032 546938 110268 547174
rect 110352 546938 110588 547174
rect 110032 546618 110268 546854
rect 110352 546618 110588 546854
rect 146032 546938 146268 547174
rect 146352 546938 146588 547174
rect 146032 546618 146268 546854
rect 146352 546618 146588 546854
rect 182032 546938 182268 547174
rect 182352 546938 182588 547174
rect 182032 546618 182268 546854
rect 182352 546618 182588 546854
rect 218032 546938 218268 547174
rect 218352 546938 218588 547174
rect 218032 546618 218268 546854
rect 218352 546618 218588 546854
rect 254032 546938 254268 547174
rect 254352 546938 254588 547174
rect 254032 546618 254268 546854
rect 254352 546618 254588 546854
rect 290032 546938 290268 547174
rect 290352 546938 290588 547174
rect 290032 546618 290268 546854
rect 290352 546618 290588 546854
rect 326032 546938 326268 547174
rect 326352 546938 326588 547174
rect 326032 546618 326268 546854
rect 326352 546618 326588 546854
rect 362032 546938 362268 547174
rect 362352 546938 362588 547174
rect 362032 546618 362268 546854
rect 362352 546618 362588 546854
rect 398032 546938 398268 547174
rect 398352 546938 398588 547174
rect 398032 546618 398268 546854
rect 398352 546618 398588 546854
rect 434032 546938 434268 547174
rect 434352 546938 434588 547174
rect 434032 546618 434268 546854
rect 434352 546618 434588 546854
rect 470032 546938 470268 547174
rect 470352 546938 470588 547174
rect 470032 546618 470268 546854
rect 470352 546618 470588 546854
rect 506032 546938 506268 547174
rect 506352 546938 506588 547174
rect 506032 546618 506268 546854
rect 506352 546618 506588 546854
rect 542032 546938 542268 547174
rect 542352 546938 542588 547174
rect 542032 546618 542268 546854
rect 542352 546618 542588 546854
rect 571532 546938 571768 547174
rect 571852 546938 572088 547174
rect 571532 546618 571768 546854
rect 571852 546618 572088 546854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect 9116 543218 9352 543454
rect 9436 543218 9672 543454
rect 9116 542898 9352 543134
rect 9436 542898 9672 543134
rect 56652 543218 56888 543454
rect 56972 543218 57208 543454
rect 56652 542898 56888 543134
rect 56972 542898 57208 543134
rect 92652 543218 92888 543454
rect 92972 543218 93208 543454
rect 92652 542898 92888 543134
rect 92972 542898 93208 543134
rect 128652 543218 128888 543454
rect 128972 543218 129208 543454
rect 128652 542898 128888 543134
rect 128972 542898 129208 543134
rect 164652 543218 164888 543454
rect 164972 543218 165208 543454
rect 164652 542898 164888 543134
rect 164972 542898 165208 543134
rect 200652 543218 200888 543454
rect 200972 543218 201208 543454
rect 200652 542898 200888 543134
rect 200972 542898 201208 543134
rect 236652 543218 236888 543454
rect 236972 543218 237208 543454
rect 236652 542898 236888 543134
rect 236972 542898 237208 543134
rect 272652 543218 272888 543454
rect 272972 543218 273208 543454
rect 272652 542898 272888 543134
rect 272972 542898 273208 543134
rect 308652 543218 308888 543454
rect 308972 543218 309208 543454
rect 308652 542898 308888 543134
rect 308972 542898 309208 543134
rect 344652 543218 344888 543454
rect 344972 543218 345208 543454
rect 344652 542898 344888 543134
rect 344972 542898 345208 543134
rect 380652 543218 380888 543454
rect 380972 543218 381208 543454
rect 380652 542898 380888 543134
rect 380972 542898 381208 543134
rect 416652 543218 416888 543454
rect 416972 543218 417208 543454
rect 416652 542898 416888 543134
rect 416972 542898 417208 543134
rect 452652 543218 452888 543454
rect 452972 543218 453208 543454
rect 452652 542898 452888 543134
rect 452972 542898 453208 543134
rect 488652 543218 488888 543454
rect 488972 543218 489208 543454
rect 488652 542898 488888 543134
rect 488972 542898 489208 543134
rect 524652 543218 524888 543454
rect 524972 543218 525208 543454
rect 524652 542898 524888 543134
rect 524972 542898 525208 543134
rect 560652 543218 560888 543454
rect 560972 543218 561208 543454
rect 560652 542898 560888 543134
rect 560972 542898 561208 543134
rect 570292 543218 570528 543454
rect 570612 543218 570848 543454
rect 570292 542898 570528 543134
rect 570612 542898 570848 543134
rect 7876 510938 8112 511174
rect 8196 510938 8432 511174
rect 7876 510618 8112 510854
rect 8196 510618 8432 510854
rect 38032 510938 38268 511174
rect 38352 510938 38588 511174
rect 38032 510618 38268 510854
rect 38352 510618 38588 510854
rect 60622 510938 60858 511174
rect 60622 510618 60858 510854
rect 159098 510938 159334 511174
rect 159098 510618 159334 510854
rect 182032 510938 182268 511174
rect 182352 510938 182588 511174
rect 182032 510618 182268 510854
rect 182352 510618 182588 510854
rect 185622 510938 185858 511174
rect 185622 510618 185858 510854
rect 284098 510938 284334 511174
rect 284098 510618 284334 510854
rect 290032 510938 290268 511174
rect 290352 510938 290588 511174
rect 290032 510618 290268 510854
rect 290352 510618 290588 510854
rect 310622 510938 310858 511174
rect 310622 510618 310858 510854
rect 409098 510938 409334 511174
rect 409098 510618 409334 510854
rect 434032 510938 434268 511174
rect 434352 510938 434588 511174
rect 434032 510618 434268 510854
rect 434352 510618 434588 510854
rect 436622 510938 436858 511174
rect 436622 510618 436858 510854
rect 535098 510938 535334 511174
rect 535098 510618 535334 510854
rect 542032 510938 542268 511174
rect 542352 510938 542588 511174
rect 542032 510618 542268 510854
rect 542352 510618 542588 510854
rect 571532 510938 571768 511174
rect 571852 510938 572088 511174
rect 571532 510618 571768 510854
rect 571852 510618 572088 510854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect 9116 507218 9352 507454
rect 9436 507218 9672 507454
rect 9116 506898 9352 507134
rect 9436 506898 9672 507134
rect 56652 507218 56888 507454
rect 56972 507218 57208 507454
rect 56652 506898 56888 507134
rect 56972 506898 57208 507134
rect 61342 507218 61578 507454
rect 61342 506898 61578 507134
rect 158378 507218 158614 507454
rect 158378 506898 158614 507134
rect 164652 507218 164888 507454
rect 164972 507218 165208 507454
rect 164652 506898 164888 507134
rect 164972 506898 165208 507134
rect 186342 507218 186578 507454
rect 186342 506898 186578 507134
rect 283378 507218 283614 507454
rect 283378 506898 283614 507134
rect 308652 507218 308888 507454
rect 308972 507218 309208 507454
rect 308652 506898 308888 507134
rect 308972 506898 309208 507134
rect 311342 507218 311578 507454
rect 311342 506898 311578 507134
rect 408378 507218 408614 507454
rect 408378 506898 408614 507134
rect 416652 507218 416888 507454
rect 416972 507218 417208 507454
rect 416652 506898 416888 507134
rect 416972 506898 417208 507134
rect 437342 507218 437578 507454
rect 437342 506898 437578 507134
rect 534378 507218 534614 507454
rect 534378 506898 534614 507134
rect 560652 507218 560888 507454
rect 560972 507218 561208 507454
rect 560652 506898 560888 507134
rect 560972 506898 561208 507134
rect 570292 507218 570528 507454
rect 570612 507218 570848 507454
rect 570292 506898 570528 507134
rect 570612 506898 570848 507134
rect 7876 474938 8112 475174
rect 8196 474938 8432 475174
rect 7876 474618 8112 474854
rect 8196 474618 8432 474854
rect 38032 474938 38268 475174
rect 38352 474938 38588 475174
rect 38032 474618 38268 474854
rect 38352 474618 38588 474854
rect 60622 474938 60858 475174
rect 60622 474618 60858 474854
rect 159098 474938 159334 475174
rect 159098 474618 159334 474854
rect 182032 474938 182268 475174
rect 182352 474938 182588 475174
rect 182032 474618 182268 474854
rect 182352 474618 182588 474854
rect 185622 474938 185858 475174
rect 185622 474618 185858 474854
rect 284098 474938 284334 475174
rect 284098 474618 284334 474854
rect 290032 474938 290268 475174
rect 290352 474938 290588 475174
rect 290032 474618 290268 474854
rect 290352 474618 290588 474854
rect 310622 474938 310858 475174
rect 310622 474618 310858 474854
rect 409098 474938 409334 475174
rect 409098 474618 409334 474854
rect 434032 474938 434268 475174
rect 434352 474938 434588 475174
rect 434032 474618 434268 474854
rect 434352 474618 434588 474854
rect 436622 474938 436858 475174
rect 436622 474618 436858 474854
rect 535098 474938 535334 475174
rect 535098 474618 535334 474854
rect 542032 474938 542268 475174
rect 542352 474938 542588 475174
rect 542032 474618 542268 474854
rect 542352 474618 542588 474854
rect 571532 474938 571768 475174
rect 571852 474938 572088 475174
rect 571532 474618 571768 474854
rect 571852 474618 572088 474854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect 9116 471218 9352 471454
rect 9436 471218 9672 471454
rect 9116 470898 9352 471134
rect 9436 470898 9672 471134
rect 56652 471218 56888 471454
rect 56972 471218 57208 471454
rect 56652 470898 56888 471134
rect 56972 470898 57208 471134
rect 61342 471218 61578 471454
rect 61342 470898 61578 471134
rect 158378 471218 158614 471454
rect 158378 470898 158614 471134
rect 164652 471218 164888 471454
rect 164972 471218 165208 471454
rect 164652 470898 164888 471134
rect 164972 470898 165208 471134
rect 186342 471218 186578 471454
rect 186342 470898 186578 471134
rect 283378 471218 283614 471454
rect 283378 470898 283614 471134
rect 308652 471218 308888 471454
rect 308972 471218 309208 471454
rect 308652 470898 308888 471134
rect 308972 470898 309208 471134
rect 311342 471218 311578 471454
rect 311342 470898 311578 471134
rect 408378 471218 408614 471454
rect 408378 470898 408614 471134
rect 416652 471218 416888 471454
rect 416972 471218 417208 471454
rect 416652 470898 416888 471134
rect 416972 470898 417208 471134
rect 437342 471218 437578 471454
rect 437342 470898 437578 471134
rect 534378 471218 534614 471454
rect 534378 470898 534614 471134
rect 560652 471218 560888 471454
rect 560972 471218 561208 471454
rect 560652 470898 560888 471134
rect 560972 470898 561208 471134
rect 570292 471218 570528 471454
rect 570612 471218 570848 471454
rect 570292 470898 570528 471134
rect 570612 470898 570848 471134
rect 7876 438938 8112 439174
rect 8196 438938 8432 439174
rect 7876 438618 8112 438854
rect 8196 438618 8432 438854
rect 38032 438938 38268 439174
rect 38352 438938 38588 439174
rect 38032 438618 38268 438854
rect 38352 438618 38588 438854
rect 60622 438938 60858 439174
rect 60622 438618 60858 438854
rect 159098 438938 159334 439174
rect 159098 438618 159334 438854
rect 182032 438938 182268 439174
rect 182352 438938 182588 439174
rect 182032 438618 182268 438854
rect 182352 438618 182588 438854
rect 185622 438938 185858 439174
rect 185622 438618 185858 438854
rect 284098 438938 284334 439174
rect 284098 438618 284334 438854
rect 290032 438938 290268 439174
rect 290352 438938 290588 439174
rect 290032 438618 290268 438854
rect 290352 438618 290588 438854
rect 310622 438938 310858 439174
rect 310622 438618 310858 438854
rect 409098 438938 409334 439174
rect 409098 438618 409334 438854
rect 434032 438938 434268 439174
rect 434352 438938 434588 439174
rect 434032 438618 434268 438854
rect 434352 438618 434588 438854
rect 436622 438938 436858 439174
rect 436622 438618 436858 438854
rect 535098 438938 535334 439174
rect 535098 438618 535334 438854
rect 542032 438938 542268 439174
rect 542352 438938 542588 439174
rect 542032 438618 542268 438854
rect 542352 438618 542588 438854
rect 571532 438938 571768 439174
rect 571852 438938 572088 439174
rect 571532 438618 571768 438854
rect 571852 438618 572088 438854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect 9116 435218 9352 435454
rect 9436 435218 9672 435454
rect 9116 434898 9352 435134
rect 9436 434898 9672 435134
rect 56652 435218 56888 435454
rect 56972 435218 57208 435454
rect 56652 434898 56888 435134
rect 56972 434898 57208 435134
rect 61342 435218 61578 435454
rect 61342 434898 61578 435134
rect 158378 435218 158614 435454
rect 158378 434898 158614 435134
rect 164652 435218 164888 435454
rect 164972 435218 165208 435454
rect 164652 434898 164888 435134
rect 164972 434898 165208 435134
rect 186342 435218 186578 435454
rect 186342 434898 186578 435134
rect 283378 435218 283614 435454
rect 283378 434898 283614 435134
rect 308652 435218 308888 435454
rect 308972 435218 309208 435454
rect 308652 434898 308888 435134
rect 308972 434898 309208 435134
rect 311342 435218 311578 435454
rect 311342 434898 311578 435134
rect 408378 435218 408614 435454
rect 408378 434898 408614 435134
rect 416652 435218 416888 435454
rect 416972 435218 417208 435454
rect 416652 434898 416888 435134
rect 416972 434898 417208 435134
rect 437342 435218 437578 435454
rect 437342 434898 437578 435134
rect 534378 435218 534614 435454
rect 534378 434898 534614 435134
rect 560652 435218 560888 435454
rect 560972 435218 561208 435454
rect 560652 434898 560888 435134
rect 560972 434898 561208 435134
rect 570292 435218 570528 435454
rect 570612 435218 570848 435454
rect 570292 434898 570528 435134
rect 570612 434898 570848 435134
rect 61342 433008 61578 433244
rect 63008 433008 63244 433244
rect 281712 433008 281948 433244
rect 283378 433008 283614 433244
rect 311342 433008 311578 433244
rect 313008 433008 313244 433244
rect 532712 433008 532948 433244
rect 534378 433008 534614 433244
rect 157392 432328 157628 432564
rect 159098 432328 159334 432564
rect 185622 432328 185858 432564
rect 187328 432328 187564 432564
rect 407392 432328 407628 432564
rect 409098 432328 409334 432564
rect 436622 432328 436858 432564
rect 438328 432328 438564 432564
rect 7876 402938 8112 403174
rect 8196 402938 8432 403174
rect 7876 402618 8112 402854
rect 8196 402618 8432 402854
rect 38032 402938 38268 403174
rect 38352 402938 38588 403174
rect 38032 402618 38268 402854
rect 38352 402618 38588 402854
rect 74032 402938 74268 403174
rect 74352 402938 74588 403174
rect 74032 402618 74268 402854
rect 74352 402618 74588 402854
rect 110032 402938 110268 403174
rect 110352 402938 110588 403174
rect 110032 402618 110268 402854
rect 110352 402618 110588 402854
rect 146032 402938 146268 403174
rect 146352 402938 146588 403174
rect 146032 402618 146268 402854
rect 146352 402618 146588 402854
rect 182032 402938 182268 403174
rect 182352 402938 182588 403174
rect 182032 402618 182268 402854
rect 182352 402618 182588 402854
rect 218032 402938 218268 403174
rect 218352 402938 218588 403174
rect 218032 402618 218268 402854
rect 218352 402618 218588 402854
rect 254032 402938 254268 403174
rect 254352 402938 254588 403174
rect 254032 402618 254268 402854
rect 254352 402618 254588 402854
rect 290032 402938 290268 403174
rect 290352 402938 290588 403174
rect 290032 402618 290268 402854
rect 290352 402618 290588 402854
rect 326032 402938 326268 403174
rect 326352 402938 326588 403174
rect 326032 402618 326268 402854
rect 326352 402618 326588 402854
rect 362032 402938 362268 403174
rect 362352 402938 362588 403174
rect 362032 402618 362268 402854
rect 362352 402618 362588 402854
rect 398032 402938 398268 403174
rect 398352 402938 398588 403174
rect 398032 402618 398268 402854
rect 398352 402618 398588 402854
rect 434032 402938 434268 403174
rect 434352 402938 434588 403174
rect 434032 402618 434268 402854
rect 434352 402618 434588 402854
rect 470032 402938 470268 403174
rect 470352 402938 470588 403174
rect 470032 402618 470268 402854
rect 470352 402618 470588 402854
rect 506032 402938 506268 403174
rect 506352 402938 506588 403174
rect 506032 402618 506268 402854
rect 506352 402618 506588 402854
rect 542032 402938 542268 403174
rect 542352 402938 542588 403174
rect 542032 402618 542268 402854
rect 542352 402618 542588 402854
rect 571532 402938 571768 403174
rect 571852 402938 572088 403174
rect 571532 402618 571768 402854
rect 571852 402618 572088 402854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect 9116 399218 9352 399454
rect 9436 399218 9672 399454
rect 9116 398898 9352 399134
rect 9436 398898 9672 399134
rect 56652 399218 56888 399454
rect 56972 399218 57208 399454
rect 56652 398898 56888 399134
rect 56972 398898 57208 399134
rect 92652 399218 92888 399454
rect 92972 399218 93208 399454
rect 92652 398898 92888 399134
rect 92972 398898 93208 399134
rect 128652 399218 128888 399454
rect 128972 399218 129208 399454
rect 128652 398898 128888 399134
rect 128972 398898 129208 399134
rect 164652 399218 164888 399454
rect 164972 399218 165208 399454
rect 164652 398898 164888 399134
rect 164972 398898 165208 399134
rect 200652 399218 200888 399454
rect 200972 399218 201208 399454
rect 200652 398898 200888 399134
rect 200972 398898 201208 399134
rect 236652 399218 236888 399454
rect 236972 399218 237208 399454
rect 236652 398898 236888 399134
rect 236972 398898 237208 399134
rect 272652 399218 272888 399454
rect 272972 399218 273208 399454
rect 272652 398898 272888 399134
rect 272972 398898 273208 399134
rect 308652 399218 308888 399454
rect 308972 399218 309208 399454
rect 308652 398898 308888 399134
rect 308972 398898 309208 399134
rect 344652 399218 344888 399454
rect 344972 399218 345208 399454
rect 344652 398898 344888 399134
rect 344972 398898 345208 399134
rect 380652 399218 380888 399454
rect 380972 399218 381208 399454
rect 380652 398898 380888 399134
rect 380972 398898 381208 399134
rect 416652 399218 416888 399454
rect 416972 399218 417208 399454
rect 416652 398898 416888 399134
rect 416972 398898 417208 399134
rect 452652 399218 452888 399454
rect 452972 399218 453208 399454
rect 452652 398898 452888 399134
rect 452972 398898 453208 399134
rect 488652 399218 488888 399454
rect 488972 399218 489208 399454
rect 488652 398898 488888 399134
rect 488972 398898 489208 399134
rect 524652 399218 524888 399454
rect 524972 399218 525208 399454
rect 524652 398898 524888 399134
rect 524972 398898 525208 399134
rect 560652 399218 560888 399454
rect 560972 399218 561208 399454
rect 560652 398898 560888 399134
rect 560972 398898 561208 399134
rect 570292 399218 570528 399454
rect 570612 399218 570848 399454
rect 570292 398898 570528 399134
rect 570612 398898 570848 399134
rect 7876 366938 8112 367174
rect 8196 366938 8432 367174
rect 7876 366618 8112 366854
rect 8196 366618 8432 366854
rect 38032 366938 38268 367174
rect 38352 366938 38588 367174
rect 38032 366618 38268 366854
rect 38352 366618 38588 366854
rect 74032 366938 74268 367174
rect 74352 366938 74588 367174
rect 74032 366618 74268 366854
rect 74352 366618 74588 366854
rect 110032 366938 110268 367174
rect 110352 366938 110588 367174
rect 110032 366618 110268 366854
rect 110352 366618 110588 366854
rect 146032 366938 146268 367174
rect 146352 366938 146588 367174
rect 146032 366618 146268 366854
rect 146352 366618 146588 366854
rect 182032 366938 182268 367174
rect 182352 366938 182588 367174
rect 182032 366618 182268 366854
rect 182352 366618 182588 366854
rect 218032 366938 218268 367174
rect 218352 366938 218588 367174
rect 218032 366618 218268 366854
rect 218352 366618 218588 366854
rect 254032 366938 254268 367174
rect 254352 366938 254588 367174
rect 254032 366618 254268 366854
rect 254352 366618 254588 366854
rect 290032 366938 290268 367174
rect 290352 366938 290588 367174
rect 290032 366618 290268 366854
rect 290352 366618 290588 366854
rect 326032 366938 326268 367174
rect 326352 366938 326588 367174
rect 326032 366618 326268 366854
rect 326352 366618 326588 366854
rect 362032 366938 362268 367174
rect 362352 366938 362588 367174
rect 362032 366618 362268 366854
rect 362352 366618 362588 366854
rect 398032 366938 398268 367174
rect 398352 366938 398588 367174
rect 398032 366618 398268 366854
rect 398352 366618 398588 366854
rect 434032 366938 434268 367174
rect 434352 366938 434588 367174
rect 434032 366618 434268 366854
rect 434352 366618 434588 366854
rect 470032 366938 470268 367174
rect 470352 366938 470588 367174
rect 470032 366618 470268 366854
rect 470352 366618 470588 366854
rect 506032 366938 506268 367174
rect 506352 366938 506588 367174
rect 506032 366618 506268 366854
rect 506352 366618 506588 366854
rect 542032 366938 542268 367174
rect 542352 366938 542588 367174
rect 542032 366618 542268 366854
rect 542352 366618 542588 366854
rect 571532 366938 571768 367174
rect 571852 366938 572088 367174
rect 571532 366618 571768 366854
rect 571852 366618 572088 366854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect 9116 363218 9352 363454
rect 9436 363218 9672 363454
rect 9116 362898 9352 363134
rect 9436 362898 9672 363134
rect 56652 363218 56888 363454
rect 56972 363218 57208 363454
rect 56652 362898 56888 363134
rect 56972 362898 57208 363134
rect 92652 363218 92888 363454
rect 92972 363218 93208 363454
rect 92652 362898 92888 363134
rect 92972 362898 93208 363134
rect 128652 363218 128888 363454
rect 128972 363218 129208 363454
rect 128652 362898 128888 363134
rect 128972 362898 129208 363134
rect 164652 363218 164888 363454
rect 164972 363218 165208 363454
rect 164652 362898 164888 363134
rect 164972 362898 165208 363134
rect 200652 363218 200888 363454
rect 200972 363218 201208 363454
rect 200652 362898 200888 363134
rect 200972 362898 201208 363134
rect 236652 363218 236888 363454
rect 236972 363218 237208 363454
rect 236652 362898 236888 363134
rect 236972 362898 237208 363134
rect 272652 363218 272888 363454
rect 272972 363218 273208 363454
rect 272652 362898 272888 363134
rect 272972 362898 273208 363134
rect 308652 363218 308888 363454
rect 308972 363218 309208 363454
rect 308652 362898 308888 363134
rect 308972 362898 309208 363134
rect 344652 363218 344888 363454
rect 344972 363218 345208 363454
rect 344652 362898 344888 363134
rect 344972 362898 345208 363134
rect 380652 363218 380888 363454
rect 380972 363218 381208 363454
rect 380652 362898 380888 363134
rect 380972 362898 381208 363134
rect 416652 363218 416888 363454
rect 416972 363218 417208 363454
rect 416652 362898 416888 363134
rect 416972 362898 417208 363134
rect 452652 363218 452888 363454
rect 452972 363218 453208 363454
rect 452652 362898 452888 363134
rect 452972 362898 453208 363134
rect 488652 363218 488888 363454
rect 488972 363218 489208 363454
rect 488652 362898 488888 363134
rect 488972 362898 489208 363134
rect 524652 363218 524888 363454
rect 524972 363218 525208 363454
rect 524652 362898 524888 363134
rect 524972 362898 525208 363134
rect 560652 363218 560888 363454
rect 560972 363218 561208 363454
rect 560652 362898 560888 363134
rect 560972 362898 561208 363134
rect 570292 363218 570528 363454
rect 570612 363218 570848 363454
rect 570292 362898 570528 363134
rect 570612 362898 570848 363134
rect 7876 330938 8112 331174
rect 8196 330938 8432 331174
rect 7876 330618 8112 330854
rect 8196 330618 8432 330854
rect 38032 330938 38268 331174
rect 38352 330938 38588 331174
rect 38032 330618 38268 330854
rect 38352 330618 38588 330854
rect 74032 330938 74268 331174
rect 74352 330938 74588 331174
rect 74032 330618 74268 330854
rect 74352 330618 74588 330854
rect 110032 330938 110268 331174
rect 110352 330938 110588 331174
rect 110032 330618 110268 330854
rect 110352 330618 110588 330854
rect 146032 330938 146268 331174
rect 146352 330938 146588 331174
rect 146032 330618 146268 330854
rect 146352 330618 146588 330854
rect 182032 330938 182268 331174
rect 182352 330938 182588 331174
rect 182032 330618 182268 330854
rect 182352 330618 182588 330854
rect 218032 330938 218268 331174
rect 218352 330938 218588 331174
rect 218032 330618 218268 330854
rect 218352 330618 218588 330854
rect 254032 330938 254268 331174
rect 254352 330938 254588 331174
rect 254032 330618 254268 330854
rect 254352 330618 254588 330854
rect 290032 330938 290268 331174
rect 290352 330938 290588 331174
rect 290032 330618 290268 330854
rect 290352 330618 290588 330854
rect 326032 330938 326268 331174
rect 326352 330938 326588 331174
rect 326032 330618 326268 330854
rect 326352 330618 326588 330854
rect 362032 330938 362268 331174
rect 362352 330938 362588 331174
rect 362032 330618 362268 330854
rect 362352 330618 362588 330854
rect 398032 330938 398268 331174
rect 398352 330938 398588 331174
rect 398032 330618 398268 330854
rect 398352 330618 398588 330854
rect 434032 330938 434268 331174
rect 434352 330938 434588 331174
rect 434032 330618 434268 330854
rect 434352 330618 434588 330854
rect 470032 330938 470268 331174
rect 470352 330938 470588 331174
rect 470032 330618 470268 330854
rect 470352 330618 470588 330854
rect 506032 330938 506268 331174
rect 506352 330938 506588 331174
rect 506032 330618 506268 330854
rect 506352 330618 506588 330854
rect 542032 330938 542268 331174
rect 542352 330938 542588 331174
rect 542032 330618 542268 330854
rect 542352 330618 542588 330854
rect 571532 330938 571768 331174
rect 571852 330938 572088 331174
rect 571532 330618 571768 330854
rect 571852 330618 572088 330854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect 9116 327218 9352 327454
rect 9436 327218 9672 327454
rect 9116 326898 9352 327134
rect 9436 326898 9672 327134
rect 56652 327218 56888 327454
rect 56972 327218 57208 327454
rect 56652 326898 56888 327134
rect 56972 326898 57208 327134
rect 92652 327218 92888 327454
rect 92972 327218 93208 327454
rect 92652 326898 92888 327134
rect 92972 326898 93208 327134
rect 128652 327218 128888 327454
rect 128972 327218 129208 327454
rect 128652 326898 128888 327134
rect 128972 326898 129208 327134
rect 164652 327218 164888 327454
rect 164972 327218 165208 327454
rect 164652 326898 164888 327134
rect 164972 326898 165208 327134
rect 200652 327218 200888 327454
rect 200972 327218 201208 327454
rect 200652 326898 200888 327134
rect 200972 326898 201208 327134
rect 236652 327218 236888 327454
rect 236972 327218 237208 327454
rect 236652 326898 236888 327134
rect 236972 326898 237208 327134
rect 272652 327218 272888 327454
rect 272972 327218 273208 327454
rect 272652 326898 272888 327134
rect 272972 326898 273208 327134
rect 308652 327218 308888 327454
rect 308972 327218 309208 327454
rect 308652 326898 308888 327134
rect 308972 326898 309208 327134
rect 344652 327218 344888 327454
rect 344972 327218 345208 327454
rect 344652 326898 344888 327134
rect 344972 326898 345208 327134
rect 380652 327218 380888 327454
rect 380972 327218 381208 327454
rect 380652 326898 380888 327134
rect 380972 326898 381208 327134
rect 416652 327218 416888 327454
rect 416972 327218 417208 327454
rect 416652 326898 416888 327134
rect 416972 326898 417208 327134
rect 452652 327218 452888 327454
rect 452972 327218 453208 327454
rect 452652 326898 452888 327134
rect 452972 326898 453208 327134
rect 488652 327218 488888 327454
rect 488972 327218 489208 327454
rect 488652 326898 488888 327134
rect 488972 326898 489208 327134
rect 524652 327218 524888 327454
rect 524972 327218 525208 327454
rect 524652 326898 524888 327134
rect 524972 326898 525208 327134
rect 560652 327218 560888 327454
rect 560972 327218 561208 327454
rect 560652 326898 560888 327134
rect 560972 326898 561208 327134
rect 570292 327218 570528 327454
rect 570612 327218 570848 327454
rect 570292 326898 570528 327134
rect 570612 326898 570848 327134
rect 7876 294938 8112 295174
rect 8196 294938 8432 295174
rect 7876 294618 8112 294854
rect 8196 294618 8432 294854
rect 38032 294938 38268 295174
rect 38352 294938 38588 295174
rect 38032 294618 38268 294854
rect 38352 294618 38588 294854
rect 74032 294938 74268 295174
rect 74352 294938 74588 295174
rect 74032 294618 74268 294854
rect 74352 294618 74588 294854
rect 110032 294938 110268 295174
rect 110352 294938 110588 295174
rect 110032 294618 110268 294854
rect 110352 294618 110588 294854
rect 146032 294938 146268 295174
rect 146352 294938 146588 295174
rect 146032 294618 146268 294854
rect 146352 294618 146588 294854
rect 182032 294938 182268 295174
rect 182352 294938 182588 295174
rect 182032 294618 182268 294854
rect 182352 294618 182588 294854
rect 218032 294938 218268 295174
rect 218352 294938 218588 295174
rect 218032 294618 218268 294854
rect 218352 294618 218588 294854
rect 254032 294938 254268 295174
rect 254352 294938 254588 295174
rect 254032 294618 254268 294854
rect 254352 294618 254588 294854
rect 290032 294938 290268 295174
rect 290352 294938 290588 295174
rect 290032 294618 290268 294854
rect 290352 294618 290588 294854
rect 326032 294938 326268 295174
rect 326352 294938 326588 295174
rect 326032 294618 326268 294854
rect 326352 294618 326588 294854
rect 362032 294938 362268 295174
rect 362352 294938 362588 295174
rect 362032 294618 362268 294854
rect 362352 294618 362588 294854
rect 398032 294938 398268 295174
rect 398352 294938 398588 295174
rect 398032 294618 398268 294854
rect 398352 294618 398588 294854
rect 434032 294938 434268 295174
rect 434352 294938 434588 295174
rect 434032 294618 434268 294854
rect 434352 294618 434588 294854
rect 470032 294938 470268 295174
rect 470352 294938 470588 295174
rect 470032 294618 470268 294854
rect 470352 294618 470588 294854
rect 506032 294938 506268 295174
rect 506352 294938 506588 295174
rect 506032 294618 506268 294854
rect 506352 294618 506588 294854
rect 542032 294938 542268 295174
rect 542352 294938 542588 295174
rect 542032 294618 542268 294854
rect 542352 294618 542588 294854
rect 571532 294938 571768 295174
rect 571852 294938 572088 295174
rect 571532 294618 571768 294854
rect 571852 294618 572088 294854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect 9116 291218 9352 291454
rect 9436 291218 9672 291454
rect 9116 290898 9352 291134
rect 9436 290898 9672 291134
rect 56652 291218 56888 291454
rect 56972 291218 57208 291454
rect 56652 290898 56888 291134
rect 56972 290898 57208 291134
rect 92652 291218 92888 291454
rect 92972 291218 93208 291454
rect 92652 290898 92888 291134
rect 92972 290898 93208 291134
rect 128652 291218 128888 291454
rect 128972 291218 129208 291454
rect 128652 290898 128888 291134
rect 128972 290898 129208 291134
rect 164652 291218 164888 291454
rect 164972 291218 165208 291454
rect 164652 290898 164888 291134
rect 164972 290898 165208 291134
rect 200652 291218 200888 291454
rect 200972 291218 201208 291454
rect 200652 290898 200888 291134
rect 200972 290898 201208 291134
rect 236652 291218 236888 291454
rect 236972 291218 237208 291454
rect 236652 290898 236888 291134
rect 236972 290898 237208 291134
rect 272652 291218 272888 291454
rect 272972 291218 273208 291454
rect 272652 290898 272888 291134
rect 272972 290898 273208 291134
rect 308652 291218 308888 291454
rect 308972 291218 309208 291454
rect 308652 290898 308888 291134
rect 308972 290898 309208 291134
rect 344652 291218 344888 291454
rect 344972 291218 345208 291454
rect 344652 290898 344888 291134
rect 344972 290898 345208 291134
rect 380652 291218 380888 291454
rect 380972 291218 381208 291454
rect 380652 290898 380888 291134
rect 380972 290898 381208 291134
rect 416652 291218 416888 291454
rect 416972 291218 417208 291454
rect 416652 290898 416888 291134
rect 416972 290898 417208 291134
rect 452652 291218 452888 291454
rect 452972 291218 453208 291454
rect 452652 290898 452888 291134
rect 452972 290898 453208 291134
rect 488652 291218 488888 291454
rect 488972 291218 489208 291454
rect 488652 290898 488888 291134
rect 488972 290898 489208 291134
rect 524652 291218 524888 291454
rect 524972 291218 525208 291454
rect 524652 290898 524888 291134
rect 524972 290898 525208 291134
rect 560652 291218 560888 291454
rect 560972 291218 561208 291454
rect 560652 290898 560888 291134
rect 560972 290898 561208 291134
rect 570292 291218 570528 291454
rect 570612 291218 570848 291454
rect 570292 290898 570528 291134
rect 570612 290898 570848 291134
rect 7876 258938 8112 259174
rect 8196 258938 8432 259174
rect 7876 258618 8112 258854
rect 8196 258618 8432 258854
rect 38032 258938 38268 259174
rect 38352 258938 38588 259174
rect 38032 258618 38268 258854
rect 38352 258618 38588 258854
rect 74032 258938 74268 259174
rect 74352 258938 74588 259174
rect 74032 258618 74268 258854
rect 74352 258618 74588 258854
rect 110032 258938 110268 259174
rect 110352 258938 110588 259174
rect 110032 258618 110268 258854
rect 110352 258618 110588 258854
rect 146032 258938 146268 259174
rect 146352 258938 146588 259174
rect 146032 258618 146268 258854
rect 146352 258618 146588 258854
rect 182032 258938 182268 259174
rect 182352 258938 182588 259174
rect 182032 258618 182268 258854
rect 182352 258618 182588 258854
rect 218032 258938 218268 259174
rect 218352 258938 218588 259174
rect 218032 258618 218268 258854
rect 218352 258618 218588 258854
rect 254032 258938 254268 259174
rect 254352 258938 254588 259174
rect 254032 258618 254268 258854
rect 254352 258618 254588 258854
rect 290032 258938 290268 259174
rect 290352 258938 290588 259174
rect 290032 258618 290268 258854
rect 290352 258618 290588 258854
rect 326032 258938 326268 259174
rect 326352 258938 326588 259174
rect 326032 258618 326268 258854
rect 326352 258618 326588 258854
rect 362032 258938 362268 259174
rect 362352 258938 362588 259174
rect 362032 258618 362268 258854
rect 362352 258618 362588 258854
rect 398032 258938 398268 259174
rect 398352 258938 398588 259174
rect 398032 258618 398268 258854
rect 398352 258618 398588 258854
rect 434032 258938 434268 259174
rect 434352 258938 434588 259174
rect 434032 258618 434268 258854
rect 434352 258618 434588 258854
rect 470032 258938 470268 259174
rect 470352 258938 470588 259174
rect 470032 258618 470268 258854
rect 470352 258618 470588 258854
rect 506032 258938 506268 259174
rect 506352 258938 506588 259174
rect 506032 258618 506268 258854
rect 506352 258618 506588 258854
rect 542032 258938 542268 259174
rect 542352 258938 542588 259174
rect 542032 258618 542268 258854
rect 542352 258618 542588 258854
rect 571532 258938 571768 259174
rect 571852 258938 572088 259174
rect 571532 258618 571768 258854
rect 571852 258618 572088 258854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect 9116 255218 9352 255454
rect 9436 255218 9672 255454
rect 9116 254898 9352 255134
rect 9436 254898 9672 255134
rect 56652 255218 56888 255454
rect 56972 255218 57208 255454
rect 56652 254898 56888 255134
rect 56972 254898 57208 255134
rect 92652 255218 92888 255454
rect 92972 255218 93208 255454
rect 92652 254898 92888 255134
rect 92972 254898 93208 255134
rect 128652 255218 128888 255454
rect 128972 255218 129208 255454
rect 128652 254898 128888 255134
rect 128972 254898 129208 255134
rect 164652 255218 164888 255454
rect 164972 255218 165208 255454
rect 164652 254898 164888 255134
rect 164972 254898 165208 255134
rect 200652 255218 200888 255454
rect 200972 255218 201208 255454
rect 200652 254898 200888 255134
rect 200972 254898 201208 255134
rect 236652 255218 236888 255454
rect 236972 255218 237208 255454
rect 236652 254898 236888 255134
rect 236972 254898 237208 255134
rect 272652 255218 272888 255454
rect 272972 255218 273208 255454
rect 272652 254898 272888 255134
rect 272972 254898 273208 255134
rect 308652 255218 308888 255454
rect 308972 255218 309208 255454
rect 308652 254898 308888 255134
rect 308972 254898 309208 255134
rect 344652 255218 344888 255454
rect 344972 255218 345208 255454
rect 344652 254898 344888 255134
rect 344972 254898 345208 255134
rect 380652 255218 380888 255454
rect 380972 255218 381208 255454
rect 380652 254898 380888 255134
rect 380972 254898 381208 255134
rect 416652 255218 416888 255454
rect 416972 255218 417208 255454
rect 416652 254898 416888 255134
rect 416972 254898 417208 255134
rect 452652 255218 452888 255454
rect 452972 255218 453208 255454
rect 452652 254898 452888 255134
rect 452972 254898 453208 255134
rect 488652 255218 488888 255454
rect 488972 255218 489208 255454
rect 488652 254898 488888 255134
rect 488972 254898 489208 255134
rect 524652 255218 524888 255454
rect 524972 255218 525208 255454
rect 524652 254898 524888 255134
rect 524972 254898 525208 255134
rect 560652 255218 560888 255454
rect 560972 255218 561208 255454
rect 560652 254898 560888 255134
rect 560972 254898 561208 255134
rect 570292 255218 570528 255454
rect 570612 255218 570848 255454
rect 570292 254898 570528 255134
rect 570612 254898 570848 255134
rect 7876 222938 8112 223174
rect 8196 222938 8432 223174
rect 7876 222618 8112 222854
rect 8196 222618 8432 222854
rect 38032 222938 38268 223174
rect 38352 222938 38588 223174
rect 38032 222618 38268 222854
rect 38352 222618 38588 222854
rect 74032 222938 74268 223174
rect 74352 222938 74588 223174
rect 74032 222618 74268 222854
rect 74352 222618 74588 222854
rect 110032 222938 110268 223174
rect 110352 222938 110588 223174
rect 110032 222618 110268 222854
rect 110352 222618 110588 222854
rect 146032 222938 146268 223174
rect 146352 222938 146588 223174
rect 146032 222618 146268 222854
rect 146352 222618 146588 222854
rect 182032 222938 182268 223174
rect 182352 222938 182588 223174
rect 182032 222618 182268 222854
rect 182352 222618 182588 222854
rect 218032 222938 218268 223174
rect 218352 222938 218588 223174
rect 218032 222618 218268 222854
rect 218352 222618 218588 222854
rect 254032 222938 254268 223174
rect 254352 222938 254588 223174
rect 254032 222618 254268 222854
rect 254352 222618 254588 222854
rect 290032 222938 290268 223174
rect 290352 222938 290588 223174
rect 290032 222618 290268 222854
rect 290352 222618 290588 222854
rect 326032 222938 326268 223174
rect 326352 222938 326588 223174
rect 326032 222618 326268 222854
rect 326352 222618 326588 222854
rect 362032 222938 362268 223174
rect 362352 222938 362588 223174
rect 362032 222618 362268 222854
rect 362352 222618 362588 222854
rect 398032 222938 398268 223174
rect 398352 222938 398588 223174
rect 398032 222618 398268 222854
rect 398352 222618 398588 222854
rect 434032 222938 434268 223174
rect 434352 222938 434588 223174
rect 434032 222618 434268 222854
rect 434352 222618 434588 222854
rect 470032 222938 470268 223174
rect 470352 222938 470588 223174
rect 470032 222618 470268 222854
rect 470352 222618 470588 222854
rect 506032 222938 506268 223174
rect 506352 222938 506588 223174
rect 506032 222618 506268 222854
rect 506352 222618 506588 222854
rect 542032 222938 542268 223174
rect 542352 222938 542588 223174
rect 542032 222618 542268 222854
rect 542352 222618 542588 222854
rect 571532 222938 571768 223174
rect 571852 222938 572088 223174
rect 571532 222618 571768 222854
rect 571852 222618 572088 222854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect 9116 219218 9352 219454
rect 9436 219218 9672 219454
rect 9116 218898 9352 219134
rect 9436 218898 9672 219134
rect 56652 219218 56888 219454
rect 56972 219218 57208 219454
rect 56652 218898 56888 219134
rect 56972 218898 57208 219134
rect 92652 219218 92888 219454
rect 92972 219218 93208 219454
rect 92652 218898 92888 219134
rect 92972 218898 93208 219134
rect 128652 219218 128888 219454
rect 128972 219218 129208 219454
rect 128652 218898 128888 219134
rect 128972 218898 129208 219134
rect 164652 219218 164888 219454
rect 164972 219218 165208 219454
rect 164652 218898 164888 219134
rect 164972 218898 165208 219134
rect 200652 219218 200888 219454
rect 200972 219218 201208 219454
rect 200652 218898 200888 219134
rect 200972 218898 201208 219134
rect 236652 219218 236888 219454
rect 236972 219218 237208 219454
rect 236652 218898 236888 219134
rect 236972 218898 237208 219134
rect 272652 219218 272888 219454
rect 272972 219218 273208 219454
rect 272652 218898 272888 219134
rect 272972 218898 273208 219134
rect 308652 219218 308888 219454
rect 308972 219218 309208 219454
rect 308652 218898 308888 219134
rect 308972 218898 309208 219134
rect 344652 219218 344888 219454
rect 344972 219218 345208 219454
rect 344652 218898 344888 219134
rect 344972 218898 345208 219134
rect 380652 219218 380888 219454
rect 380972 219218 381208 219454
rect 380652 218898 380888 219134
rect 380972 218898 381208 219134
rect 416652 219218 416888 219454
rect 416972 219218 417208 219454
rect 416652 218898 416888 219134
rect 416972 218898 417208 219134
rect 452652 219218 452888 219454
rect 452972 219218 453208 219454
rect 452652 218898 452888 219134
rect 452972 218898 453208 219134
rect 488652 219218 488888 219454
rect 488972 219218 489208 219454
rect 488652 218898 488888 219134
rect 488972 218898 489208 219134
rect 524652 219218 524888 219454
rect 524972 219218 525208 219454
rect 524652 218898 524888 219134
rect 524972 218898 525208 219134
rect 560652 219218 560888 219454
rect 560972 219218 561208 219454
rect 560652 218898 560888 219134
rect 560972 218898 561208 219134
rect 570292 219218 570528 219454
rect 570612 219218 570848 219454
rect 570292 218898 570528 219134
rect 570612 218898 570848 219134
rect 7876 186938 8112 187174
rect 8196 186938 8432 187174
rect 7876 186618 8112 186854
rect 8196 186618 8432 186854
rect 38032 186938 38268 187174
rect 38352 186938 38588 187174
rect 38032 186618 38268 186854
rect 38352 186618 38588 186854
rect 60622 186938 60858 187174
rect 60622 186618 60858 186854
rect 159098 186938 159334 187174
rect 159098 186618 159334 186854
rect 182032 186938 182268 187174
rect 182352 186938 182588 187174
rect 182032 186618 182268 186854
rect 182352 186618 182588 186854
rect 185622 186938 185858 187174
rect 185622 186618 185858 186854
rect 284098 186938 284334 187174
rect 284098 186618 284334 186854
rect 290032 186938 290268 187174
rect 290352 186938 290588 187174
rect 290032 186618 290268 186854
rect 290352 186618 290588 186854
rect 310622 186938 310858 187174
rect 310622 186618 310858 186854
rect 409098 186938 409334 187174
rect 409098 186618 409334 186854
rect 434032 186938 434268 187174
rect 434352 186938 434588 187174
rect 434032 186618 434268 186854
rect 434352 186618 434588 186854
rect 436622 186938 436858 187174
rect 436622 186618 436858 186854
rect 535098 186938 535334 187174
rect 535098 186618 535334 186854
rect 542032 186938 542268 187174
rect 542352 186938 542588 187174
rect 542032 186618 542268 186854
rect 542352 186618 542588 186854
rect 571532 186938 571768 187174
rect 571852 186938 572088 187174
rect 571532 186618 571768 186854
rect 571852 186618 572088 186854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect 9116 183218 9352 183454
rect 9436 183218 9672 183454
rect 9116 182898 9352 183134
rect 9436 182898 9672 183134
rect 56652 183218 56888 183454
rect 56972 183218 57208 183454
rect 56652 182898 56888 183134
rect 56972 182898 57208 183134
rect 61342 183218 61578 183454
rect 61342 182898 61578 183134
rect 158378 183218 158614 183454
rect 158378 182898 158614 183134
rect 164652 183218 164888 183454
rect 164972 183218 165208 183454
rect 164652 182898 164888 183134
rect 164972 182898 165208 183134
rect 186342 183218 186578 183454
rect 186342 182898 186578 183134
rect 283378 183218 283614 183454
rect 283378 182898 283614 183134
rect 308652 183218 308888 183454
rect 308972 183218 309208 183454
rect 308652 182898 308888 183134
rect 308972 182898 309208 183134
rect 311342 183218 311578 183454
rect 311342 182898 311578 183134
rect 408378 183218 408614 183454
rect 408378 182898 408614 183134
rect 416652 183218 416888 183454
rect 416972 183218 417208 183454
rect 416652 182898 416888 183134
rect 416972 182898 417208 183134
rect 437342 183218 437578 183454
rect 437342 182898 437578 183134
rect 534378 183218 534614 183454
rect 534378 182898 534614 183134
rect 560652 183218 560888 183454
rect 560972 183218 561208 183454
rect 560652 182898 560888 183134
rect 560972 182898 561208 183134
rect 570292 183218 570528 183454
rect 570612 183218 570848 183454
rect 570292 182898 570528 183134
rect 570612 182898 570848 183134
rect 7876 150938 8112 151174
rect 8196 150938 8432 151174
rect 7876 150618 8112 150854
rect 8196 150618 8432 150854
rect 38032 150938 38268 151174
rect 38352 150938 38588 151174
rect 38032 150618 38268 150854
rect 38352 150618 38588 150854
rect 60622 150938 60858 151174
rect 60622 150618 60858 150854
rect 159098 150938 159334 151174
rect 159098 150618 159334 150854
rect 182032 150938 182268 151174
rect 182352 150938 182588 151174
rect 182032 150618 182268 150854
rect 182352 150618 182588 150854
rect 185622 150938 185858 151174
rect 185622 150618 185858 150854
rect 284098 150938 284334 151174
rect 284098 150618 284334 150854
rect 290032 150938 290268 151174
rect 290352 150938 290588 151174
rect 290032 150618 290268 150854
rect 290352 150618 290588 150854
rect 310622 150938 310858 151174
rect 310622 150618 310858 150854
rect 409098 150938 409334 151174
rect 409098 150618 409334 150854
rect 434032 150938 434268 151174
rect 434352 150938 434588 151174
rect 434032 150618 434268 150854
rect 434352 150618 434588 150854
rect 436622 150938 436858 151174
rect 436622 150618 436858 150854
rect 535098 150938 535334 151174
rect 535098 150618 535334 150854
rect 542032 150938 542268 151174
rect 542352 150938 542588 151174
rect 542032 150618 542268 150854
rect 542352 150618 542588 150854
rect 571532 150938 571768 151174
rect 571852 150938 572088 151174
rect 571532 150618 571768 150854
rect 571852 150618 572088 150854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect 9116 147218 9352 147454
rect 9436 147218 9672 147454
rect 9116 146898 9352 147134
rect 9436 146898 9672 147134
rect 56652 147218 56888 147454
rect 56972 147218 57208 147454
rect 56652 146898 56888 147134
rect 56972 146898 57208 147134
rect 61342 147218 61578 147454
rect 61342 146898 61578 147134
rect 158378 147218 158614 147454
rect 158378 146898 158614 147134
rect 164652 147218 164888 147454
rect 164972 147218 165208 147454
rect 164652 146898 164888 147134
rect 164972 146898 165208 147134
rect 186342 147218 186578 147454
rect 186342 146898 186578 147134
rect 283378 147218 283614 147454
rect 283378 146898 283614 147134
rect 308652 147218 308888 147454
rect 308972 147218 309208 147454
rect 308652 146898 308888 147134
rect 308972 146898 309208 147134
rect 311342 147218 311578 147454
rect 311342 146898 311578 147134
rect 408378 147218 408614 147454
rect 408378 146898 408614 147134
rect 416652 147218 416888 147454
rect 416972 147218 417208 147454
rect 416652 146898 416888 147134
rect 416972 146898 417208 147134
rect 437342 147218 437578 147454
rect 437342 146898 437578 147134
rect 534378 147218 534614 147454
rect 534378 146898 534614 147134
rect 560652 147218 560888 147454
rect 560972 147218 561208 147454
rect 560652 146898 560888 147134
rect 560972 146898 561208 147134
rect 570292 147218 570528 147454
rect 570612 147218 570848 147454
rect 570292 146898 570528 147134
rect 570612 146898 570848 147134
rect 61342 121008 61578 121244
rect 63008 121008 63244 121244
rect 281712 121008 281948 121244
rect 283378 121008 283614 121244
rect 311342 121008 311578 121244
rect 313008 121008 313244 121244
rect 532712 121008 532948 121244
rect 534378 121008 534614 121244
rect 157392 120328 157628 120564
rect 159098 120328 159334 120564
rect 185622 120328 185858 120564
rect 187328 120328 187564 120564
rect 407392 120328 407628 120564
rect 409098 120328 409334 120564
rect 436622 120328 436858 120564
rect 438328 120328 438564 120564
rect 7876 114938 8112 115174
rect 8196 114938 8432 115174
rect 7876 114618 8112 114854
rect 8196 114618 8432 114854
rect 38032 114938 38268 115174
rect 38352 114938 38588 115174
rect 38032 114618 38268 114854
rect 38352 114618 38588 114854
rect 74032 114938 74268 115174
rect 74352 114938 74588 115174
rect 74032 114618 74268 114854
rect 74352 114618 74588 114854
rect 110032 114938 110268 115174
rect 110352 114938 110588 115174
rect 110032 114618 110268 114854
rect 110352 114618 110588 114854
rect 146032 114938 146268 115174
rect 146352 114938 146588 115174
rect 146032 114618 146268 114854
rect 146352 114618 146588 114854
rect 182032 114938 182268 115174
rect 182352 114938 182588 115174
rect 182032 114618 182268 114854
rect 182352 114618 182588 114854
rect 218032 114938 218268 115174
rect 218352 114938 218588 115174
rect 218032 114618 218268 114854
rect 218352 114618 218588 114854
rect 254032 114938 254268 115174
rect 254352 114938 254588 115174
rect 254032 114618 254268 114854
rect 254352 114618 254588 114854
rect 290032 114938 290268 115174
rect 290352 114938 290588 115174
rect 290032 114618 290268 114854
rect 290352 114618 290588 114854
rect 326032 114938 326268 115174
rect 326352 114938 326588 115174
rect 326032 114618 326268 114854
rect 326352 114618 326588 114854
rect 362032 114938 362268 115174
rect 362352 114938 362588 115174
rect 362032 114618 362268 114854
rect 362352 114618 362588 114854
rect 398032 114938 398268 115174
rect 398352 114938 398588 115174
rect 398032 114618 398268 114854
rect 398352 114618 398588 114854
rect 434032 114938 434268 115174
rect 434352 114938 434588 115174
rect 434032 114618 434268 114854
rect 434352 114618 434588 114854
rect 470032 114938 470268 115174
rect 470352 114938 470588 115174
rect 470032 114618 470268 114854
rect 470352 114618 470588 114854
rect 506032 114938 506268 115174
rect 506352 114938 506588 115174
rect 506032 114618 506268 114854
rect 506352 114618 506588 114854
rect 542032 114938 542268 115174
rect 542352 114938 542588 115174
rect 542032 114618 542268 114854
rect 542352 114618 542588 114854
rect 571532 114938 571768 115174
rect 571852 114938 572088 115174
rect 571532 114618 571768 114854
rect 571852 114618 572088 114854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect 9116 111218 9352 111454
rect 9436 111218 9672 111454
rect 9116 110898 9352 111134
rect 9436 110898 9672 111134
rect 56652 111218 56888 111454
rect 56972 111218 57208 111454
rect 56652 110898 56888 111134
rect 56972 110898 57208 111134
rect 92652 111218 92888 111454
rect 92972 111218 93208 111454
rect 92652 110898 92888 111134
rect 92972 110898 93208 111134
rect 128652 111218 128888 111454
rect 128972 111218 129208 111454
rect 128652 110898 128888 111134
rect 128972 110898 129208 111134
rect 164652 111218 164888 111454
rect 164972 111218 165208 111454
rect 164652 110898 164888 111134
rect 164972 110898 165208 111134
rect 200652 111218 200888 111454
rect 200972 111218 201208 111454
rect 200652 110898 200888 111134
rect 200972 110898 201208 111134
rect 236652 111218 236888 111454
rect 236972 111218 237208 111454
rect 236652 110898 236888 111134
rect 236972 110898 237208 111134
rect 272652 111218 272888 111454
rect 272972 111218 273208 111454
rect 272652 110898 272888 111134
rect 272972 110898 273208 111134
rect 308652 111218 308888 111454
rect 308972 111218 309208 111454
rect 308652 110898 308888 111134
rect 308972 110898 309208 111134
rect 344652 111218 344888 111454
rect 344972 111218 345208 111454
rect 344652 110898 344888 111134
rect 344972 110898 345208 111134
rect 380652 111218 380888 111454
rect 380972 111218 381208 111454
rect 380652 110898 380888 111134
rect 380972 110898 381208 111134
rect 416652 111218 416888 111454
rect 416972 111218 417208 111454
rect 416652 110898 416888 111134
rect 416972 110898 417208 111134
rect 452652 111218 452888 111454
rect 452972 111218 453208 111454
rect 452652 110898 452888 111134
rect 452972 110898 453208 111134
rect 488652 111218 488888 111454
rect 488972 111218 489208 111454
rect 488652 110898 488888 111134
rect 488972 110898 489208 111134
rect 524652 111218 524888 111454
rect 524972 111218 525208 111454
rect 524652 110898 524888 111134
rect 524972 110898 525208 111134
rect 560652 111218 560888 111454
rect 560972 111218 561208 111454
rect 560652 110898 560888 111134
rect 560972 110898 561208 111134
rect 570292 111218 570528 111454
rect 570612 111218 570848 111454
rect 570292 110898 570528 111134
rect 570612 110898 570848 111134
rect 7876 78938 8112 79174
rect 8196 78938 8432 79174
rect 7876 78618 8112 78854
rect 8196 78618 8432 78854
rect 38032 78938 38268 79174
rect 38352 78938 38588 79174
rect 38032 78618 38268 78854
rect 38352 78618 38588 78854
rect 60622 78938 60858 79174
rect 60622 78618 60858 78854
rect 159098 78938 159334 79174
rect 159098 78618 159334 78854
rect 182032 78938 182268 79174
rect 182352 78938 182588 79174
rect 182032 78618 182268 78854
rect 182352 78618 182588 78854
rect 185622 78938 185858 79174
rect 185622 78618 185858 78854
rect 284098 78938 284334 79174
rect 284098 78618 284334 78854
rect 290032 78938 290268 79174
rect 290352 78938 290588 79174
rect 290032 78618 290268 78854
rect 290352 78618 290588 78854
rect 310622 78938 310858 79174
rect 310622 78618 310858 78854
rect 409098 78938 409334 79174
rect 409098 78618 409334 78854
rect 434032 78938 434268 79174
rect 434352 78938 434588 79174
rect 434032 78618 434268 78854
rect 434352 78618 434588 78854
rect 436622 78938 436858 79174
rect 436622 78618 436858 78854
rect 535098 78938 535334 79174
rect 535098 78618 535334 78854
rect 542032 78938 542268 79174
rect 542352 78938 542588 79174
rect 542032 78618 542268 78854
rect 542352 78618 542588 78854
rect 571532 78938 571768 79174
rect 571852 78938 572088 79174
rect 571532 78618 571768 78854
rect 571852 78618 572088 78854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect 9116 75218 9352 75454
rect 9436 75218 9672 75454
rect 9116 74898 9352 75134
rect 9436 74898 9672 75134
rect 56652 75218 56888 75454
rect 56972 75218 57208 75454
rect 56652 74898 56888 75134
rect 56972 74898 57208 75134
rect 61342 75218 61578 75454
rect 61342 74898 61578 75134
rect 158378 75218 158614 75454
rect 158378 74898 158614 75134
rect 164652 75218 164888 75454
rect 164972 75218 165208 75454
rect 164652 74898 164888 75134
rect 164972 74898 165208 75134
rect 186342 75218 186578 75454
rect 186342 74898 186578 75134
rect 283378 75218 283614 75454
rect 283378 74898 283614 75134
rect 308652 75218 308888 75454
rect 308972 75218 309208 75454
rect 308652 74898 308888 75134
rect 308972 74898 309208 75134
rect 311342 75218 311578 75454
rect 311342 74898 311578 75134
rect 408378 75218 408614 75454
rect 408378 74898 408614 75134
rect 416652 75218 416888 75454
rect 416972 75218 417208 75454
rect 416652 74898 416888 75134
rect 416972 74898 417208 75134
rect 437342 75218 437578 75454
rect 437342 74898 437578 75134
rect 534378 75218 534614 75454
rect 534378 74898 534614 75134
rect 560652 75218 560888 75454
rect 560972 75218 561208 75454
rect 560652 74898 560888 75134
rect 560972 74898 561208 75134
rect 570292 75218 570528 75454
rect 570612 75218 570848 75454
rect 570292 74898 570528 75134
rect 570612 74898 570848 75134
rect 7876 42938 8112 43174
rect 8196 42938 8432 43174
rect 7876 42618 8112 42854
rect 8196 42618 8432 42854
rect 38032 42938 38268 43174
rect 38352 42938 38588 43174
rect 38032 42618 38268 42854
rect 38352 42618 38588 42854
rect 60622 42938 60858 43174
rect 60622 42618 60858 42854
rect 159098 42938 159334 43174
rect 159098 42618 159334 42854
rect 182032 42938 182268 43174
rect 182352 42938 182588 43174
rect 182032 42618 182268 42854
rect 182352 42618 182588 42854
rect 185622 42938 185858 43174
rect 185622 42618 185858 42854
rect 284098 42938 284334 43174
rect 284098 42618 284334 42854
rect 290032 42938 290268 43174
rect 290352 42938 290588 43174
rect 290032 42618 290268 42854
rect 290352 42618 290588 42854
rect 310622 42938 310858 43174
rect 310622 42618 310858 42854
rect 409098 42938 409334 43174
rect 409098 42618 409334 42854
rect 434032 42938 434268 43174
rect 434352 42938 434588 43174
rect 434032 42618 434268 42854
rect 434352 42618 434588 42854
rect 436622 42938 436858 43174
rect 436622 42618 436858 42854
rect 535098 42938 535334 43174
rect 535098 42618 535334 42854
rect 542032 42938 542268 43174
rect 542352 42938 542588 43174
rect 542032 42618 542268 42854
rect 542352 42618 542588 42854
rect 571532 42938 571768 43174
rect 571852 42938 572088 43174
rect 571532 42618 571768 42854
rect 571852 42618 572088 42854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect 9116 39218 9352 39454
rect 9436 39218 9672 39454
rect 9116 38898 9352 39134
rect 9436 38898 9672 39134
rect 56652 39218 56888 39454
rect 56972 39218 57208 39454
rect 56652 38898 56888 39134
rect 56972 38898 57208 39134
rect 61342 39218 61578 39454
rect 61342 38898 61578 39134
rect 158378 39218 158614 39454
rect 158378 38898 158614 39134
rect 164652 39218 164888 39454
rect 164972 39218 165208 39454
rect 164652 38898 164888 39134
rect 164972 38898 165208 39134
rect 186342 39218 186578 39454
rect 186342 38898 186578 39134
rect 283378 39218 283614 39454
rect 283378 38898 283614 39134
rect 308652 39218 308888 39454
rect 308972 39218 309208 39454
rect 308652 38898 308888 39134
rect 308972 38898 309208 39134
rect 311342 39218 311578 39454
rect 311342 38898 311578 39134
rect 408378 39218 408614 39454
rect 408378 38898 408614 39134
rect 416652 39218 416888 39454
rect 416972 39218 417208 39454
rect 416652 38898 416888 39134
rect 416972 38898 417208 39134
rect 437342 39218 437578 39454
rect 437342 38898 437578 39134
rect 534378 39218 534614 39454
rect 534378 38898 534614 39134
rect 560652 39218 560888 39454
rect 560972 39218 561208 39454
rect 560652 38898 560888 39134
rect 560972 38898 561208 39134
rect 570292 39218 570528 39454
rect 570612 39218 570848 39454
rect 570292 38898 570528 39134
rect 570612 38898 570848 39134
rect 61342 21008 61578 21244
rect 63008 21008 63244 21244
rect 188008 21008 188244 21244
rect 311342 21008 311578 21244
rect 313008 21008 313244 21244
rect 439008 21008 439244 21244
rect 62328 20328 62564 20564
rect 185622 20328 185858 20564
rect 187328 20328 187564 20564
rect 312328 20328 312564 20564
rect 436622 20328 436858 20564
rect 438328 20328 438564 20564
rect 62328 19598 62564 19834
rect 188008 19342 188244 19578
rect 312328 19598 312564 19834
rect 439008 19342 439244 19578
rect 9116 9444 9352 9680
rect 9436 9444 9672 9680
rect 9116 9124 9352 9360
rect 9436 9124 9672 9360
rect 56652 9444 56888 9680
rect 56972 9444 57208 9680
rect 56652 9124 56888 9360
rect 56972 9124 57208 9360
rect 92652 9444 92888 9680
rect 92972 9444 93208 9680
rect 92652 9124 92888 9360
rect 92972 9124 93208 9360
rect 128652 9444 128888 9680
rect 128972 9444 129208 9680
rect 128652 9124 128888 9360
rect 128972 9124 129208 9360
rect 164652 9444 164888 9680
rect 164972 9444 165208 9680
rect 164652 9124 164888 9360
rect 164972 9124 165208 9360
rect 200652 9444 200888 9680
rect 200972 9444 201208 9680
rect 200652 9124 200888 9360
rect 200972 9124 201208 9360
rect 236652 9444 236888 9680
rect 236972 9444 237208 9680
rect 236652 9124 236888 9360
rect 236972 9124 237208 9360
rect 272652 9444 272888 9680
rect 272972 9444 273208 9680
rect 272652 9124 272888 9360
rect 272972 9124 273208 9360
rect 308652 9444 308888 9680
rect 308972 9444 309208 9680
rect 308652 9124 308888 9360
rect 308972 9124 309208 9360
rect 344652 9444 344888 9680
rect 344972 9444 345208 9680
rect 344652 9124 344888 9360
rect 344972 9124 345208 9360
rect 380652 9444 380888 9680
rect 380972 9444 381208 9680
rect 380652 9124 380888 9360
rect 380972 9124 381208 9360
rect 416652 9444 416888 9680
rect 416972 9444 417208 9680
rect 416652 9124 416888 9360
rect 416972 9124 417208 9360
rect 452652 9444 452888 9680
rect 452972 9444 453208 9680
rect 452652 9124 452888 9360
rect 452972 9124 453208 9360
rect 488652 9444 488888 9680
rect 488972 9444 489208 9680
rect 488652 9124 488888 9360
rect 488972 9124 489208 9360
rect 524652 9444 524888 9680
rect 524972 9444 525208 9680
rect 524652 9124 524888 9360
rect 524972 9124 525208 9360
rect 560652 9444 560888 9680
rect 560972 9444 561208 9680
rect 560652 9124 560888 9360
rect 560972 9124 561208 9360
rect 570292 9444 570528 9680
rect 570612 9444 570848 9680
rect 570292 9124 570528 9360
rect 570612 9124 570848 9360
rect 7876 8204 8112 8440
rect 8196 8204 8432 8440
rect 7876 7884 8112 8120
rect 8196 7884 8432 8120
rect 38032 8204 38268 8440
rect 38352 8204 38588 8440
rect 38032 7884 38268 8120
rect 38352 7884 38588 8120
rect 74032 8204 74268 8440
rect 74352 8204 74588 8440
rect 74032 7884 74268 8120
rect 74352 7884 74588 8120
rect 110032 8204 110268 8440
rect 110352 8204 110588 8440
rect 110032 7884 110268 8120
rect 110352 7884 110588 8120
rect 146032 8204 146268 8440
rect 146352 8204 146588 8440
rect 146032 7884 146268 8120
rect 146352 7884 146588 8120
rect 182032 8204 182268 8440
rect 182352 8204 182588 8440
rect 182032 7884 182268 8120
rect 182352 7884 182588 8120
rect 218032 8204 218268 8440
rect 218352 8204 218588 8440
rect 218032 7884 218268 8120
rect 218352 7884 218588 8120
rect 254032 8204 254268 8440
rect 254352 8204 254588 8440
rect 254032 7884 254268 8120
rect 254352 7884 254588 8120
rect 290032 8204 290268 8440
rect 290352 8204 290588 8440
rect 290032 7884 290268 8120
rect 290352 7884 290588 8120
rect 326032 8204 326268 8440
rect 326352 8204 326588 8440
rect 326032 7884 326268 8120
rect 326352 7884 326588 8120
rect 362032 8204 362268 8440
rect 362352 8204 362588 8440
rect 362032 7884 362268 8120
rect 362352 7884 362588 8120
rect 398032 8204 398268 8440
rect 398352 8204 398588 8440
rect 398032 7884 398268 8120
rect 398352 7884 398588 8120
rect 434032 8204 434268 8440
rect 434352 8204 434588 8440
rect 434032 7884 434268 8120
rect 434352 7884 434588 8120
rect 470032 8204 470268 8440
rect 470352 8204 470588 8440
rect 470032 7884 470268 8120
rect 470352 7884 470588 8120
rect 506032 8204 506268 8440
rect 506352 8204 506588 8440
rect 506032 7884 506268 8120
rect 506352 7884 506588 8120
rect 542032 8204 542268 8440
rect 542352 8204 542588 8440
rect 542032 7884 542268 8120
rect 542352 7884 542588 8120
rect 571532 8204 571768 8440
rect 571852 8204 572088 8440
rect 571532 7884 571768 8120
rect 571852 7884 572088 8120
rect 7876 6938 8112 7174
rect 8196 6938 8432 7174
rect 7876 6618 8112 6854
rect 8196 6618 8432 6854
rect 571532 6938 571768 7174
rect 571852 6938 572088 7174
rect 571532 6618 571768 6854
rect 571852 6618 572088 6854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect -5084 -3692 -4848 -3456
rect -4764 -3692 -4528 -3456
rect -5084 -4012 -4848 -3776
rect -4764 -4012 -4528 -3776
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 588452 690938 588688 691174
rect 588772 690938 589008 691174
rect 588452 690618 588688 690854
rect 588772 690618 589008 690854
rect 588452 654938 588688 655174
rect 588772 654938 589008 655174
rect 588452 654618 588688 654854
rect 588772 654618 589008 654854
rect 588452 618938 588688 619174
rect 588772 618938 589008 619174
rect 588452 618618 588688 618854
rect 588772 618618 589008 618854
rect 588452 582938 588688 583174
rect 588772 582938 589008 583174
rect 588452 582618 588688 582854
rect 588772 582618 589008 582854
rect 588452 546938 588688 547174
rect 588772 546938 589008 547174
rect 588452 546618 588688 546854
rect 588772 546618 589008 546854
rect 588452 510938 588688 511174
rect 588772 510938 589008 511174
rect 588452 510618 588688 510854
rect 588772 510618 589008 510854
rect 588452 474938 588688 475174
rect 588772 474938 589008 475174
rect 588452 474618 588688 474854
rect 588772 474618 589008 474854
rect 588452 438938 588688 439174
rect 588772 438938 589008 439174
rect 588452 438618 588688 438854
rect 588772 438618 589008 438854
rect 588452 402938 588688 403174
rect 588772 402938 589008 403174
rect 588452 402618 588688 402854
rect 588772 402618 589008 402854
rect 588452 366938 588688 367174
rect 588772 366938 589008 367174
rect 588452 366618 588688 366854
rect 588772 366618 589008 366854
rect 588452 330938 588688 331174
rect 588772 330938 589008 331174
rect 588452 330618 588688 330854
rect 588772 330618 589008 330854
rect 588452 294938 588688 295174
rect 588772 294938 589008 295174
rect 588452 294618 588688 294854
rect 588772 294618 589008 294854
rect 588452 258938 588688 259174
rect 588772 258938 589008 259174
rect 588452 258618 588688 258854
rect 588772 258618 589008 258854
rect 588452 222938 588688 223174
rect 588772 222938 589008 223174
rect 588452 222618 588688 222854
rect 588772 222618 589008 222854
rect 588452 186938 588688 187174
rect 588772 186938 589008 187174
rect 588452 186618 588688 186854
rect 588772 186618 589008 186854
rect 588452 150938 588688 151174
rect 588772 150938 589008 151174
rect 588452 150618 588688 150854
rect 588772 150618 589008 150854
rect 588452 114938 588688 115174
rect 588772 114938 589008 115174
rect 588452 114618 588688 114854
rect 588772 114618 589008 114854
rect 588452 78938 588688 79174
rect 588772 78938 589008 79174
rect 588452 78618 588688 78854
rect 588772 78618 589008 78854
rect 588452 42938 588688 43174
rect 588772 42938 589008 43174
rect 588452 42618 588688 42854
rect 588772 42618 589008 42854
rect 588452 6938 588688 7174
rect 588772 6938 589008 7174
rect 588452 6618 588688 6854
rect 588772 6618 589008 6854
rect 581546 -3692 581782 -3456
rect 581866 -3692 582102 -3456
rect 581546 -4012 581782 -3776
rect 581866 -4012 582102 -3776
rect -8194 -6802 -7958 -6566
rect -7874 -6802 -7638 -6566
rect -8194 -7122 -7958 -6886
rect -7874 -7122 -7638 -6886
rect -11304 -9912 -11068 -9676
rect -10984 -9912 -10748 -9676
rect -11304 -10232 -11068 -9996
rect -10984 -10232 -10748 -9996
rect -14414 -13022 -14178 -12786
rect -14094 -13022 -13858 -12786
rect -14414 -13342 -14178 -13106
rect -14094 -13342 -13858 -13106
rect -17524 -16132 -17288 -15896
rect -17204 -16132 -16968 -15896
rect -17524 -16452 -17288 -16216
rect -17204 -16452 -16968 -16216
rect -20634 -19242 -20398 -19006
rect -20314 -19242 -20078 -19006
rect -20634 -19562 -20398 -19326
rect -20314 -19562 -20078 -19326
rect -23744 -22352 -23508 -22116
rect -23424 -22352 -23188 -22116
rect -23744 -22672 -23508 -22436
rect -23424 -22672 -23188 -22436
rect 588452 -3692 588688 -3456
rect 588772 -3692 589008 -3456
rect 588452 -4012 588688 -3776
rect 588772 -4012 589008 -3776
rect 591562 694658 591798 694894
rect 591882 694658 592118 694894
rect 591562 694338 591798 694574
rect 591882 694338 592118 694574
rect 591562 658658 591798 658894
rect 591882 658658 592118 658894
rect 591562 658338 591798 658574
rect 591882 658338 592118 658574
rect 591562 622658 591798 622894
rect 591882 622658 592118 622894
rect 591562 622338 591798 622574
rect 591882 622338 592118 622574
rect 591562 586658 591798 586894
rect 591882 586658 592118 586894
rect 591562 586338 591798 586574
rect 591882 586338 592118 586574
rect 591562 550658 591798 550894
rect 591882 550658 592118 550894
rect 591562 550338 591798 550574
rect 591882 550338 592118 550574
rect 591562 514658 591798 514894
rect 591882 514658 592118 514894
rect 591562 514338 591798 514574
rect 591882 514338 592118 514574
rect 591562 478658 591798 478894
rect 591882 478658 592118 478894
rect 591562 478338 591798 478574
rect 591882 478338 592118 478574
rect 591562 442658 591798 442894
rect 591882 442658 592118 442894
rect 591562 442338 591798 442574
rect 591882 442338 592118 442574
rect 591562 406658 591798 406894
rect 591882 406658 592118 406894
rect 591562 406338 591798 406574
rect 591882 406338 592118 406574
rect 591562 370658 591798 370894
rect 591882 370658 592118 370894
rect 591562 370338 591798 370574
rect 591882 370338 592118 370574
rect 591562 334658 591798 334894
rect 591882 334658 592118 334894
rect 591562 334338 591798 334574
rect 591882 334338 592118 334574
rect 591562 298658 591798 298894
rect 591882 298658 592118 298894
rect 591562 298338 591798 298574
rect 591882 298338 592118 298574
rect 591562 262658 591798 262894
rect 591882 262658 592118 262894
rect 591562 262338 591798 262574
rect 591882 262338 592118 262574
rect 591562 226658 591798 226894
rect 591882 226658 592118 226894
rect 591562 226338 591798 226574
rect 591882 226338 592118 226574
rect 591562 190658 591798 190894
rect 591882 190658 592118 190894
rect 591562 190338 591798 190574
rect 591882 190338 592118 190574
rect 591562 154658 591798 154894
rect 591882 154658 592118 154894
rect 591562 154338 591798 154574
rect 591882 154338 592118 154574
rect 591562 118658 591798 118894
rect 591882 118658 592118 118894
rect 591562 118338 591798 118574
rect 591882 118338 592118 118574
rect 591562 82658 591798 82894
rect 591882 82658 592118 82894
rect 591562 82338 591798 82574
rect 591882 82338 592118 82574
rect 591562 46658 591798 46894
rect 591882 46658 592118 46894
rect 591562 46338 591798 46574
rect 591882 46338 592118 46574
rect 591562 10658 591798 10894
rect 591882 10658 592118 10894
rect 591562 10338 591798 10574
rect 591882 10338 592118 10574
rect 591562 -6802 591798 -6566
rect 591882 -6802 592118 -6566
rect 591562 -7122 591798 -6886
rect 591882 -7122 592118 -6886
rect 594672 698378 594908 698614
rect 594992 698378 595228 698614
rect 594672 698058 594908 698294
rect 594992 698058 595228 698294
rect 594672 662378 594908 662614
rect 594992 662378 595228 662614
rect 594672 662058 594908 662294
rect 594992 662058 595228 662294
rect 594672 626378 594908 626614
rect 594992 626378 595228 626614
rect 594672 626058 594908 626294
rect 594992 626058 595228 626294
rect 594672 590378 594908 590614
rect 594992 590378 595228 590614
rect 594672 590058 594908 590294
rect 594992 590058 595228 590294
rect 594672 554378 594908 554614
rect 594992 554378 595228 554614
rect 594672 554058 594908 554294
rect 594992 554058 595228 554294
rect 594672 518378 594908 518614
rect 594992 518378 595228 518614
rect 594672 518058 594908 518294
rect 594992 518058 595228 518294
rect 594672 482378 594908 482614
rect 594992 482378 595228 482614
rect 594672 482058 594908 482294
rect 594992 482058 595228 482294
rect 594672 446378 594908 446614
rect 594992 446378 595228 446614
rect 594672 446058 594908 446294
rect 594992 446058 595228 446294
rect 594672 410378 594908 410614
rect 594992 410378 595228 410614
rect 594672 410058 594908 410294
rect 594992 410058 595228 410294
rect 594672 374378 594908 374614
rect 594992 374378 595228 374614
rect 594672 374058 594908 374294
rect 594992 374058 595228 374294
rect 594672 338378 594908 338614
rect 594992 338378 595228 338614
rect 594672 338058 594908 338294
rect 594992 338058 595228 338294
rect 594672 302378 594908 302614
rect 594992 302378 595228 302614
rect 594672 302058 594908 302294
rect 594992 302058 595228 302294
rect 594672 266378 594908 266614
rect 594992 266378 595228 266614
rect 594672 266058 594908 266294
rect 594992 266058 595228 266294
rect 594672 230378 594908 230614
rect 594992 230378 595228 230614
rect 594672 230058 594908 230294
rect 594992 230058 595228 230294
rect 594672 194378 594908 194614
rect 594992 194378 595228 194614
rect 594672 194058 594908 194294
rect 594992 194058 595228 194294
rect 594672 158378 594908 158614
rect 594992 158378 595228 158614
rect 594672 158058 594908 158294
rect 594992 158058 595228 158294
rect 594672 122378 594908 122614
rect 594992 122378 595228 122614
rect 594672 122058 594908 122294
rect 594992 122058 595228 122294
rect 594672 86378 594908 86614
rect 594992 86378 595228 86614
rect 594672 86058 594908 86294
rect 594992 86058 595228 86294
rect 594672 50378 594908 50614
rect 594992 50378 595228 50614
rect 594672 50058 594908 50294
rect 594992 50058 595228 50294
rect 594672 14378 594908 14614
rect 594992 14378 595228 14614
rect 594672 14058 594908 14294
rect 594992 14058 595228 14294
rect 594672 -9912 594908 -9676
rect 594992 -9912 595228 -9676
rect 594672 -10232 594908 -9996
rect 594992 -10232 595228 -9996
rect 597782 666098 598018 666334
rect 598102 666098 598338 666334
rect 597782 665778 598018 666014
rect 598102 665778 598338 666014
rect 597782 630098 598018 630334
rect 598102 630098 598338 630334
rect 597782 629778 598018 630014
rect 598102 629778 598338 630014
rect 597782 594098 598018 594334
rect 598102 594098 598338 594334
rect 597782 593778 598018 594014
rect 598102 593778 598338 594014
rect 597782 558098 598018 558334
rect 598102 558098 598338 558334
rect 597782 557778 598018 558014
rect 598102 557778 598338 558014
rect 597782 522098 598018 522334
rect 598102 522098 598338 522334
rect 597782 521778 598018 522014
rect 598102 521778 598338 522014
rect 597782 486098 598018 486334
rect 598102 486098 598338 486334
rect 597782 485778 598018 486014
rect 598102 485778 598338 486014
rect 597782 450098 598018 450334
rect 598102 450098 598338 450334
rect 597782 449778 598018 450014
rect 598102 449778 598338 450014
rect 597782 414098 598018 414334
rect 598102 414098 598338 414334
rect 597782 413778 598018 414014
rect 598102 413778 598338 414014
rect 597782 378098 598018 378334
rect 598102 378098 598338 378334
rect 597782 377778 598018 378014
rect 598102 377778 598338 378014
rect 597782 342098 598018 342334
rect 598102 342098 598338 342334
rect 597782 341778 598018 342014
rect 598102 341778 598338 342014
rect 597782 306098 598018 306334
rect 598102 306098 598338 306334
rect 597782 305778 598018 306014
rect 598102 305778 598338 306014
rect 597782 270098 598018 270334
rect 598102 270098 598338 270334
rect 597782 269778 598018 270014
rect 598102 269778 598338 270014
rect 597782 234098 598018 234334
rect 598102 234098 598338 234334
rect 597782 233778 598018 234014
rect 598102 233778 598338 234014
rect 597782 198098 598018 198334
rect 598102 198098 598338 198334
rect 597782 197778 598018 198014
rect 598102 197778 598338 198014
rect 597782 162098 598018 162334
rect 598102 162098 598338 162334
rect 597782 161778 598018 162014
rect 598102 161778 598338 162014
rect 597782 126098 598018 126334
rect 598102 126098 598338 126334
rect 597782 125778 598018 126014
rect 598102 125778 598338 126014
rect 597782 90098 598018 90334
rect 598102 90098 598338 90334
rect 597782 89778 598018 90014
rect 598102 89778 598338 90014
rect 597782 54098 598018 54334
rect 598102 54098 598338 54334
rect 597782 53778 598018 54014
rect 598102 53778 598338 54014
rect 597782 18098 598018 18334
rect 598102 18098 598338 18334
rect 597782 17778 598018 18014
rect 598102 17778 598338 18014
rect 597782 -13022 598018 -12786
rect 598102 -13022 598338 -12786
rect 597782 -13342 598018 -13106
rect 598102 -13342 598338 -13106
rect 600892 669818 601128 670054
rect 601212 669818 601448 670054
rect 600892 669498 601128 669734
rect 601212 669498 601448 669734
rect 600892 633818 601128 634054
rect 601212 633818 601448 634054
rect 600892 633498 601128 633734
rect 601212 633498 601448 633734
rect 600892 597818 601128 598054
rect 601212 597818 601448 598054
rect 600892 597498 601128 597734
rect 601212 597498 601448 597734
rect 600892 561818 601128 562054
rect 601212 561818 601448 562054
rect 600892 561498 601128 561734
rect 601212 561498 601448 561734
rect 600892 525818 601128 526054
rect 601212 525818 601448 526054
rect 600892 525498 601128 525734
rect 601212 525498 601448 525734
rect 600892 489818 601128 490054
rect 601212 489818 601448 490054
rect 600892 489498 601128 489734
rect 601212 489498 601448 489734
rect 600892 453818 601128 454054
rect 601212 453818 601448 454054
rect 600892 453498 601128 453734
rect 601212 453498 601448 453734
rect 600892 417818 601128 418054
rect 601212 417818 601448 418054
rect 600892 417498 601128 417734
rect 601212 417498 601448 417734
rect 600892 381818 601128 382054
rect 601212 381818 601448 382054
rect 600892 381498 601128 381734
rect 601212 381498 601448 381734
rect 600892 345818 601128 346054
rect 601212 345818 601448 346054
rect 600892 345498 601128 345734
rect 601212 345498 601448 345734
rect 600892 309818 601128 310054
rect 601212 309818 601448 310054
rect 600892 309498 601128 309734
rect 601212 309498 601448 309734
rect 600892 273818 601128 274054
rect 601212 273818 601448 274054
rect 600892 273498 601128 273734
rect 601212 273498 601448 273734
rect 600892 237818 601128 238054
rect 601212 237818 601448 238054
rect 600892 237498 601128 237734
rect 601212 237498 601448 237734
rect 600892 201818 601128 202054
rect 601212 201818 601448 202054
rect 600892 201498 601128 201734
rect 601212 201498 601448 201734
rect 600892 165818 601128 166054
rect 601212 165818 601448 166054
rect 600892 165498 601128 165734
rect 601212 165498 601448 165734
rect 600892 129818 601128 130054
rect 601212 129818 601448 130054
rect 600892 129498 601128 129734
rect 601212 129498 601448 129734
rect 600892 93818 601128 94054
rect 601212 93818 601448 94054
rect 600892 93498 601128 93734
rect 601212 93498 601448 93734
rect 600892 57818 601128 58054
rect 601212 57818 601448 58054
rect 600892 57498 601128 57734
rect 601212 57498 601448 57734
rect 600892 -16132 601128 -15896
rect 601212 -16132 601448 -15896
rect 600892 -16452 601128 -16216
rect 601212 -16452 601448 -16216
rect 604002 673538 604238 673774
rect 604322 673538 604558 673774
rect 604002 673218 604238 673454
rect 604322 673218 604558 673454
rect 604002 637538 604238 637774
rect 604322 637538 604558 637774
rect 604002 637218 604238 637454
rect 604322 637218 604558 637454
rect 604002 601538 604238 601774
rect 604322 601538 604558 601774
rect 604002 601218 604238 601454
rect 604322 601218 604558 601454
rect 604002 565538 604238 565774
rect 604322 565538 604558 565774
rect 604002 565218 604238 565454
rect 604322 565218 604558 565454
rect 604002 529538 604238 529774
rect 604322 529538 604558 529774
rect 604002 529218 604238 529454
rect 604322 529218 604558 529454
rect 604002 493538 604238 493774
rect 604322 493538 604558 493774
rect 604002 493218 604238 493454
rect 604322 493218 604558 493454
rect 604002 457538 604238 457774
rect 604322 457538 604558 457774
rect 604002 457218 604238 457454
rect 604322 457218 604558 457454
rect 604002 421538 604238 421774
rect 604322 421538 604558 421774
rect 604002 421218 604238 421454
rect 604322 421218 604558 421454
rect 604002 385538 604238 385774
rect 604322 385538 604558 385774
rect 604002 385218 604238 385454
rect 604322 385218 604558 385454
rect 604002 349538 604238 349774
rect 604322 349538 604558 349774
rect 604002 349218 604238 349454
rect 604322 349218 604558 349454
rect 604002 313538 604238 313774
rect 604322 313538 604558 313774
rect 604002 313218 604238 313454
rect 604322 313218 604558 313454
rect 604002 277538 604238 277774
rect 604322 277538 604558 277774
rect 604002 277218 604238 277454
rect 604322 277218 604558 277454
rect 604002 241538 604238 241774
rect 604322 241538 604558 241774
rect 604002 241218 604238 241454
rect 604322 241218 604558 241454
rect 604002 205538 604238 205774
rect 604322 205538 604558 205774
rect 604002 205218 604238 205454
rect 604322 205218 604558 205454
rect 604002 169538 604238 169774
rect 604322 169538 604558 169774
rect 604002 169218 604238 169454
rect 604322 169218 604558 169454
rect 604002 133538 604238 133774
rect 604322 133538 604558 133774
rect 604002 133218 604238 133454
rect 604322 133218 604558 133454
rect 604002 97538 604238 97774
rect 604322 97538 604558 97774
rect 604002 97218 604238 97454
rect 604322 97218 604558 97454
rect 604002 61538 604238 61774
rect 604322 61538 604558 61774
rect 604002 61218 604238 61454
rect 604322 61218 604558 61454
rect 604002 25538 604238 25774
rect 604322 25538 604558 25774
rect 604002 25218 604238 25454
rect 604322 25218 604558 25454
rect 604002 -19242 604238 -19006
rect 604322 -19242 604558 -19006
rect 604002 -19562 604238 -19326
rect 604322 -19562 604558 -19326
rect 607112 677258 607348 677494
rect 607432 677258 607668 677494
rect 607112 676938 607348 677174
rect 607432 676938 607668 677174
rect 607112 641258 607348 641494
rect 607432 641258 607668 641494
rect 607112 640938 607348 641174
rect 607432 640938 607668 641174
rect 607112 605258 607348 605494
rect 607432 605258 607668 605494
rect 607112 604938 607348 605174
rect 607432 604938 607668 605174
rect 607112 569258 607348 569494
rect 607432 569258 607668 569494
rect 607112 568938 607348 569174
rect 607432 568938 607668 569174
rect 607112 533258 607348 533494
rect 607432 533258 607668 533494
rect 607112 532938 607348 533174
rect 607432 532938 607668 533174
rect 607112 497258 607348 497494
rect 607432 497258 607668 497494
rect 607112 496938 607348 497174
rect 607432 496938 607668 497174
rect 607112 461258 607348 461494
rect 607432 461258 607668 461494
rect 607112 460938 607348 461174
rect 607432 460938 607668 461174
rect 607112 425258 607348 425494
rect 607432 425258 607668 425494
rect 607112 424938 607348 425174
rect 607432 424938 607668 425174
rect 607112 389258 607348 389494
rect 607432 389258 607668 389494
rect 607112 388938 607348 389174
rect 607432 388938 607668 389174
rect 607112 353258 607348 353494
rect 607432 353258 607668 353494
rect 607112 352938 607348 353174
rect 607432 352938 607668 353174
rect 607112 317258 607348 317494
rect 607432 317258 607668 317494
rect 607112 316938 607348 317174
rect 607432 316938 607668 317174
rect 607112 281258 607348 281494
rect 607432 281258 607668 281494
rect 607112 280938 607348 281174
rect 607432 280938 607668 281174
rect 607112 245258 607348 245494
rect 607432 245258 607668 245494
rect 607112 244938 607348 245174
rect 607432 244938 607668 245174
rect 607112 209258 607348 209494
rect 607432 209258 607668 209494
rect 607112 208938 607348 209174
rect 607432 208938 607668 209174
rect 607112 173258 607348 173494
rect 607432 173258 607668 173494
rect 607112 172938 607348 173174
rect 607432 172938 607668 173174
rect 607112 137258 607348 137494
rect 607432 137258 607668 137494
rect 607112 136938 607348 137174
rect 607432 136938 607668 137174
rect 607112 101258 607348 101494
rect 607432 101258 607668 101494
rect 607112 100938 607348 101174
rect 607432 100938 607668 101174
rect 607112 65258 607348 65494
rect 607432 65258 607668 65494
rect 607112 64938 607348 65174
rect 607432 64938 607668 65174
rect 607112 29258 607348 29494
rect 607432 29258 607668 29494
rect 607112 28938 607348 29174
rect 607432 28938 607668 29174
rect 607112 -22352 607348 -22116
rect 607432 -22352 607668 -22116
rect 607112 -22672 607348 -22436
rect 607432 -22672 607668 -22436
<< metal5 >>
rect -23776 726608 607700 726640
rect -23776 726372 -23744 726608
rect -23508 726372 -23424 726608
rect -23188 726372 607112 726608
rect 607348 726372 607432 726608
rect 607668 726372 607700 726608
rect -23776 726288 607700 726372
rect -23776 726052 -23744 726288
rect -23508 726052 -23424 726288
rect -23188 726052 607112 726288
rect 607348 726052 607432 726288
rect 607668 726052 607700 726288
rect -23776 726020 607700 726052
rect -20666 723498 604590 723530
rect -20666 723262 -20634 723498
rect -20398 723262 -20314 723498
rect -20078 723262 604002 723498
rect 604238 723262 604322 723498
rect 604558 723262 604590 723498
rect -20666 723178 604590 723262
rect -20666 722942 -20634 723178
rect -20398 722942 -20314 723178
rect -20078 722942 604002 723178
rect 604238 722942 604322 723178
rect 604558 722942 604590 723178
rect -20666 722910 604590 722942
rect -17556 720388 601480 720420
rect -17556 720152 -17524 720388
rect -17288 720152 -17204 720388
rect -16968 720152 600892 720388
rect 601128 720152 601212 720388
rect 601448 720152 601480 720388
rect -17556 720068 601480 720152
rect -17556 719832 -17524 720068
rect -17288 719832 -17204 720068
rect -16968 719832 600892 720068
rect 601128 719832 601212 720068
rect 601448 719832 601480 720068
rect -17556 719800 601480 719832
rect -14446 717278 598370 717310
rect -14446 717042 -14414 717278
rect -14178 717042 -14094 717278
rect -13858 717042 597782 717278
rect 598018 717042 598102 717278
rect 598338 717042 598370 717278
rect -14446 716958 598370 717042
rect -14446 716722 -14414 716958
rect -14178 716722 -14094 716958
rect -13858 716722 597782 716958
rect 598018 716722 598102 716958
rect 598338 716722 598370 716958
rect -14446 716690 598370 716722
rect -11336 714168 595260 714200
rect -11336 713932 -11304 714168
rect -11068 713932 -10984 714168
rect -10748 713932 594672 714168
rect 594908 713932 594992 714168
rect 595228 713932 595260 714168
rect -11336 713848 595260 713932
rect -11336 713612 -11304 713848
rect -11068 713612 -10984 713848
rect -10748 713612 594672 713848
rect 594908 713612 594992 713848
rect 595228 713612 595260 713848
rect -11336 713580 595260 713612
rect -8226 711058 592150 711090
rect -8226 710822 -8194 711058
rect -7958 710822 -7874 711058
rect -7638 710822 591562 711058
rect 591798 710822 591882 711058
rect 592118 710822 592150 711058
rect -8226 710738 592150 710822
rect -8226 710502 -8194 710738
rect -7958 710502 -7874 710738
rect -7638 710502 591562 710738
rect 591798 710502 591882 710738
rect 592118 710502 592150 710738
rect -8226 710470 592150 710502
rect -5116 707948 589040 707980
rect -5116 707712 -5084 707948
rect -4848 707712 -4764 707948
rect -4528 707712 581546 707948
rect 581782 707712 581866 707948
rect 582102 707712 588452 707948
rect 588688 707712 588772 707948
rect 589008 707712 589040 707948
rect -5116 707628 589040 707712
rect -5116 707392 -5084 707628
rect -4848 707392 -4764 707628
rect -4528 707392 581546 707628
rect 581782 707392 581866 707628
rect 582102 707392 588452 707628
rect 588688 707392 588772 707628
rect 589008 707392 589040 707628
rect -5116 707360 589040 707392
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -23776 698614 607700 698646
rect -23776 698378 -11304 698614
rect -11068 698378 -10984 698614
rect -10748 698378 594672 698614
rect 594908 698378 594992 698614
rect 595228 698378 607700 698614
rect -23776 698294 607700 698378
rect -23776 698058 -11304 698294
rect -11068 698058 -10984 698294
rect -10748 698058 594672 698294
rect 594908 698058 594992 698294
rect 595228 698058 607700 698294
rect -23776 698026 607700 698058
rect -23776 694894 607700 694926
rect -23776 694658 -8194 694894
rect -7958 694658 -7874 694894
rect -7638 694658 591562 694894
rect 591798 694658 591882 694894
rect 592118 694658 607700 694894
rect -23776 694574 607700 694658
rect -23776 694338 -8194 694574
rect -7958 694338 -7874 694574
rect -7638 694338 591562 694574
rect 591798 694338 591882 694574
rect 592118 694338 607700 694574
rect -23776 694306 607700 694338
rect 7852 693716 8456 693748
rect 7852 693480 7876 693716
rect 8112 693480 8196 693716
rect 8432 693480 8456 693716
rect 7852 693396 8456 693480
rect 7852 693160 7876 693396
rect 8112 693160 8196 693396
rect 8432 693160 8456 693396
rect 7852 693128 8456 693160
rect 38008 693716 38612 693748
rect 38008 693480 38032 693716
rect 38268 693480 38352 693716
rect 38588 693480 38612 693716
rect 38008 693396 38612 693480
rect 38008 693160 38032 693396
rect 38268 693160 38352 693396
rect 38588 693160 38612 693396
rect 38008 693128 38612 693160
rect 74008 693716 74612 693748
rect 74008 693480 74032 693716
rect 74268 693480 74352 693716
rect 74588 693480 74612 693716
rect 74008 693396 74612 693480
rect 74008 693160 74032 693396
rect 74268 693160 74352 693396
rect 74588 693160 74612 693396
rect 74008 693128 74612 693160
rect 110008 693716 110612 693748
rect 110008 693480 110032 693716
rect 110268 693480 110352 693716
rect 110588 693480 110612 693716
rect 110008 693396 110612 693480
rect 110008 693160 110032 693396
rect 110268 693160 110352 693396
rect 110588 693160 110612 693396
rect 110008 693128 110612 693160
rect 146008 693716 146612 693748
rect 146008 693480 146032 693716
rect 146268 693480 146352 693716
rect 146588 693480 146612 693716
rect 146008 693396 146612 693480
rect 146008 693160 146032 693396
rect 146268 693160 146352 693396
rect 146588 693160 146612 693396
rect 146008 693128 146612 693160
rect 182008 693716 182612 693748
rect 182008 693480 182032 693716
rect 182268 693480 182352 693716
rect 182588 693480 182612 693716
rect 182008 693396 182612 693480
rect 182008 693160 182032 693396
rect 182268 693160 182352 693396
rect 182588 693160 182612 693396
rect 182008 693128 182612 693160
rect 218008 693716 218612 693748
rect 218008 693480 218032 693716
rect 218268 693480 218352 693716
rect 218588 693480 218612 693716
rect 218008 693396 218612 693480
rect 218008 693160 218032 693396
rect 218268 693160 218352 693396
rect 218588 693160 218612 693396
rect 218008 693128 218612 693160
rect 254008 693716 254612 693748
rect 254008 693480 254032 693716
rect 254268 693480 254352 693716
rect 254588 693480 254612 693716
rect 254008 693396 254612 693480
rect 254008 693160 254032 693396
rect 254268 693160 254352 693396
rect 254588 693160 254612 693396
rect 254008 693128 254612 693160
rect 290008 693716 290612 693748
rect 290008 693480 290032 693716
rect 290268 693480 290352 693716
rect 290588 693480 290612 693716
rect 290008 693396 290612 693480
rect 290008 693160 290032 693396
rect 290268 693160 290352 693396
rect 290588 693160 290612 693396
rect 290008 693128 290612 693160
rect 326008 693716 326612 693748
rect 326008 693480 326032 693716
rect 326268 693480 326352 693716
rect 326588 693480 326612 693716
rect 326008 693396 326612 693480
rect 326008 693160 326032 693396
rect 326268 693160 326352 693396
rect 326588 693160 326612 693396
rect 326008 693128 326612 693160
rect 362008 693716 362612 693748
rect 362008 693480 362032 693716
rect 362268 693480 362352 693716
rect 362588 693480 362612 693716
rect 362008 693396 362612 693480
rect 362008 693160 362032 693396
rect 362268 693160 362352 693396
rect 362588 693160 362612 693396
rect 362008 693128 362612 693160
rect 398008 693716 398612 693748
rect 398008 693480 398032 693716
rect 398268 693480 398352 693716
rect 398588 693480 398612 693716
rect 398008 693396 398612 693480
rect 398008 693160 398032 693396
rect 398268 693160 398352 693396
rect 398588 693160 398612 693396
rect 398008 693128 398612 693160
rect 434008 693716 434612 693748
rect 434008 693480 434032 693716
rect 434268 693480 434352 693716
rect 434588 693480 434612 693716
rect 434008 693396 434612 693480
rect 434008 693160 434032 693396
rect 434268 693160 434352 693396
rect 434588 693160 434612 693396
rect 434008 693128 434612 693160
rect 470008 693716 470612 693748
rect 470008 693480 470032 693716
rect 470268 693480 470352 693716
rect 470588 693480 470612 693716
rect 470008 693396 470612 693480
rect 470008 693160 470032 693396
rect 470268 693160 470352 693396
rect 470588 693160 470612 693396
rect 470008 693128 470612 693160
rect 506008 693716 506612 693748
rect 506008 693480 506032 693716
rect 506268 693480 506352 693716
rect 506588 693480 506612 693716
rect 506008 693396 506612 693480
rect 506008 693160 506032 693396
rect 506268 693160 506352 693396
rect 506588 693160 506612 693396
rect 506008 693128 506612 693160
rect 542008 693716 542612 693748
rect 542008 693480 542032 693716
rect 542268 693480 542352 693716
rect 542588 693480 542612 693716
rect 542008 693396 542612 693480
rect 542008 693160 542032 693396
rect 542268 693160 542352 693396
rect 542588 693160 542612 693396
rect 542008 693128 542612 693160
rect 571508 693716 572112 693748
rect 571508 693480 571532 693716
rect 571768 693480 571852 693716
rect 572088 693480 572112 693716
rect 571508 693396 572112 693480
rect 571508 693160 571532 693396
rect 571768 693160 571852 693396
rect 572088 693160 572112 693396
rect 571508 693128 572112 693160
rect 9092 692476 9696 692508
rect 9092 692240 9116 692476
rect 9352 692240 9436 692476
rect 9672 692240 9696 692476
rect 9092 692156 9696 692240
rect 9092 691920 9116 692156
rect 9352 691920 9436 692156
rect 9672 691920 9696 692156
rect 9092 691888 9696 691920
rect 56628 692476 57232 692508
rect 56628 692240 56652 692476
rect 56888 692240 56972 692476
rect 57208 692240 57232 692476
rect 56628 692156 57232 692240
rect 56628 691920 56652 692156
rect 56888 691920 56972 692156
rect 57208 691920 57232 692156
rect 56628 691888 57232 691920
rect 92628 692476 93232 692508
rect 92628 692240 92652 692476
rect 92888 692240 92972 692476
rect 93208 692240 93232 692476
rect 92628 692156 93232 692240
rect 92628 691920 92652 692156
rect 92888 691920 92972 692156
rect 93208 691920 93232 692156
rect 92628 691888 93232 691920
rect 128628 692476 129232 692508
rect 128628 692240 128652 692476
rect 128888 692240 128972 692476
rect 129208 692240 129232 692476
rect 128628 692156 129232 692240
rect 128628 691920 128652 692156
rect 128888 691920 128972 692156
rect 129208 691920 129232 692156
rect 128628 691888 129232 691920
rect 164628 692476 165232 692508
rect 164628 692240 164652 692476
rect 164888 692240 164972 692476
rect 165208 692240 165232 692476
rect 164628 692156 165232 692240
rect 164628 691920 164652 692156
rect 164888 691920 164972 692156
rect 165208 691920 165232 692156
rect 164628 691888 165232 691920
rect 200628 692476 201232 692508
rect 200628 692240 200652 692476
rect 200888 692240 200972 692476
rect 201208 692240 201232 692476
rect 200628 692156 201232 692240
rect 200628 691920 200652 692156
rect 200888 691920 200972 692156
rect 201208 691920 201232 692156
rect 200628 691888 201232 691920
rect 236628 692476 237232 692508
rect 236628 692240 236652 692476
rect 236888 692240 236972 692476
rect 237208 692240 237232 692476
rect 236628 692156 237232 692240
rect 236628 691920 236652 692156
rect 236888 691920 236972 692156
rect 237208 691920 237232 692156
rect 236628 691888 237232 691920
rect 272628 692476 273232 692508
rect 272628 692240 272652 692476
rect 272888 692240 272972 692476
rect 273208 692240 273232 692476
rect 272628 692156 273232 692240
rect 272628 691920 272652 692156
rect 272888 691920 272972 692156
rect 273208 691920 273232 692156
rect 272628 691888 273232 691920
rect 308628 692476 309232 692508
rect 308628 692240 308652 692476
rect 308888 692240 308972 692476
rect 309208 692240 309232 692476
rect 308628 692156 309232 692240
rect 308628 691920 308652 692156
rect 308888 691920 308972 692156
rect 309208 691920 309232 692156
rect 308628 691888 309232 691920
rect 344628 692476 345232 692508
rect 344628 692240 344652 692476
rect 344888 692240 344972 692476
rect 345208 692240 345232 692476
rect 344628 692156 345232 692240
rect 344628 691920 344652 692156
rect 344888 691920 344972 692156
rect 345208 691920 345232 692156
rect 344628 691888 345232 691920
rect 380628 692476 381232 692508
rect 380628 692240 380652 692476
rect 380888 692240 380972 692476
rect 381208 692240 381232 692476
rect 380628 692156 381232 692240
rect 380628 691920 380652 692156
rect 380888 691920 380972 692156
rect 381208 691920 381232 692156
rect 380628 691888 381232 691920
rect 416628 692476 417232 692508
rect 416628 692240 416652 692476
rect 416888 692240 416972 692476
rect 417208 692240 417232 692476
rect 416628 692156 417232 692240
rect 416628 691920 416652 692156
rect 416888 691920 416972 692156
rect 417208 691920 417232 692156
rect 416628 691888 417232 691920
rect 452628 692476 453232 692508
rect 452628 692240 452652 692476
rect 452888 692240 452972 692476
rect 453208 692240 453232 692476
rect 452628 692156 453232 692240
rect 452628 691920 452652 692156
rect 452888 691920 452972 692156
rect 453208 691920 453232 692156
rect 452628 691888 453232 691920
rect 488628 692476 489232 692508
rect 488628 692240 488652 692476
rect 488888 692240 488972 692476
rect 489208 692240 489232 692476
rect 488628 692156 489232 692240
rect 488628 691920 488652 692156
rect 488888 691920 488972 692156
rect 489208 691920 489232 692156
rect 488628 691888 489232 691920
rect 524628 692476 525232 692508
rect 524628 692240 524652 692476
rect 524888 692240 524972 692476
rect 525208 692240 525232 692476
rect 524628 692156 525232 692240
rect 524628 691920 524652 692156
rect 524888 691920 524972 692156
rect 525208 691920 525232 692156
rect 524628 691888 525232 691920
rect 560628 692476 561232 692508
rect 560628 692240 560652 692476
rect 560888 692240 560972 692476
rect 561208 692240 561232 692476
rect 560628 692156 561232 692240
rect 560628 691920 560652 692156
rect 560888 691920 560972 692156
rect 561208 691920 561232 692156
rect 560628 691888 561232 691920
rect 570268 692476 570872 692508
rect 570268 692240 570292 692476
rect 570528 692240 570612 692476
rect 570848 692240 570872 692476
rect 570268 692156 570872 692240
rect 570268 691920 570292 692156
rect 570528 691920 570612 692156
rect 570848 691920 570872 692156
rect 570268 691888 570872 691920
rect -23776 691174 607700 691206
rect -23776 690938 -5084 691174
rect -4848 690938 -4764 691174
rect -4528 690938 7876 691174
rect 8112 690938 8196 691174
rect 8432 690938 38032 691174
rect 38268 690938 38352 691174
rect 38588 690938 74032 691174
rect 74268 690938 74352 691174
rect 74588 690938 110032 691174
rect 110268 690938 110352 691174
rect 110588 690938 146032 691174
rect 146268 690938 146352 691174
rect 146588 690938 182032 691174
rect 182268 690938 182352 691174
rect 182588 690938 218032 691174
rect 218268 690938 218352 691174
rect 218588 690938 254032 691174
rect 254268 690938 254352 691174
rect 254588 690938 290032 691174
rect 290268 690938 290352 691174
rect 290588 690938 326032 691174
rect 326268 690938 326352 691174
rect 326588 690938 362032 691174
rect 362268 690938 362352 691174
rect 362588 690938 398032 691174
rect 398268 690938 398352 691174
rect 398588 690938 434032 691174
rect 434268 690938 434352 691174
rect 434588 690938 470032 691174
rect 470268 690938 470352 691174
rect 470588 690938 506032 691174
rect 506268 690938 506352 691174
rect 506588 690938 542032 691174
rect 542268 690938 542352 691174
rect 542588 690938 571532 691174
rect 571768 690938 571852 691174
rect 572088 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 588452 691174
rect 588688 690938 588772 691174
rect 589008 690938 607700 691174
rect -23776 690854 607700 690938
rect -23776 690618 -5084 690854
rect -4848 690618 -4764 690854
rect -4528 690618 7876 690854
rect 8112 690618 8196 690854
rect 8432 690618 38032 690854
rect 38268 690618 38352 690854
rect 38588 690618 74032 690854
rect 74268 690618 74352 690854
rect 74588 690618 110032 690854
rect 110268 690618 110352 690854
rect 110588 690618 146032 690854
rect 146268 690618 146352 690854
rect 146588 690618 182032 690854
rect 182268 690618 182352 690854
rect 182588 690618 218032 690854
rect 218268 690618 218352 690854
rect 218588 690618 254032 690854
rect 254268 690618 254352 690854
rect 254588 690618 290032 690854
rect 290268 690618 290352 690854
rect 290588 690618 326032 690854
rect 326268 690618 326352 690854
rect 326588 690618 362032 690854
rect 362268 690618 362352 690854
rect 362588 690618 398032 690854
rect 398268 690618 398352 690854
rect 398588 690618 434032 690854
rect 434268 690618 434352 690854
rect 434588 690618 470032 690854
rect 470268 690618 470352 690854
rect 470588 690618 506032 690854
rect 506268 690618 506352 690854
rect 506588 690618 542032 690854
rect 542268 690618 542352 690854
rect 542588 690618 571532 690854
rect 571768 690618 571852 690854
rect 572088 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 588452 690854
rect 588688 690618 588772 690854
rect 589008 690618 607700 690854
rect -23776 690586 607700 690618
rect -23776 687454 607700 687486
rect -23776 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 9116 687454
rect 9352 687218 9436 687454
rect 9672 687218 56652 687454
rect 56888 687218 56972 687454
rect 57208 687218 92652 687454
rect 92888 687218 92972 687454
rect 93208 687218 128652 687454
rect 128888 687218 128972 687454
rect 129208 687218 164652 687454
rect 164888 687218 164972 687454
rect 165208 687218 200652 687454
rect 200888 687218 200972 687454
rect 201208 687218 236652 687454
rect 236888 687218 236972 687454
rect 237208 687218 272652 687454
rect 272888 687218 272972 687454
rect 273208 687218 308652 687454
rect 308888 687218 308972 687454
rect 309208 687218 344652 687454
rect 344888 687218 344972 687454
rect 345208 687218 380652 687454
rect 380888 687218 380972 687454
rect 381208 687218 416652 687454
rect 416888 687218 416972 687454
rect 417208 687218 452652 687454
rect 452888 687218 452972 687454
rect 453208 687218 488652 687454
rect 488888 687218 488972 687454
rect 489208 687218 524652 687454
rect 524888 687218 524972 687454
rect 525208 687218 560652 687454
rect 560888 687218 560972 687454
rect 561208 687218 570292 687454
rect 570528 687218 570612 687454
rect 570848 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 607700 687454
rect -23776 687134 607700 687218
rect -23776 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 9116 687134
rect 9352 686898 9436 687134
rect 9672 686898 56652 687134
rect 56888 686898 56972 687134
rect 57208 686898 92652 687134
rect 92888 686898 92972 687134
rect 93208 686898 128652 687134
rect 128888 686898 128972 687134
rect 129208 686898 164652 687134
rect 164888 686898 164972 687134
rect 165208 686898 200652 687134
rect 200888 686898 200972 687134
rect 201208 686898 236652 687134
rect 236888 686898 236972 687134
rect 237208 686898 272652 687134
rect 272888 686898 272972 687134
rect 273208 686898 308652 687134
rect 308888 686898 308972 687134
rect 309208 686898 344652 687134
rect 344888 686898 344972 687134
rect 345208 686898 380652 687134
rect 380888 686898 380972 687134
rect 381208 686898 416652 687134
rect 416888 686898 416972 687134
rect 417208 686898 452652 687134
rect 452888 686898 452972 687134
rect 453208 686898 488652 687134
rect 488888 686898 488972 687134
rect 489208 686898 524652 687134
rect 524888 686898 524972 687134
rect 525208 686898 560652 687134
rect 560888 686898 560972 687134
rect 561208 686898 570292 687134
rect 570528 686898 570612 687134
rect 570848 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 607700 687134
rect -23776 686866 607700 686898
rect -23776 677494 607700 677526
rect -23776 677258 -23744 677494
rect -23508 677258 -23424 677494
rect -23188 677258 607112 677494
rect 607348 677258 607432 677494
rect 607668 677258 607700 677494
rect -23776 677174 607700 677258
rect -23776 676938 -23744 677174
rect -23508 676938 -23424 677174
rect -23188 676938 607112 677174
rect 607348 676938 607432 677174
rect 607668 676938 607700 677174
rect -23776 676906 607700 676938
rect -23776 673774 607700 673806
rect -23776 673538 -20634 673774
rect -20398 673538 -20314 673774
rect -20078 673538 604002 673774
rect 604238 673538 604322 673774
rect 604558 673538 607700 673774
rect -23776 673454 607700 673538
rect -23776 673218 -20634 673454
rect -20398 673218 -20314 673454
rect -20078 673218 604002 673454
rect 604238 673218 604322 673454
rect 604558 673218 607700 673454
rect -23776 673186 607700 673218
rect -23776 670054 607700 670086
rect -23776 669818 -17524 670054
rect -17288 669818 -17204 670054
rect -16968 669818 600892 670054
rect 601128 669818 601212 670054
rect 601448 669818 607700 670054
rect -23776 669734 607700 669818
rect -23776 669498 -17524 669734
rect -17288 669498 -17204 669734
rect -16968 669498 600892 669734
rect 601128 669498 601212 669734
rect 601448 669498 607700 669734
rect -23776 669466 607700 669498
rect -23776 666334 607700 666366
rect -23776 666098 -14414 666334
rect -14178 666098 -14094 666334
rect -13858 666098 597782 666334
rect 598018 666098 598102 666334
rect 598338 666098 607700 666334
rect -23776 666014 607700 666098
rect -23776 665778 -14414 666014
rect -14178 665778 -14094 666014
rect -13858 665778 597782 666014
rect 598018 665778 598102 666014
rect 598338 665778 607700 666014
rect -23776 665746 607700 665778
rect -23776 662614 607700 662646
rect -23776 662378 -11304 662614
rect -11068 662378 -10984 662614
rect -10748 662378 594672 662614
rect 594908 662378 594992 662614
rect 595228 662378 607700 662614
rect -23776 662294 607700 662378
rect -23776 662058 -11304 662294
rect -11068 662058 -10984 662294
rect -10748 662058 594672 662294
rect 594908 662058 594992 662294
rect 595228 662058 607700 662294
rect -23776 662026 607700 662058
rect -23776 658894 607700 658926
rect -23776 658658 -8194 658894
rect -7958 658658 -7874 658894
rect -7638 658658 591562 658894
rect 591798 658658 591882 658894
rect 592118 658658 607700 658894
rect -23776 658574 607700 658658
rect -23776 658338 -8194 658574
rect -7958 658338 -7874 658574
rect -7638 658338 591562 658574
rect 591798 658338 591882 658574
rect 592118 658338 607700 658574
rect -23776 658306 607700 658338
rect -23776 655174 607700 655206
rect -23776 654938 -5084 655174
rect -4848 654938 -4764 655174
rect -4528 654938 7876 655174
rect 8112 654938 8196 655174
rect 8432 654938 38032 655174
rect 38268 654938 38352 655174
rect 38588 654938 74032 655174
rect 74268 654938 74352 655174
rect 74588 654938 110032 655174
rect 110268 654938 110352 655174
rect 110588 654938 146032 655174
rect 146268 654938 146352 655174
rect 146588 654938 182032 655174
rect 182268 654938 182352 655174
rect 182588 654938 218032 655174
rect 218268 654938 218352 655174
rect 218588 654938 254032 655174
rect 254268 654938 254352 655174
rect 254588 654938 290032 655174
rect 290268 654938 290352 655174
rect 290588 654938 326032 655174
rect 326268 654938 326352 655174
rect 326588 654938 362032 655174
rect 362268 654938 362352 655174
rect 362588 654938 398032 655174
rect 398268 654938 398352 655174
rect 398588 654938 434032 655174
rect 434268 654938 434352 655174
rect 434588 654938 470032 655174
rect 470268 654938 470352 655174
rect 470588 654938 506032 655174
rect 506268 654938 506352 655174
rect 506588 654938 542032 655174
rect 542268 654938 542352 655174
rect 542588 654938 571532 655174
rect 571768 654938 571852 655174
rect 572088 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 588452 655174
rect 588688 654938 588772 655174
rect 589008 654938 607700 655174
rect -23776 654854 607700 654938
rect -23776 654618 -5084 654854
rect -4848 654618 -4764 654854
rect -4528 654618 7876 654854
rect 8112 654618 8196 654854
rect 8432 654618 38032 654854
rect 38268 654618 38352 654854
rect 38588 654618 74032 654854
rect 74268 654618 74352 654854
rect 74588 654618 110032 654854
rect 110268 654618 110352 654854
rect 110588 654618 146032 654854
rect 146268 654618 146352 654854
rect 146588 654618 182032 654854
rect 182268 654618 182352 654854
rect 182588 654618 218032 654854
rect 218268 654618 218352 654854
rect 218588 654618 254032 654854
rect 254268 654618 254352 654854
rect 254588 654618 290032 654854
rect 290268 654618 290352 654854
rect 290588 654618 326032 654854
rect 326268 654618 326352 654854
rect 326588 654618 362032 654854
rect 362268 654618 362352 654854
rect 362588 654618 398032 654854
rect 398268 654618 398352 654854
rect 398588 654618 434032 654854
rect 434268 654618 434352 654854
rect 434588 654618 470032 654854
rect 470268 654618 470352 654854
rect 470588 654618 506032 654854
rect 506268 654618 506352 654854
rect 506588 654618 542032 654854
rect 542268 654618 542352 654854
rect 542588 654618 571532 654854
rect 571768 654618 571852 654854
rect 572088 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 588452 654854
rect 588688 654618 588772 654854
rect 589008 654618 607700 654854
rect -23776 654586 607700 654618
rect -23776 651454 607700 651486
rect -23776 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 9116 651454
rect 9352 651218 9436 651454
rect 9672 651218 56652 651454
rect 56888 651218 56972 651454
rect 57208 651218 92652 651454
rect 92888 651218 92972 651454
rect 93208 651218 128652 651454
rect 128888 651218 128972 651454
rect 129208 651218 164652 651454
rect 164888 651218 164972 651454
rect 165208 651218 200652 651454
rect 200888 651218 200972 651454
rect 201208 651218 236652 651454
rect 236888 651218 236972 651454
rect 237208 651218 272652 651454
rect 272888 651218 272972 651454
rect 273208 651218 308652 651454
rect 308888 651218 308972 651454
rect 309208 651218 344652 651454
rect 344888 651218 344972 651454
rect 345208 651218 380652 651454
rect 380888 651218 380972 651454
rect 381208 651218 416652 651454
rect 416888 651218 416972 651454
rect 417208 651218 452652 651454
rect 452888 651218 452972 651454
rect 453208 651218 488652 651454
rect 488888 651218 488972 651454
rect 489208 651218 524652 651454
rect 524888 651218 524972 651454
rect 525208 651218 560652 651454
rect 560888 651218 560972 651454
rect 561208 651218 570292 651454
rect 570528 651218 570612 651454
rect 570848 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 607700 651454
rect -23776 651134 607700 651218
rect -23776 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 9116 651134
rect 9352 650898 9436 651134
rect 9672 650898 56652 651134
rect 56888 650898 56972 651134
rect 57208 650898 92652 651134
rect 92888 650898 92972 651134
rect 93208 650898 128652 651134
rect 128888 650898 128972 651134
rect 129208 650898 164652 651134
rect 164888 650898 164972 651134
rect 165208 650898 200652 651134
rect 200888 650898 200972 651134
rect 201208 650898 236652 651134
rect 236888 650898 236972 651134
rect 237208 650898 272652 651134
rect 272888 650898 272972 651134
rect 273208 650898 308652 651134
rect 308888 650898 308972 651134
rect 309208 650898 344652 651134
rect 344888 650898 344972 651134
rect 345208 650898 380652 651134
rect 380888 650898 380972 651134
rect 381208 650898 416652 651134
rect 416888 650898 416972 651134
rect 417208 650898 452652 651134
rect 452888 650898 452972 651134
rect 453208 650898 488652 651134
rect 488888 650898 488972 651134
rect 489208 650898 524652 651134
rect 524888 650898 524972 651134
rect 525208 650898 560652 651134
rect 560888 650898 560972 651134
rect 561208 650898 570292 651134
rect 570528 650898 570612 651134
rect 570848 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 607700 651134
rect -23776 650866 607700 650898
rect -23776 641494 607700 641526
rect -23776 641258 -23744 641494
rect -23508 641258 -23424 641494
rect -23188 641258 607112 641494
rect 607348 641258 607432 641494
rect 607668 641258 607700 641494
rect -23776 641174 607700 641258
rect -23776 640938 -23744 641174
rect -23508 640938 -23424 641174
rect -23188 640938 607112 641174
rect 607348 640938 607432 641174
rect 607668 640938 607700 641174
rect -23776 640906 607700 640938
rect -23776 637774 607700 637806
rect -23776 637538 -20634 637774
rect -20398 637538 -20314 637774
rect -20078 637538 604002 637774
rect 604238 637538 604322 637774
rect 604558 637538 607700 637774
rect -23776 637454 607700 637538
rect -23776 637218 -20634 637454
rect -20398 637218 -20314 637454
rect -20078 637218 604002 637454
rect 604238 637218 604322 637454
rect 604558 637218 607700 637454
rect -23776 637186 607700 637218
rect -23776 634054 607700 634086
rect -23776 633818 -17524 634054
rect -17288 633818 -17204 634054
rect -16968 633818 600892 634054
rect 601128 633818 601212 634054
rect 601448 633818 607700 634054
rect -23776 633734 607700 633818
rect -23776 633498 -17524 633734
rect -17288 633498 -17204 633734
rect -16968 633498 600892 633734
rect 601128 633498 601212 633734
rect 601448 633498 607700 633734
rect -23776 633466 607700 633498
rect -23776 630334 607700 630366
rect -23776 630098 -14414 630334
rect -14178 630098 -14094 630334
rect -13858 630098 597782 630334
rect 598018 630098 598102 630334
rect 598338 630098 607700 630334
rect -23776 630014 607700 630098
rect -23776 629778 -14414 630014
rect -14178 629778 -14094 630014
rect -13858 629778 597782 630014
rect 598018 629778 598102 630014
rect 598338 629778 607700 630014
rect -23776 629746 607700 629778
rect -23776 626614 607700 626646
rect -23776 626378 -11304 626614
rect -11068 626378 -10984 626614
rect -10748 626378 594672 626614
rect 594908 626378 594992 626614
rect 595228 626378 607700 626614
rect -23776 626294 607700 626378
rect -23776 626058 -11304 626294
rect -11068 626058 -10984 626294
rect -10748 626058 594672 626294
rect 594908 626058 594992 626294
rect 595228 626058 607700 626294
rect -23776 626026 607700 626058
rect -23776 622894 607700 622926
rect -23776 622658 -8194 622894
rect -7958 622658 -7874 622894
rect -7638 622658 591562 622894
rect 591798 622658 591882 622894
rect 592118 622658 607700 622894
rect -23776 622574 607700 622658
rect -23776 622338 -8194 622574
rect -7958 622338 -7874 622574
rect -7638 622338 591562 622574
rect 591798 622338 591882 622574
rect 592118 622338 607700 622574
rect -23776 622306 607700 622338
rect -23776 619174 607700 619206
rect -23776 618938 -5084 619174
rect -4848 618938 -4764 619174
rect -4528 618938 7876 619174
rect 8112 618938 8196 619174
rect 8432 618938 38032 619174
rect 38268 618938 38352 619174
rect 38588 618938 74032 619174
rect 74268 618938 74352 619174
rect 74588 618938 110032 619174
rect 110268 618938 110352 619174
rect 110588 618938 146032 619174
rect 146268 618938 146352 619174
rect 146588 618938 182032 619174
rect 182268 618938 182352 619174
rect 182588 618938 218032 619174
rect 218268 618938 218352 619174
rect 218588 618938 254032 619174
rect 254268 618938 254352 619174
rect 254588 618938 290032 619174
rect 290268 618938 290352 619174
rect 290588 618938 326032 619174
rect 326268 618938 326352 619174
rect 326588 618938 362032 619174
rect 362268 618938 362352 619174
rect 362588 618938 398032 619174
rect 398268 618938 398352 619174
rect 398588 618938 434032 619174
rect 434268 618938 434352 619174
rect 434588 618938 470032 619174
rect 470268 618938 470352 619174
rect 470588 618938 506032 619174
rect 506268 618938 506352 619174
rect 506588 618938 542032 619174
rect 542268 618938 542352 619174
rect 542588 618938 571532 619174
rect 571768 618938 571852 619174
rect 572088 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 588452 619174
rect 588688 618938 588772 619174
rect 589008 618938 607700 619174
rect -23776 618854 607700 618938
rect -23776 618618 -5084 618854
rect -4848 618618 -4764 618854
rect -4528 618618 7876 618854
rect 8112 618618 8196 618854
rect 8432 618618 38032 618854
rect 38268 618618 38352 618854
rect 38588 618618 74032 618854
rect 74268 618618 74352 618854
rect 74588 618618 110032 618854
rect 110268 618618 110352 618854
rect 110588 618618 146032 618854
rect 146268 618618 146352 618854
rect 146588 618618 182032 618854
rect 182268 618618 182352 618854
rect 182588 618618 218032 618854
rect 218268 618618 218352 618854
rect 218588 618618 254032 618854
rect 254268 618618 254352 618854
rect 254588 618618 290032 618854
rect 290268 618618 290352 618854
rect 290588 618618 326032 618854
rect 326268 618618 326352 618854
rect 326588 618618 362032 618854
rect 362268 618618 362352 618854
rect 362588 618618 398032 618854
rect 398268 618618 398352 618854
rect 398588 618618 434032 618854
rect 434268 618618 434352 618854
rect 434588 618618 470032 618854
rect 470268 618618 470352 618854
rect 470588 618618 506032 618854
rect 506268 618618 506352 618854
rect 506588 618618 542032 618854
rect 542268 618618 542352 618854
rect 542588 618618 571532 618854
rect 571768 618618 571852 618854
rect 572088 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 588452 618854
rect 588688 618618 588772 618854
rect 589008 618618 607700 618854
rect -23776 618586 607700 618618
rect -23776 615454 607700 615486
rect -23776 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 9116 615454
rect 9352 615218 9436 615454
rect 9672 615218 56652 615454
rect 56888 615218 56972 615454
rect 57208 615218 92652 615454
rect 92888 615218 92972 615454
rect 93208 615218 128652 615454
rect 128888 615218 128972 615454
rect 129208 615218 164652 615454
rect 164888 615218 164972 615454
rect 165208 615218 200652 615454
rect 200888 615218 200972 615454
rect 201208 615218 236652 615454
rect 236888 615218 236972 615454
rect 237208 615218 272652 615454
rect 272888 615218 272972 615454
rect 273208 615218 308652 615454
rect 308888 615218 308972 615454
rect 309208 615218 344652 615454
rect 344888 615218 344972 615454
rect 345208 615218 380652 615454
rect 380888 615218 380972 615454
rect 381208 615218 416652 615454
rect 416888 615218 416972 615454
rect 417208 615218 452652 615454
rect 452888 615218 452972 615454
rect 453208 615218 488652 615454
rect 488888 615218 488972 615454
rect 489208 615218 524652 615454
rect 524888 615218 524972 615454
rect 525208 615218 560652 615454
rect 560888 615218 560972 615454
rect 561208 615218 570292 615454
rect 570528 615218 570612 615454
rect 570848 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 607700 615454
rect -23776 615134 607700 615218
rect -23776 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 9116 615134
rect 9352 614898 9436 615134
rect 9672 614898 56652 615134
rect 56888 614898 56972 615134
rect 57208 614898 92652 615134
rect 92888 614898 92972 615134
rect 93208 614898 128652 615134
rect 128888 614898 128972 615134
rect 129208 614898 164652 615134
rect 164888 614898 164972 615134
rect 165208 614898 200652 615134
rect 200888 614898 200972 615134
rect 201208 614898 236652 615134
rect 236888 614898 236972 615134
rect 237208 614898 272652 615134
rect 272888 614898 272972 615134
rect 273208 614898 308652 615134
rect 308888 614898 308972 615134
rect 309208 614898 344652 615134
rect 344888 614898 344972 615134
rect 345208 614898 380652 615134
rect 380888 614898 380972 615134
rect 381208 614898 416652 615134
rect 416888 614898 416972 615134
rect 417208 614898 452652 615134
rect 452888 614898 452972 615134
rect 453208 614898 488652 615134
rect 488888 614898 488972 615134
rect 489208 614898 524652 615134
rect 524888 614898 524972 615134
rect 525208 614898 560652 615134
rect 560888 614898 560972 615134
rect 561208 614898 570292 615134
rect 570528 614898 570612 615134
rect 570848 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 607700 615134
rect -23776 614866 607700 614898
rect -23776 605494 607700 605526
rect -23776 605258 -23744 605494
rect -23508 605258 -23424 605494
rect -23188 605258 607112 605494
rect 607348 605258 607432 605494
rect 607668 605258 607700 605494
rect -23776 605174 607700 605258
rect -23776 604938 -23744 605174
rect -23508 604938 -23424 605174
rect -23188 604938 607112 605174
rect 607348 604938 607432 605174
rect 607668 604938 607700 605174
rect -23776 604906 607700 604938
rect -23776 601774 607700 601806
rect -23776 601538 -20634 601774
rect -20398 601538 -20314 601774
rect -20078 601538 604002 601774
rect 604238 601538 604322 601774
rect 604558 601538 607700 601774
rect -23776 601454 607700 601538
rect -23776 601218 -20634 601454
rect -20398 601218 -20314 601454
rect -20078 601218 604002 601454
rect 604238 601218 604322 601454
rect 604558 601218 607700 601454
rect -23776 601186 607700 601218
rect -23776 598054 607700 598086
rect -23776 597818 -17524 598054
rect -17288 597818 -17204 598054
rect -16968 597818 600892 598054
rect 601128 597818 601212 598054
rect 601448 597818 607700 598054
rect -23776 597734 607700 597818
rect -23776 597498 -17524 597734
rect -17288 597498 -17204 597734
rect -16968 597498 600892 597734
rect 601128 597498 601212 597734
rect 601448 597498 607700 597734
rect -23776 597466 607700 597498
rect -23776 594334 607700 594366
rect -23776 594098 -14414 594334
rect -14178 594098 -14094 594334
rect -13858 594098 597782 594334
rect 598018 594098 598102 594334
rect 598338 594098 607700 594334
rect -23776 594014 607700 594098
rect -23776 593778 -14414 594014
rect -14178 593778 -14094 594014
rect -13858 593778 597782 594014
rect 598018 593778 598102 594014
rect 598338 593778 607700 594014
rect -23776 593746 607700 593778
rect -23776 590614 607700 590646
rect -23776 590378 -11304 590614
rect -11068 590378 -10984 590614
rect -10748 590378 594672 590614
rect 594908 590378 594992 590614
rect 595228 590378 607700 590614
rect -23776 590294 607700 590378
rect -23776 590058 -11304 590294
rect -11068 590058 -10984 590294
rect -10748 590058 594672 590294
rect 594908 590058 594992 590294
rect 595228 590058 607700 590294
rect -23776 590026 607700 590058
rect -23776 586894 607700 586926
rect -23776 586658 -8194 586894
rect -7958 586658 -7874 586894
rect -7638 586658 591562 586894
rect 591798 586658 591882 586894
rect 592118 586658 607700 586894
rect -23776 586574 607700 586658
rect -23776 586338 -8194 586574
rect -7958 586338 -7874 586574
rect -7638 586338 591562 586574
rect 591798 586338 591882 586574
rect 592118 586338 607700 586574
rect -23776 586306 607700 586338
rect -23776 583174 607700 583206
rect -23776 582938 -5084 583174
rect -4848 582938 -4764 583174
rect -4528 582938 7876 583174
rect 8112 582938 8196 583174
rect 8432 582938 38032 583174
rect 38268 582938 38352 583174
rect 38588 582938 74032 583174
rect 74268 582938 74352 583174
rect 74588 582938 110032 583174
rect 110268 582938 110352 583174
rect 110588 582938 146032 583174
rect 146268 582938 146352 583174
rect 146588 582938 182032 583174
rect 182268 582938 182352 583174
rect 182588 582938 218032 583174
rect 218268 582938 218352 583174
rect 218588 582938 254032 583174
rect 254268 582938 254352 583174
rect 254588 582938 290032 583174
rect 290268 582938 290352 583174
rect 290588 582938 326032 583174
rect 326268 582938 326352 583174
rect 326588 582938 362032 583174
rect 362268 582938 362352 583174
rect 362588 582938 398032 583174
rect 398268 582938 398352 583174
rect 398588 582938 434032 583174
rect 434268 582938 434352 583174
rect 434588 582938 470032 583174
rect 470268 582938 470352 583174
rect 470588 582938 506032 583174
rect 506268 582938 506352 583174
rect 506588 582938 542032 583174
rect 542268 582938 542352 583174
rect 542588 582938 571532 583174
rect 571768 582938 571852 583174
rect 572088 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 588452 583174
rect 588688 582938 588772 583174
rect 589008 582938 607700 583174
rect -23776 582854 607700 582938
rect -23776 582618 -5084 582854
rect -4848 582618 -4764 582854
rect -4528 582618 7876 582854
rect 8112 582618 8196 582854
rect 8432 582618 38032 582854
rect 38268 582618 38352 582854
rect 38588 582618 74032 582854
rect 74268 582618 74352 582854
rect 74588 582618 110032 582854
rect 110268 582618 110352 582854
rect 110588 582618 146032 582854
rect 146268 582618 146352 582854
rect 146588 582618 182032 582854
rect 182268 582618 182352 582854
rect 182588 582618 218032 582854
rect 218268 582618 218352 582854
rect 218588 582618 254032 582854
rect 254268 582618 254352 582854
rect 254588 582618 290032 582854
rect 290268 582618 290352 582854
rect 290588 582618 326032 582854
rect 326268 582618 326352 582854
rect 326588 582618 362032 582854
rect 362268 582618 362352 582854
rect 362588 582618 398032 582854
rect 398268 582618 398352 582854
rect 398588 582618 434032 582854
rect 434268 582618 434352 582854
rect 434588 582618 470032 582854
rect 470268 582618 470352 582854
rect 470588 582618 506032 582854
rect 506268 582618 506352 582854
rect 506588 582618 542032 582854
rect 542268 582618 542352 582854
rect 542588 582618 571532 582854
rect 571768 582618 571852 582854
rect 572088 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 588452 582854
rect 588688 582618 588772 582854
rect 589008 582618 607700 582854
rect -23776 582586 607700 582618
rect -23776 579454 607700 579486
rect -23776 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 9116 579454
rect 9352 579218 9436 579454
rect 9672 579218 56652 579454
rect 56888 579218 56972 579454
rect 57208 579218 92652 579454
rect 92888 579218 92972 579454
rect 93208 579218 128652 579454
rect 128888 579218 128972 579454
rect 129208 579218 164652 579454
rect 164888 579218 164972 579454
rect 165208 579218 200652 579454
rect 200888 579218 200972 579454
rect 201208 579218 236652 579454
rect 236888 579218 236972 579454
rect 237208 579218 272652 579454
rect 272888 579218 272972 579454
rect 273208 579218 308652 579454
rect 308888 579218 308972 579454
rect 309208 579218 344652 579454
rect 344888 579218 344972 579454
rect 345208 579218 380652 579454
rect 380888 579218 380972 579454
rect 381208 579218 416652 579454
rect 416888 579218 416972 579454
rect 417208 579218 452652 579454
rect 452888 579218 452972 579454
rect 453208 579218 488652 579454
rect 488888 579218 488972 579454
rect 489208 579218 524652 579454
rect 524888 579218 524972 579454
rect 525208 579218 560652 579454
rect 560888 579218 560972 579454
rect 561208 579218 570292 579454
rect 570528 579218 570612 579454
rect 570848 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 607700 579454
rect -23776 579134 607700 579218
rect -23776 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 9116 579134
rect 9352 578898 9436 579134
rect 9672 578898 56652 579134
rect 56888 578898 56972 579134
rect 57208 578898 92652 579134
rect 92888 578898 92972 579134
rect 93208 578898 128652 579134
rect 128888 578898 128972 579134
rect 129208 578898 164652 579134
rect 164888 578898 164972 579134
rect 165208 578898 200652 579134
rect 200888 578898 200972 579134
rect 201208 578898 236652 579134
rect 236888 578898 236972 579134
rect 237208 578898 272652 579134
rect 272888 578898 272972 579134
rect 273208 578898 308652 579134
rect 308888 578898 308972 579134
rect 309208 578898 344652 579134
rect 344888 578898 344972 579134
rect 345208 578898 380652 579134
rect 380888 578898 380972 579134
rect 381208 578898 416652 579134
rect 416888 578898 416972 579134
rect 417208 578898 452652 579134
rect 452888 578898 452972 579134
rect 453208 578898 488652 579134
rect 488888 578898 488972 579134
rect 489208 578898 524652 579134
rect 524888 578898 524972 579134
rect 525208 578898 560652 579134
rect 560888 578898 560972 579134
rect 561208 578898 570292 579134
rect 570528 578898 570612 579134
rect 570848 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 607700 579134
rect -23776 578866 607700 578898
rect -23776 569494 607700 569526
rect -23776 569258 -23744 569494
rect -23508 569258 -23424 569494
rect -23188 569258 607112 569494
rect 607348 569258 607432 569494
rect 607668 569258 607700 569494
rect -23776 569174 607700 569258
rect -23776 568938 -23744 569174
rect -23508 568938 -23424 569174
rect -23188 568938 607112 569174
rect 607348 568938 607432 569174
rect 607668 568938 607700 569174
rect -23776 568906 607700 568938
rect -23776 565774 607700 565806
rect -23776 565538 -20634 565774
rect -20398 565538 -20314 565774
rect -20078 565538 604002 565774
rect 604238 565538 604322 565774
rect 604558 565538 607700 565774
rect -23776 565454 607700 565538
rect -23776 565218 -20634 565454
rect -20398 565218 -20314 565454
rect -20078 565218 604002 565454
rect 604238 565218 604322 565454
rect 604558 565218 607700 565454
rect -23776 565186 607700 565218
rect -23776 562054 607700 562086
rect -23776 561818 -17524 562054
rect -17288 561818 -17204 562054
rect -16968 561818 600892 562054
rect 601128 561818 601212 562054
rect 601448 561818 607700 562054
rect -23776 561734 607700 561818
rect -23776 561498 -17524 561734
rect -17288 561498 -17204 561734
rect -16968 561498 600892 561734
rect 601128 561498 601212 561734
rect 601448 561498 607700 561734
rect -23776 561466 607700 561498
rect -23776 558334 607700 558366
rect -23776 558098 -14414 558334
rect -14178 558098 -14094 558334
rect -13858 558098 597782 558334
rect 598018 558098 598102 558334
rect 598338 558098 607700 558334
rect -23776 558014 607700 558098
rect -23776 557778 -14414 558014
rect -14178 557778 -14094 558014
rect -13858 557778 597782 558014
rect 598018 557778 598102 558014
rect 598338 557778 607700 558014
rect -23776 557746 607700 557778
rect -23776 554614 607700 554646
rect -23776 554378 -11304 554614
rect -11068 554378 -10984 554614
rect -10748 554378 594672 554614
rect 594908 554378 594992 554614
rect 595228 554378 607700 554614
rect -23776 554294 607700 554378
rect -23776 554058 -11304 554294
rect -11068 554058 -10984 554294
rect -10748 554058 594672 554294
rect 594908 554058 594992 554294
rect 595228 554058 607700 554294
rect -23776 554026 607700 554058
rect -23776 550894 607700 550926
rect -23776 550658 -8194 550894
rect -7958 550658 -7874 550894
rect -7638 550658 591562 550894
rect 591798 550658 591882 550894
rect 592118 550658 607700 550894
rect -23776 550574 607700 550658
rect -23776 550338 -8194 550574
rect -7958 550338 -7874 550574
rect -7638 550338 591562 550574
rect 591798 550338 591882 550574
rect 592118 550338 607700 550574
rect -23776 550306 607700 550338
rect -23776 547174 607700 547206
rect -23776 546938 -5084 547174
rect -4848 546938 -4764 547174
rect -4528 546938 7876 547174
rect 8112 546938 8196 547174
rect 8432 546938 38032 547174
rect 38268 546938 38352 547174
rect 38588 546938 74032 547174
rect 74268 546938 74352 547174
rect 74588 546938 110032 547174
rect 110268 546938 110352 547174
rect 110588 546938 146032 547174
rect 146268 546938 146352 547174
rect 146588 546938 182032 547174
rect 182268 546938 182352 547174
rect 182588 546938 218032 547174
rect 218268 546938 218352 547174
rect 218588 546938 254032 547174
rect 254268 546938 254352 547174
rect 254588 546938 290032 547174
rect 290268 546938 290352 547174
rect 290588 546938 326032 547174
rect 326268 546938 326352 547174
rect 326588 546938 362032 547174
rect 362268 546938 362352 547174
rect 362588 546938 398032 547174
rect 398268 546938 398352 547174
rect 398588 546938 434032 547174
rect 434268 546938 434352 547174
rect 434588 546938 470032 547174
rect 470268 546938 470352 547174
rect 470588 546938 506032 547174
rect 506268 546938 506352 547174
rect 506588 546938 542032 547174
rect 542268 546938 542352 547174
rect 542588 546938 571532 547174
rect 571768 546938 571852 547174
rect 572088 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 588452 547174
rect 588688 546938 588772 547174
rect 589008 546938 607700 547174
rect -23776 546854 607700 546938
rect -23776 546618 -5084 546854
rect -4848 546618 -4764 546854
rect -4528 546618 7876 546854
rect 8112 546618 8196 546854
rect 8432 546618 38032 546854
rect 38268 546618 38352 546854
rect 38588 546618 74032 546854
rect 74268 546618 74352 546854
rect 74588 546618 110032 546854
rect 110268 546618 110352 546854
rect 110588 546618 146032 546854
rect 146268 546618 146352 546854
rect 146588 546618 182032 546854
rect 182268 546618 182352 546854
rect 182588 546618 218032 546854
rect 218268 546618 218352 546854
rect 218588 546618 254032 546854
rect 254268 546618 254352 546854
rect 254588 546618 290032 546854
rect 290268 546618 290352 546854
rect 290588 546618 326032 546854
rect 326268 546618 326352 546854
rect 326588 546618 362032 546854
rect 362268 546618 362352 546854
rect 362588 546618 398032 546854
rect 398268 546618 398352 546854
rect 398588 546618 434032 546854
rect 434268 546618 434352 546854
rect 434588 546618 470032 546854
rect 470268 546618 470352 546854
rect 470588 546618 506032 546854
rect 506268 546618 506352 546854
rect 506588 546618 542032 546854
rect 542268 546618 542352 546854
rect 542588 546618 571532 546854
rect 571768 546618 571852 546854
rect 572088 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 588452 546854
rect 588688 546618 588772 546854
rect 589008 546618 607700 546854
rect -23776 546586 607700 546618
rect -23776 543454 607700 543486
rect -23776 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 9116 543454
rect 9352 543218 9436 543454
rect 9672 543218 56652 543454
rect 56888 543218 56972 543454
rect 57208 543218 92652 543454
rect 92888 543218 92972 543454
rect 93208 543218 128652 543454
rect 128888 543218 128972 543454
rect 129208 543218 164652 543454
rect 164888 543218 164972 543454
rect 165208 543218 200652 543454
rect 200888 543218 200972 543454
rect 201208 543218 236652 543454
rect 236888 543218 236972 543454
rect 237208 543218 272652 543454
rect 272888 543218 272972 543454
rect 273208 543218 308652 543454
rect 308888 543218 308972 543454
rect 309208 543218 344652 543454
rect 344888 543218 344972 543454
rect 345208 543218 380652 543454
rect 380888 543218 380972 543454
rect 381208 543218 416652 543454
rect 416888 543218 416972 543454
rect 417208 543218 452652 543454
rect 452888 543218 452972 543454
rect 453208 543218 488652 543454
rect 488888 543218 488972 543454
rect 489208 543218 524652 543454
rect 524888 543218 524972 543454
rect 525208 543218 560652 543454
rect 560888 543218 560972 543454
rect 561208 543218 570292 543454
rect 570528 543218 570612 543454
rect 570848 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 607700 543454
rect -23776 543134 607700 543218
rect -23776 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 9116 543134
rect 9352 542898 9436 543134
rect 9672 542898 56652 543134
rect 56888 542898 56972 543134
rect 57208 542898 92652 543134
rect 92888 542898 92972 543134
rect 93208 542898 128652 543134
rect 128888 542898 128972 543134
rect 129208 542898 164652 543134
rect 164888 542898 164972 543134
rect 165208 542898 200652 543134
rect 200888 542898 200972 543134
rect 201208 542898 236652 543134
rect 236888 542898 236972 543134
rect 237208 542898 272652 543134
rect 272888 542898 272972 543134
rect 273208 542898 308652 543134
rect 308888 542898 308972 543134
rect 309208 542898 344652 543134
rect 344888 542898 344972 543134
rect 345208 542898 380652 543134
rect 380888 542898 380972 543134
rect 381208 542898 416652 543134
rect 416888 542898 416972 543134
rect 417208 542898 452652 543134
rect 452888 542898 452972 543134
rect 453208 542898 488652 543134
rect 488888 542898 488972 543134
rect 489208 542898 524652 543134
rect 524888 542898 524972 543134
rect 525208 542898 560652 543134
rect 560888 542898 560972 543134
rect 561208 542898 570292 543134
rect 570528 542898 570612 543134
rect 570848 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 607700 543134
rect -23776 542866 607700 542898
rect -23776 533494 607700 533526
rect -23776 533258 -23744 533494
rect -23508 533258 -23424 533494
rect -23188 533258 607112 533494
rect 607348 533258 607432 533494
rect 607668 533258 607700 533494
rect -23776 533174 607700 533258
rect -23776 532938 -23744 533174
rect -23508 532938 -23424 533174
rect -23188 532938 607112 533174
rect 607348 532938 607432 533174
rect 607668 532938 607700 533174
rect -23776 532906 607700 532938
rect -23776 529774 607700 529806
rect -23776 529538 -20634 529774
rect -20398 529538 -20314 529774
rect -20078 529538 604002 529774
rect 604238 529538 604322 529774
rect 604558 529538 607700 529774
rect -23776 529454 607700 529538
rect -23776 529218 -20634 529454
rect -20398 529218 -20314 529454
rect -20078 529218 604002 529454
rect 604238 529218 604322 529454
rect 604558 529218 607700 529454
rect -23776 529186 607700 529218
rect -23776 526054 607700 526086
rect -23776 525818 -17524 526054
rect -17288 525818 -17204 526054
rect -16968 525818 600892 526054
rect 601128 525818 601212 526054
rect 601448 525818 607700 526054
rect -23776 525734 607700 525818
rect -23776 525498 -17524 525734
rect -17288 525498 -17204 525734
rect -16968 525498 600892 525734
rect 601128 525498 601212 525734
rect 601448 525498 607700 525734
rect -23776 525466 607700 525498
rect -23776 522334 607700 522366
rect -23776 522098 -14414 522334
rect -14178 522098 -14094 522334
rect -13858 522098 597782 522334
rect 598018 522098 598102 522334
rect 598338 522098 607700 522334
rect -23776 522014 607700 522098
rect -23776 521778 -14414 522014
rect -14178 521778 -14094 522014
rect -13858 521778 597782 522014
rect 598018 521778 598102 522014
rect 598338 521778 607700 522014
rect -23776 521746 607700 521778
rect -23776 518614 607700 518646
rect -23776 518378 -11304 518614
rect -11068 518378 -10984 518614
rect -10748 518378 594672 518614
rect 594908 518378 594992 518614
rect 595228 518378 607700 518614
rect -23776 518294 607700 518378
rect -23776 518058 -11304 518294
rect -11068 518058 -10984 518294
rect -10748 518058 594672 518294
rect 594908 518058 594992 518294
rect 595228 518058 607700 518294
rect -23776 518026 607700 518058
rect -23776 514894 607700 514926
rect -23776 514658 -8194 514894
rect -7958 514658 -7874 514894
rect -7638 514658 591562 514894
rect 591798 514658 591882 514894
rect 592118 514658 607700 514894
rect -23776 514574 607700 514658
rect -23776 514338 -8194 514574
rect -7958 514338 -7874 514574
rect -7638 514338 591562 514574
rect 591798 514338 591882 514574
rect 592118 514338 607700 514574
rect -23776 514306 607700 514338
rect -23776 511174 607700 511206
rect -23776 510938 -5084 511174
rect -4848 510938 -4764 511174
rect -4528 510938 7876 511174
rect 8112 510938 8196 511174
rect 8432 510938 38032 511174
rect 38268 510938 38352 511174
rect 38588 510938 60622 511174
rect 60858 510938 159098 511174
rect 159334 510938 182032 511174
rect 182268 510938 182352 511174
rect 182588 510938 185622 511174
rect 185858 510938 284098 511174
rect 284334 510938 290032 511174
rect 290268 510938 290352 511174
rect 290588 510938 310622 511174
rect 310858 510938 409098 511174
rect 409334 510938 434032 511174
rect 434268 510938 434352 511174
rect 434588 510938 436622 511174
rect 436858 510938 535098 511174
rect 535334 510938 542032 511174
rect 542268 510938 542352 511174
rect 542588 510938 571532 511174
rect 571768 510938 571852 511174
rect 572088 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 588452 511174
rect 588688 510938 588772 511174
rect 589008 510938 607700 511174
rect -23776 510854 607700 510938
rect -23776 510618 -5084 510854
rect -4848 510618 -4764 510854
rect -4528 510618 7876 510854
rect 8112 510618 8196 510854
rect 8432 510618 38032 510854
rect 38268 510618 38352 510854
rect 38588 510618 60622 510854
rect 60858 510618 159098 510854
rect 159334 510618 182032 510854
rect 182268 510618 182352 510854
rect 182588 510618 185622 510854
rect 185858 510618 284098 510854
rect 284334 510618 290032 510854
rect 290268 510618 290352 510854
rect 290588 510618 310622 510854
rect 310858 510618 409098 510854
rect 409334 510618 434032 510854
rect 434268 510618 434352 510854
rect 434588 510618 436622 510854
rect 436858 510618 535098 510854
rect 535334 510618 542032 510854
rect 542268 510618 542352 510854
rect 542588 510618 571532 510854
rect 571768 510618 571852 510854
rect 572088 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 588452 510854
rect 588688 510618 588772 510854
rect 589008 510618 607700 510854
rect -23776 510586 607700 510618
rect -23776 507454 607700 507486
rect -23776 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 9116 507454
rect 9352 507218 9436 507454
rect 9672 507218 56652 507454
rect 56888 507218 56972 507454
rect 57208 507218 61342 507454
rect 61578 507218 158378 507454
rect 158614 507218 164652 507454
rect 164888 507218 164972 507454
rect 165208 507218 186342 507454
rect 186578 507218 283378 507454
rect 283614 507218 308652 507454
rect 308888 507218 308972 507454
rect 309208 507218 311342 507454
rect 311578 507218 408378 507454
rect 408614 507218 416652 507454
rect 416888 507218 416972 507454
rect 417208 507218 437342 507454
rect 437578 507218 534378 507454
rect 534614 507218 560652 507454
rect 560888 507218 560972 507454
rect 561208 507218 570292 507454
rect 570528 507218 570612 507454
rect 570848 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 607700 507454
rect -23776 507134 607700 507218
rect -23776 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 9116 507134
rect 9352 506898 9436 507134
rect 9672 506898 56652 507134
rect 56888 506898 56972 507134
rect 57208 506898 61342 507134
rect 61578 506898 158378 507134
rect 158614 506898 164652 507134
rect 164888 506898 164972 507134
rect 165208 506898 186342 507134
rect 186578 506898 283378 507134
rect 283614 506898 308652 507134
rect 308888 506898 308972 507134
rect 309208 506898 311342 507134
rect 311578 506898 408378 507134
rect 408614 506898 416652 507134
rect 416888 506898 416972 507134
rect 417208 506898 437342 507134
rect 437578 506898 534378 507134
rect 534614 506898 560652 507134
rect 560888 506898 560972 507134
rect 561208 506898 570292 507134
rect 570528 506898 570612 507134
rect 570848 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 607700 507134
rect -23776 506866 607700 506898
rect -23776 497494 607700 497526
rect -23776 497258 -23744 497494
rect -23508 497258 -23424 497494
rect -23188 497258 607112 497494
rect 607348 497258 607432 497494
rect 607668 497258 607700 497494
rect -23776 497174 607700 497258
rect -23776 496938 -23744 497174
rect -23508 496938 -23424 497174
rect -23188 496938 607112 497174
rect 607348 496938 607432 497174
rect 607668 496938 607700 497174
rect -23776 496906 607700 496938
rect -23776 493774 607700 493806
rect -23776 493538 -20634 493774
rect -20398 493538 -20314 493774
rect -20078 493538 604002 493774
rect 604238 493538 604322 493774
rect 604558 493538 607700 493774
rect -23776 493454 607700 493538
rect -23776 493218 -20634 493454
rect -20398 493218 -20314 493454
rect -20078 493218 604002 493454
rect 604238 493218 604322 493454
rect 604558 493218 607700 493454
rect -23776 493186 607700 493218
rect -23776 490054 607700 490086
rect -23776 489818 -17524 490054
rect -17288 489818 -17204 490054
rect -16968 489818 600892 490054
rect 601128 489818 601212 490054
rect 601448 489818 607700 490054
rect -23776 489734 607700 489818
rect -23776 489498 -17524 489734
rect -17288 489498 -17204 489734
rect -16968 489498 600892 489734
rect 601128 489498 601212 489734
rect 601448 489498 607700 489734
rect -23776 489466 607700 489498
rect -23776 486334 607700 486366
rect -23776 486098 -14414 486334
rect -14178 486098 -14094 486334
rect -13858 486098 597782 486334
rect 598018 486098 598102 486334
rect 598338 486098 607700 486334
rect -23776 486014 607700 486098
rect -23776 485778 -14414 486014
rect -14178 485778 -14094 486014
rect -13858 485778 597782 486014
rect 598018 485778 598102 486014
rect 598338 485778 607700 486014
rect -23776 485746 607700 485778
rect -23776 482614 607700 482646
rect -23776 482378 -11304 482614
rect -11068 482378 -10984 482614
rect -10748 482378 594672 482614
rect 594908 482378 594992 482614
rect 595228 482378 607700 482614
rect -23776 482294 607700 482378
rect -23776 482058 -11304 482294
rect -11068 482058 -10984 482294
rect -10748 482058 594672 482294
rect 594908 482058 594992 482294
rect 595228 482058 607700 482294
rect -23776 482026 607700 482058
rect -23776 478894 607700 478926
rect -23776 478658 -8194 478894
rect -7958 478658 -7874 478894
rect -7638 478658 591562 478894
rect 591798 478658 591882 478894
rect 592118 478658 607700 478894
rect -23776 478574 607700 478658
rect -23776 478338 -8194 478574
rect -7958 478338 -7874 478574
rect -7638 478338 591562 478574
rect 591798 478338 591882 478574
rect 592118 478338 607700 478574
rect -23776 478306 607700 478338
rect -23776 475174 607700 475206
rect -23776 474938 -5084 475174
rect -4848 474938 -4764 475174
rect -4528 474938 7876 475174
rect 8112 474938 8196 475174
rect 8432 474938 38032 475174
rect 38268 474938 38352 475174
rect 38588 474938 60622 475174
rect 60858 474938 159098 475174
rect 159334 474938 182032 475174
rect 182268 474938 182352 475174
rect 182588 474938 185622 475174
rect 185858 474938 284098 475174
rect 284334 474938 290032 475174
rect 290268 474938 290352 475174
rect 290588 474938 310622 475174
rect 310858 474938 409098 475174
rect 409334 474938 434032 475174
rect 434268 474938 434352 475174
rect 434588 474938 436622 475174
rect 436858 474938 535098 475174
rect 535334 474938 542032 475174
rect 542268 474938 542352 475174
rect 542588 474938 571532 475174
rect 571768 474938 571852 475174
rect 572088 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 588452 475174
rect 588688 474938 588772 475174
rect 589008 474938 607700 475174
rect -23776 474854 607700 474938
rect -23776 474618 -5084 474854
rect -4848 474618 -4764 474854
rect -4528 474618 7876 474854
rect 8112 474618 8196 474854
rect 8432 474618 38032 474854
rect 38268 474618 38352 474854
rect 38588 474618 60622 474854
rect 60858 474618 159098 474854
rect 159334 474618 182032 474854
rect 182268 474618 182352 474854
rect 182588 474618 185622 474854
rect 185858 474618 284098 474854
rect 284334 474618 290032 474854
rect 290268 474618 290352 474854
rect 290588 474618 310622 474854
rect 310858 474618 409098 474854
rect 409334 474618 434032 474854
rect 434268 474618 434352 474854
rect 434588 474618 436622 474854
rect 436858 474618 535098 474854
rect 535334 474618 542032 474854
rect 542268 474618 542352 474854
rect 542588 474618 571532 474854
rect 571768 474618 571852 474854
rect 572088 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 588452 474854
rect 588688 474618 588772 474854
rect 589008 474618 607700 474854
rect -23776 474586 607700 474618
rect -23776 471454 607700 471486
rect -23776 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 9116 471454
rect 9352 471218 9436 471454
rect 9672 471218 56652 471454
rect 56888 471218 56972 471454
rect 57208 471218 61342 471454
rect 61578 471218 158378 471454
rect 158614 471218 164652 471454
rect 164888 471218 164972 471454
rect 165208 471218 186342 471454
rect 186578 471218 283378 471454
rect 283614 471218 308652 471454
rect 308888 471218 308972 471454
rect 309208 471218 311342 471454
rect 311578 471218 408378 471454
rect 408614 471218 416652 471454
rect 416888 471218 416972 471454
rect 417208 471218 437342 471454
rect 437578 471218 534378 471454
rect 534614 471218 560652 471454
rect 560888 471218 560972 471454
rect 561208 471218 570292 471454
rect 570528 471218 570612 471454
rect 570848 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 607700 471454
rect -23776 471134 607700 471218
rect -23776 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 9116 471134
rect 9352 470898 9436 471134
rect 9672 470898 56652 471134
rect 56888 470898 56972 471134
rect 57208 470898 61342 471134
rect 61578 470898 158378 471134
rect 158614 470898 164652 471134
rect 164888 470898 164972 471134
rect 165208 470898 186342 471134
rect 186578 470898 283378 471134
rect 283614 470898 308652 471134
rect 308888 470898 308972 471134
rect 309208 470898 311342 471134
rect 311578 470898 408378 471134
rect 408614 470898 416652 471134
rect 416888 470898 416972 471134
rect 417208 470898 437342 471134
rect 437578 470898 534378 471134
rect 534614 470898 560652 471134
rect 560888 470898 560972 471134
rect 561208 470898 570292 471134
rect 570528 470898 570612 471134
rect 570848 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 607700 471134
rect -23776 470866 607700 470898
rect -23776 461494 607700 461526
rect -23776 461258 -23744 461494
rect -23508 461258 -23424 461494
rect -23188 461258 607112 461494
rect 607348 461258 607432 461494
rect 607668 461258 607700 461494
rect -23776 461174 607700 461258
rect -23776 460938 -23744 461174
rect -23508 460938 -23424 461174
rect -23188 460938 607112 461174
rect 607348 460938 607432 461174
rect 607668 460938 607700 461174
rect -23776 460906 607700 460938
rect -23776 457774 607700 457806
rect -23776 457538 -20634 457774
rect -20398 457538 -20314 457774
rect -20078 457538 604002 457774
rect 604238 457538 604322 457774
rect 604558 457538 607700 457774
rect -23776 457454 607700 457538
rect -23776 457218 -20634 457454
rect -20398 457218 -20314 457454
rect -20078 457218 604002 457454
rect 604238 457218 604322 457454
rect 604558 457218 607700 457454
rect -23776 457186 607700 457218
rect -23776 454054 607700 454086
rect -23776 453818 -17524 454054
rect -17288 453818 -17204 454054
rect -16968 453818 600892 454054
rect 601128 453818 601212 454054
rect 601448 453818 607700 454054
rect -23776 453734 607700 453818
rect -23776 453498 -17524 453734
rect -17288 453498 -17204 453734
rect -16968 453498 600892 453734
rect 601128 453498 601212 453734
rect 601448 453498 607700 453734
rect -23776 453466 607700 453498
rect -23776 450334 607700 450366
rect -23776 450098 -14414 450334
rect -14178 450098 -14094 450334
rect -13858 450098 597782 450334
rect 598018 450098 598102 450334
rect 598338 450098 607700 450334
rect -23776 450014 607700 450098
rect -23776 449778 -14414 450014
rect -14178 449778 -14094 450014
rect -13858 449778 597782 450014
rect 598018 449778 598102 450014
rect 598338 449778 607700 450014
rect -23776 449746 607700 449778
rect -23776 446614 607700 446646
rect -23776 446378 -11304 446614
rect -11068 446378 -10984 446614
rect -10748 446378 594672 446614
rect 594908 446378 594992 446614
rect 595228 446378 607700 446614
rect -23776 446294 607700 446378
rect -23776 446058 -11304 446294
rect -11068 446058 -10984 446294
rect -10748 446058 594672 446294
rect 594908 446058 594992 446294
rect 595228 446058 607700 446294
rect -23776 446026 607700 446058
rect -23776 442894 607700 442926
rect -23776 442658 -8194 442894
rect -7958 442658 -7874 442894
rect -7638 442658 591562 442894
rect 591798 442658 591882 442894
rect 592118 442658 607700 442894
rect -23776 442574 607700 442658
rect -23776 442338 -8194 442574
rect -7958 442338 -7874 442574
rect -7638 442338 591562 442574
rect 591798 442338 591882 442574
rect 592118 442338 607700 442574
rect -23776 442306 607700 442338
rect -23776 439174 607700 439206
rect -23776 438938 -5084 439174
rect -4848 438938 -4764 439174
rect -4528 438938 7876 439174
rect 8112 438938 8196 439174
rect 8432 438938 38032 439174
rect 38268 438938 38352 439174
rect 38588 438938 60622 439174
rect 60858 438938 159098 439174
rect 159334 438938 182032 439174
rect 182268 438938 182352 439174
rect 182588 438938 185622 439174
rect 185858 438938 284098 439174
rect 284334 438938 290032 439174
rect 290268 438938 290352 439174
rect 290588 438938 310622 439174
rect 310858 438938 409098 439174
rect 409334 438938 434032 439174
rect 434268 438938 434352 439174
rect 434588 438938 436622 439174
rect 436858 438938 535098 439174
rect 535334 438938 542032 439174
rect 542268 438938 542352 439174
rect 542588 438938 571532 439174
rect 571768 438938 571852 439174
rect 572088 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 588452 439174
rect 588688 438938 588772 439174
rect 589008 438938 607700 439174
rect -23776 438854 607700 438938
rect -23776 438618 -5084 438854
rect -4848 438618 -4764 438854
rect -4528 438618 7876 438854
rect 8112 438618 8196 438854
rect 8432 438618 38032 438854
rect 38268 438618 38352 438854
rect 38588 438618 60622 438854
rect 60858 438618 159098 438854
rect 159334 438618 182032 438854
rect 182268 438618 182352 438854
rect 182588 438618 185622 438854
rect 185858 438618 284098 438854
rect 284334 438618 290032 438854
rect 290268 438618 290352 438854
rect 290588 438618 310622 438854
rect 310858 438618 409098 438854
rect 409334 438618 434032 438854
rect 434268 438618 434352 438854
rect 434588 438618 436622 438854
rect 436858 438618 535098 438854
rect 535334 438618 542032 438854
rect 542268 438618 542352 438854
rect 542588 438618 571532 438854
rect 571768 438618 571852 438854
rect 572088 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 588452 438854
rect 588688 438618 588772 438854
rect 589008 438618 607700 438854
rect -23776 438586 607700 438618
rect -23776 435454 607700 435486
rect -23776 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 9116 435454
rect 9352 435218 9436 435454
rect 9672 435218 56652 435454
rect 56888 435218 56972 435454
rect 57208 435218 61342 435454
rect 61578 435218 158378 435454
rect 158614 435218 164652 435454
rect 164888 435218 164972 435454
rect 165208 435218 186342 435454
rect 186578 435218 283378 435454
rect 283614 435218 308652 435454
rect 308888 435218 308972 435454
rect 309208 435218 311342 435454
rect 311578 435218 408378 435454
rect 408614 435218 416652 435454
rect 416888 435218 416972 435454
rect 417208 435218 437342 435454
rect 437578 435218 534378 435454
rect 534614 435218 560652 435454
rect 560888 435218 560972 435454
rect 561208 435218 570292 435454
rect 570528 435218 570612 435454
rect 570848 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 607700 435454
rect -23776 435134 607700 435218
rect -23776 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 9116 435134
rect 9352 434898 9436 435134
rect 9672 434898 56652 435134
rect 56888 434898 56972 435134
rect 57208 434898 61342 435134
rect 61578 434898 158378 435134
rect 158614 434898 164652 435134
rect 164888 434898 164972 435134
rect 165208 434898 186342 435134
rect 186578 434898 283378 435134
rect 283614 434898 308652 435134
rect 308888 434898 308972 435134
rect 309208 434898 311342 435134
rect 311578 434898 408378 435134
rect 408614 434898 416652 435134
rect 416888 434898 416972 435134
rect 417208 434898 437342 435134
rect 437578 434898 534378 435134
rect 534614 434898 560652 435134
rect 560888 434898 560972 435134
rect 561208 434898 570292 435134
rect 570528 434898 570612 435134
rect 570848 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 607700 435134
rect -23776 434866 607700 434898
rect 61280 433244 61640 433300
rect 61280 433008 61342 433244
rect 61578 433008 61640 433244
rect 61280 432952 61640 433008
rect 62952 433244 63300 433300
rect 62952 433008 63008 433244
rect 63244 433008 63300 433244
rect 62952 432952 63300 433008
rect 281656 433244 282004 433300
rect 281656 433008 281712 433244
rect 281948 433008 282004 433244
rect 281656 432952 282004 433008
rect 283316 433244 283676 433300
rect 283316 433008 283378 433244
rect 283614 433008 283676 433244
rect 283316 432952 283676 433008
rect 311280 433244 311640 433300
rect 311280 433008 311342 433244
rect 311578 433008 311640 433244
rect 311280 432952 311640 433008
rect 312952 433244 313300 433300
rect 312952 433008 313008 433244
rect 313244 433008 313300 433244
rect 312952 432952 313300 433008
rect 532656 433244 533004 433300
rect 532656 433008 532712 433244
rect 532948 433008 533004 433244
rect 532656 432952 533004 433008
rect 534316 433244 534676 433300
rect 534316 433008 534378 433244
rect 534614 433008 534676 433244
rect 534316 432952 534676 433008
rect 157336 432564 157684 432620
rect 157336 432328 157392 432564
rect 157628 432328 157684 432564
rect 157336 432272 157684 432328
rect 159036 432564 159396 432620
rect 159036 432328 159098 432564
rect 159334 432328 159396 432564
rect 159036 432272 159396 432328
rect 185560 432564 185920 432620
rect 185560 432328 185622 432564
rect 185858 432328 185920 432564
rect 185560 432272 185920 432328
rect 187272 432564 187620 432620
rect 187272 432328 187328 432564
rect 187564 432328 187620 432564
rect 187272 432272 187620 432328
rect 407336 432564 407684 432620
rect 407336 432328 407392 432564
rect 407628 432328 407684 432564
rect 407336 432272 407684 432328
rect 409036 432564 409396 432620
rect 409036 432328 409098 432564
rect 409334 432328 409396 432564
rect 409036 432272 409396 432328
rect 436560 432564 436920 432620
rect 436560 432328 436622 432564
rect 436858 432328 436920 432564
rect 436560 432272 436920 432328
rect 438272 432564 438620 432620
rect 438272 432328 438328 432564
rect 438564 432328 438620 432564
rect 438272 432272 438620 432328
rect -23776 425494 607700 425526
rect -23776 425258 -23744 425494
rect -23508 425258 -23424 425494
rect -23188 425258 607112 425494
rect 607348 425258 607432 425494
rect 607668 425258 607700 425494
rect -23776 425174 607700 425258
rect -23776 424938 -23744 425174
rect -23508 424938 -23424 425174
rect -23188 424938 607112 425174
rect 607348 424938 607432 425174
rect 607668 424938 607700 425174
rect -23776 424906 607700 424938
rect -23776 421774 607700 421806
rect -23776 421538 -20634 421774
rect -20398 421538 -20314 421774
rect -20078 421538 604002 421774
rect 604238 421538 604322 421774
rect 604558 421538 607700 421774
rect -23776 421454 607700 421538
rect -23776 421218 -20634 421454
rect -20398 421218 -20314 421454
rect -20078 421218 604002 421454
rect 604238 421218 604322 421454
rect 604558 421218 607700 421454
rect -23776 421186 607700 421218
rect -23776 418054 607700 418086
rect -23776 417818 -17524 418054
rect -17288 417818 -17204 418054
rect -16968 417818 600892 418054
rect 601128 417818 601212 418054
rect 601448 417818 607700 418054
rect -23776 417734 607700 417818
rect -23776 417498 -17524 417734
rect -17288 417498 -17204 417734
rect -16968 417498 600892 417734
rect 601128 417498 601212 417734
rect 601448 417498 607700 417734
rect -23776 417466 607700 417498
rect -23776 414334 607700 414366
rect -23776 414098 -14414 414334
rect -14178 414098 -14094 414334
rect -13858 414098 597782 414334
rect 598018 414098 598102 414334
rect 598338 414098 607700 414334
rect -23776 414014 607700 414098
rect -23776 413778 -14414 414014
rect -14178 413778 -14094 414014
rect -13858 413778 597782 414014
rect 598018 413778 598102 414014
rect 598338 413778 607700 414014
rect -23776 413746 607700 413778
rect -23776 410614 607700 410646
rect -23776 410378 -11304 410614
rect -11068 410378 -10984 410614
rect -10748 410378 594672 410614
rect 594908 410378 594992 410614
rect 595228 410378 607700 410614
rect -23776 410294 607700 410378
rect -23776 410058 -11304 410294
rect -11068 410058 -10984 410294
rect -10748 410058 594672 410294
rect 594908 410058 594992 410294
rect 595228 410058 607700 410294
rect -23776 410026 607700 410058
rect -23776 406894 607700 406926
rect -23776 406658 -8194 406894
rect -7958 406658 -7874 406894
rect -7638 406658 591562 406894
rect 591798 406658 591882 406894
rect 592118 406658 607700 406894
rect -23776 406574 607700 406658
rect -23776 406338 -8194 406574
rect -7958 406338 -7874 406574
rect -7638 406338 591562 406574
rect 591798 406338 591882 406574
rect 592118 406338 607700 406574
rect -23776 406306 607700 406338
rect -23776 403174 607700 403206
rect -23776 402938 -5084 403174
rect -4848 402938 -4764 403174
rect -4528 402938 7876 403174
rect 8112 402938 8196 403174
rect 8432 402938 38032 403174
rect 38268 402938 38352 403174
rect 38588 402938 74032 403174
rect 74268 402938 74352 403174
rect 74588 402938 110032 403174
rect 110268 402938 110352 403174
rect 110588 402938 146032 403174
rect 146268 402938 146352 403174
rect 146588 402938 182032 403174
rect 182268 402938 182352 403174
rect 182588 402938 218032 403174
rect 218268 402938 218352 403174
rect 218588 402938 254032 403174
rect 254268 402938 254352 403174
rect 254588 402938 290032 403174
rect 290268 402938 290352 403174
rect 290588 402938 326032 403174
rect 326268 402938 326352 403174
rect 326588 402938 362032 403174
rect 362268 402938 362352 403174
rect 362588 402938 398032 403174
rect 398268 402938 398352 403174
rect 398588 402938 434032 403174
rect 434268 402938 434352 403174
rect 434588 402938 470032 403174
rect 470268 402938 470352 403174
rect 470588 402938 506032 403174
rect 506268 402938 506352 403174
rect 506588 402938 542032 403174
rect 542268 402938 542352 403174
rect 542588 402938 571532 403174
rect 571768 402938 571852 403174
rect 572088 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 588452 403174
rect 588688 402938 588772 403174
rect 589008 402938 607700 403174
rect -23776 402854 607700 402938
rect -23776 402618 -5084 402854
rect -4848 402618 -4764 402854
rect -4528 402618 7876 402854
rect 8112 402618 8196 402854
rect 8432 402618 38032 402854
rect 38268 402618 38352 402854
rect 38588 402618 74032 402854
rect 74268 402618 74352 402854
rect 74588 402618 110032 402854
rect 110268 402618 110352 402854
rect 110588 402618 146032 402854
rect 146268 402618 146352 402854
rect 146588 402618 182032 402854
rect 182268 402618 182352 402854
rect 182588 402618 218032 402854
rect 218268 402618 218352 402854
rect 218588 402618 254032 402854
rect 254268 402618 254352 402854
rect 254588 402618 290032 402854
rect 290268 402618 290352 402854
rect 290588 402618 326032 402854
rect 326268 402618 326352 402854
rect 326588 402618 362032 402854
rect 362268 402618 362352 402854
rect 362588 402618 398032 402854
rect 398268 402618 398352 402854
rect 398588 402618 434032 402854
rect 434268 402618 434352 402854
rect 434588 402618 470032 402854
rect 470268 402618 470352 402854
rect 470588 402618 506032 402854
rect 506268 402618 506352 402854
rect 506588 402618 542032 402854
rect 542268 402618 542352 402854
rect 542588 402618 571532 402854
rect 571768 402618 571852 402854
rect 572088 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 588452 402854
rect 588688 402618 588772 402854
rect 589008 402618 607700 402854
rect -23776 402586 607700 402618
rect -23776 399454 607700 399486
rect -23776 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 9116 399454
rect 9352 399218 9436 399454
rect 9672 399218 56652 399454
rect 56888 399218 56972 399454
rect 57208 399218 92652 399454
rect 92888 399218 92972 399454
rect 93208 399218 128652 399454
rect 128888 399218 128972 399454
rect 129208 399218 164652 399454
rect 164888 399218 164972 399454
rect 165208 399218 200652 399454
rect 200888 399218 200972 399454
rect 201208 399218 236652 399454
rect 236888 399218 236972 399454
rect 237208 399218 272652 399454
rect 272888 399218 272972 399454
rect 273208 399218 308652 399454
rect 308888 399218 308972 399454
rect 309208 399218 344652 399454
rect 344888 399218 344972 399454
rect 345208 399218 380652 399454
rect 380888 399218 380972 399454
rect 381208 399218 416652 399454
rect 416888 399218 416972 399454
rect 417208 399218 452652 399454
rect 452888 399218 452972 399454
rect 453208 399218 488652 399454
rect 488888 399218 488972 399454
rect 489208 399218 524652 399454
rect 524888 399218 524972 399454
rect 525208 399218 560652 399454
rect 560888 399218 560972 399454
rect 561208 399218 570292 399454
rect 570528 399218 570612 399454
rect 570848 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 607700 399454
rect -23776 399134 607700 399218
rect -23776 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 9116 399134
rect 9352 398898 9436 399134
rect 9672 398898 56652 399134
rect 56888 398898 56972 399134
rect 57208 398898 92652 399134
rect 92888 398898 92972 399134
rect 93208 398898 128652 399134
rect 128888 398898 128972 399134
rect 129208 398898 164652 399134
rect 164888 398898 164972 399134
rect 165208 398898 200652 399134
rect 200888 398898 200972 399134
rect 201208 398898 236652 399134
rect 236888 398898 236972 399134
rect 237208 398898 272652 399134
rect 272888 398898 272972 399134
rect 273208 398898 308652 399134
rect 308888 398898 308972 399134
rect 309208 398898 344652 399134
rect 344888 398898 344972 399134
rect 345208 398898 380652 399134
rect 380888 398898 380972 399134
rect 381208 398898 416652 399134
rect 416888 398898 416972 399134
rect 417208 398898 452652 399134
rect 452888 398898 452972 399134
rect 453208 398898 488652 399134
rect 488888 398898 488972 399134
rect 489208 398898 524652 399134
rect 524888 398898 524972 399134
rect 525208 398898 560652 399134
rect 560888 398898 560972 399134
rect 561208 398898 570292 399134
rect 570528 398898 570612 399134
rect 570848 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 607700 399134
rect -23776 398866 607700 398898
rect -23776 389494 607700 389526
rect -23776 389258 -23744 389494
rect -23508 389258 -23424 389494
rect -23188 389258 607112 389494
rect 607348 389258 607432 389494
rect 607668 389258 607700 389494
rect -23776 389174 607700 389258
rect -23776 388938 -23744 389174
rect -23508 388938 -23424 389174
rect -23188 388938 607112 389174
rect 607348 388938 607432 389174
rect 607668 388938 607700 389174
rect -23776 388906 607700 388938
rect -23776 385774 607700 385806
rect -23776 385538 -20634 385774
rect -20398 385538 -20314 385774
rect -20078 385538 604002 385774
rect 604238 385538 604322 385774
rect 604558 385538 607700 385774
rect -23776 385454 607700 385538
rect -23776 385218 -20634 385454
rect -20398 385218 -20314 385454
rect -20078 385218 604002 385454
rect 604238 385218 604322 385454
rect 604558 385218 607700 385454
rect -23776 385186 607700 385218
rect -23776 382054 607700 382086
rect -23776 381818 -17524 382054
rect -17288 381818 -17204 382054
rect -16968 381818 600892 382054
rect 601128 381818 601212 382054
rect 601448 381818 607700 382054
rect -23776 381734 607700 381818
rect -23776 381498 -17524 381734
rect -17288 381498 -17204 381734
rect -16968 381498 600892 381734
rect 601128 381498 601212 381734
rect 601448 381498 607700 381734
rect -23776 381466 607700 381498
rect -23776 378334 607700 378366
rect -23776 378098 -14414 378334
rect -14178 378098 -14094 378334
rect -13858 378098 597782 378334
rect 598018 378098 598102 378334
rect 598338 378098 607700 378334
rect -23776 378014 607700 378098
rect -23776 377778 -14414 378014
rect -14178 377778 -14094 378014
rect -13858 377778 597782 378014
rect 598018 377778 598102 378014
rect 598338 377778 607700 378014
rect -23776 377746 607700 377778
rect -23776 374614 607700 374646
rect -23776 374378 -11304 374614
rect -11068 374378 -10984 374614
rect -10748 374378 594672 374614
rect 594908 374378 594992 374614
rect 595228 374378 607700 374614
rect -23776 374294 607700 374378
rect -23776 374058 -11304 374294
rect -11068 374058 -10984 374294
rect -10748 374058 594672 374294
rect 594908 374058 594992 374294
rect 595228 374058 607700 374294
rect -23776 374026 607700 374058
rect -23776 370894 607700 370926
rect -23776 370658 -8194 370894
rect -7958 370658 -7874 370894
rect -7638 370658 591562 370894
rect 591798 370658 591882 370894
rect 592118 370658 607700 370894
rect -23776 370574 607700 370658
rect -23776 370338 -8194 370574
rect -7958 370338 -7874 370574
rect -7638 370338 591562 370574
rect 591798 370338 591882 370574
rect 592118 370338 607700 370574
rect -23776 370306 607700 370338
rect -23776 367174 607700 367206
rect -23776 366938 -5084 367174
rect -4848 366938 -4764 367174
rect -4528 366938 7876 367174
rect 8112 366938 8196 367174
rect 8432 366938 38032 367174
rect 38268 366938 38352 367174
rect 38588 366938 74032 367174
rect 74268 366938 74352 367174
rect 74588 366938 110032 367174
rect 110268 366938 110352 367174
rect 110588 366938 146032 367174
rect 146268 366938 146352 367174
rect 146588 366938 182032 367174
rect 182268 366938 182352 367174
rect 182588 366938 218032 367174
rect 218268 366938 218352 367174
rect 218588 366938 254032 367174
rect 254268 366938 254352 367174
rect 254588 366938 290032 367174
rect 290268 366938 290352 367174
rect 290588 366938 326032 367174
rect 326268 366938 326352 367174
rect 326588 366938 362032 367174
rect 362268 366938 362352 367174
rect 362588 366938 398032 367174
rect 398268 366938 398352 367174
rect 398588 366938 434032 367174
rect 434268 366938 434352 367174
rect 434588 366938 470032 367174
rect 470268 366938 470352 367174
rect 470588 366938 506032 367174
rect 506268 366938 506352 367174
rect 506588 366938 542032 367174
rect 542268 366938 542352 367174
rect 542588 366938 571532 367174
rect 571768 366938 571852 367174
rect 572088 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 588452 367174
rect 588688 366938 588772 367174
rect 589008 366938 607700 367174
rect -23776 366854 607700 366938
rect -23776 366618 -5084 366854
rect -4848 366618 -4764 366854
rect -4528 366618 7876 366854
rect 8112 366618 8196 366854
rect 8432 366618 38032 366854
rect 38268 366618 38352 366854
rect 38588 366618 74032 366854
rect 74268 366618 74352 366854
rect 74588 366618 110032 366854
rect 110268 366618 110352 366854
rect 110588 366618 146032 366854
rect 146268 366618 146352 366854
rect 146588 366618 182032 366854
rect 182268 366618 182352 366854
rect 182588 366618 218032 366854
rect 218268 366618 218352 366854
rect 218588 366618 254032 366854
rect 254268 366618 254352 366854
rect 254588 366618 290032 366854
rect 290268 366618 290352 366854
rect 290588 366618 326032 366854
rect 326268 366618 326352 366854
rect 326588 366618 362032 366854
rect 362268 366618 362352 366854
rect 362588 366618 398032 366854
rect 398268 366618 398352 366854
rect 398588 366618 434032 366854
rect 434268 366618 434352 366854
rect 434588 366618 470032 366854
rect 470268 366618 470352 366854
rect 470588 366618 506032 366854
rect 506268 366618 506352 366854
rect 506588 366618 542032 366854
rect 542268 366618 542352 366854
rect 542588 366618 571532 366854
rect 571768 366618 571852 366854
rect 572088 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 588452 366854
rect 588688 366618 588772 366854
rect 589008 366618 607700 366854
rect -23776 366586 607700 366618
rect -23776 363454 607700 363486
rect -23776 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 9116 363454
rect 9352 363218 9436 363454
rect 9672 363218 56652 363454
rect 56888 363218 56972 363454
rect 57208 363218 92652 363454
rect 92888 363218 92972 363454
rect 93208 363218 128652 363454
rect 128888 363218 128972 363454
rect 129208 363218 164652 363454
rect 164888 363218 164972 363454
rect 165208 363218 200652 363454
rect 200888 363218 200972 363454
rect 201208 363218 236652 363454
rect 236888 363218 236972 363454
rect 237208 363218 272652 363454
rect 272888 363218 272972 363454
rect 273208 363218 308652 363454
rect 308888 363218 308972 363454
rect 309208 363218 344652 363454
rect 344888 363218 344972 363454
rect 345208 363218 380652 363454
rect 380888 363218 380972 363454
rect 381208 363218 416652 363454
rect 416888 363218 416972 363454
rect 417208 363218 452652 363454
rect 452888 363218 452972 363454
rect 453208 363218 488652 363454
rect 488888 363218 488972 363454
rect 489208 363218 524652 363454
rect 524888 363218 524972 363454
rect 525208 363218 560652 363454
rect 560888 363218 560972 363454
rect 561208 363218 570292 363454
rect 570528 363218 570612 363454
rect 570848 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 607700 363454
rect -23776 363134 607700 363218
rect -23776 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 9116 363134
rect 9352 362898 9436 363134
rect 9672 362898 56652 363134
rect 56888 362898 56972 363134
rect 57208 362898 92652 363134
rect 92888 362898 92972 363134
rect 93208 362898 128652 363134
rect 128888 362898 128972 363134
rect 129208 362898 164652 363134
rect 164888 362898 164972 363134
rect 165208 362898 200652 363134
rect 200888 362898 200972 363134
rect 201208 362898 236652 363134
rect 236888 362898 236972 363134
rect 237208 362898 272652 363134
rect 272888 362898 272972 363134
rect 273208 362898 308652 363134
rect 308888 362898 308972 363134
rect 309208 362898 344652 363134
rect 344888 362898 344972 363134
rect 345208 362898 380652 363134
rect 380888 362898 380972 363134
rect 381208 362898 416652 363134
rect 416888 362898 416972 363134
rect 417208 362898 452652 363134
rect 452888 362898 452972 363134
rect 453208 362898 488652 363134
rect 488888 362898 488972 363134
rect 489208 362898 524652 363134
rect 524888 362898 524972 363134
rect 525208 362898 560652 363134
rect 560888 362898 560972 363134
rect 561208 362898 570292 363134
rect 570528 362898 570612 363134
rect 570848 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 607700 363134
rect -23776 362866 607700 362898
rect -23776 353494 607700 353526
rect -23776 353258 -23744 353494
rect -23508 353258 -23424 353494
rect -23188 353258 607112 353494
rect 607348 353258 607432 353494
rect 607668 353258 607700 353494
rect -23776 353174 607700 353258
rect -23776 352938 -23744 353174
rect -23508 352938 -23424 353174
rect -23188 352938 607112 353174
rect 607348 352938 607432 353174
rect 607668 352938 607700 353174
rect -23776 352906 607700 352938
rect -23776 349774 607700 349806
rect -23776 349538 -20634 349774
rect -20398 349538 -20314 349774
rect -20078 349538 604002 349774
rect 604238 349538 604322 349774
rect 604558 349538 607700 349774
rect -23776 349454 607700 349538
rect -23776 349218 -20634 349454
rect -20398 349218 -20314 349454
rect -20078 349218 604002 349454
rect 604238 349218 604322 349454
rect 604558 349218 607700 349454
rect -23776 349186 607700 349218
rect -23776 346054 607700 346086
rect -23776 345818 -17524 346054
rect -17288 345818 -17204 346054
rect -16968 345818 600892 346054
rect 601128 345818 601212 346054
rect 601448 345818 607700 346054
rect -23776 345734 607700 345818
rect -23776 345498 -17524 345734
rect -17288 345498 -17204 345734
rect -16968 345498 600892 345734
rect 601128 345498 601212 345734
rect 601448 345498 607700 345734
rect -23776 345466 607700 345498
rect -23776 342334 607700 342366
rect -23776 342098 -14414 342334
rect -14178 342098 -14094 342334
rect -13858 342098 597782 342334
rect 598018 342098 598102 342334
rect 598338 342098 607700 342334
rect -23776 342014 607700 342098
rect -23776 341778 -14414 342014
rect -14178 341778 -14094 342014
rect -13858 341778 597782 342014
rect 598018 341778 598102 342014
rect 598338 341778 607700 342014
rect -23776 341746 607700 341778
rect -23776 338614 607700 338646
rect -23776 338378 -11304 338614
rect -11068 338378 -10984 338614
rect -10748 338378 594672 338614
rect 594908 338378 594992 338614
rect 595228 338378 607700 338614
rect -23776 338294 607700 338378
rect -23776 338058 -11304 338294
rect -11068 338058 -10984 338294
rect -10748 338058 594672 338294
rect 594908 338058 594992 338294
rect 595228 338058 607700 338294
rect -23776 338026 607700 338058
rect -23776 334894 607700 334926
rect -23776 334658 -8194 334894
rect -7958 334658 -7874 334894
rect -7638 334658 591562 334894
rect 591798 334658 591882 334894
rect 592118 334658 607700 334894
rect -23776 334574 607700 334658
rect -23776 334338 -8194 334574
rect -7958 334338 -7874 334574
rect -7638 334338 591562 334574
rect 591798 334338 591882 334574
rect 592118 334338 607700 334574
rect -23776 334306 607700 334338
rect -23776 331174 607700 331206
rect -23776 330938 -5084 331174
rect -4848 330938 -4764 331174
rect -4528 330938 7876 331174
rect 8112 330938 8196 331174
rect 8432 330938 38032 331174
rect 38268 330938 38352 331174
rect 38588 330938 74032 331174
rect 74268 330938 74352 331174
rect 74588 330938 110032 331174
rect 110268 330938 110352 331174
rect 110588 330938 146032 331174
rect 146268 330938 146352 331174
rect 146588 330938 182032 331174
rect 182268 330938 182352 331174
rect 182588 330938 218032 331174
rect 218268 330938 218352 331174
rect 218588 330938 254032 331174
rect 254268 330938 254352 331174
rect 254588 330938 290032 331174
rect 290268 330938 290352 331174
rect 290588 330938 326032 331174
rect 326268 330938 326352 331174
rect 326588 330938 362032 331174
rect 362268 330938 362352 331174
rect 362588 330938 398032 331174
rect 398268 330938 398352 331174
rect 398588 330938 434032 331174
rect 434268 330938 434352 331174
rect 434588 330938 470032 331174
rect 470268 330938 470352 331174
rect 470588 330938 506032 331174
rect 506268 330938 506352 331174
rect 506588 330938 542032 331174
rect 542268 330938 542352 331174
rect 542588 330938 571532 331174
rect 571768 330938 571852 331174
rect 572088 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 588452 331174
rect 588688 330938 588772 331174
rect 589008 330938 607700 331174
rect -23776 330854 607700 330938
rect -23776 330618 -5084 330854
rect -4848 330618 -4764 330854
rect -4528 330618 7876 330854
rect 8112 330618 8196 330854
rect 8432 330618 38032 330854
rect 38268 330618 38352 330854
rect 38588 330618 74032 330854
rect 74268 330618 74352 330854
rect 74588 330618 110032 330854
rect 110268 330618 110352 330854
rect 110588 330618 146032 330854
rect 146268 330618 146352 330854
rect 146588 330618 182032 330854
rect 182268 330618 182352 330854
rect 182588 330618 218032 330854
rect 218268 330618 218352 330854
rect 218588 330618 254032 330854
rect 254268 330618 254352 330854
rect 254588 330618 290032 330854
rect 290268 330618 290352 330854
rect 290588 330618 326032 330854
rect 326268 330618 326352 330854
rect 326588 330618 362032 330854
rect 362268 330618 362352 330854
rect 362588 330618 398032 330854
rect 398268 330618 398352 330854
rect 398588 330618 434032 330854
rect 434268 330618 434352 330854
rect 434588 330618 470032 330854
rect 470268 330618 470352 330854
rect 470588 330618 506032 330854
rect 506268 330618 506352 330854
rect 506588 330618 542032 330854
rect 542268 330618 542352 330854
rect 542588 330618 571532 330854
rect 571768 330618 571852 330854
rect 572088 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 588452 330854
rect 588688 330618 588772 330854
rect 589008 330618 607700 330854
rect -23776 330586 607700 330618
rect -23776 327454 607700 327486
rect -23776 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 9116 327454
rect 9352 327218 9436 327454
rect 9672 327218 56652 327454
rect 56888 327218 56972 327454
rect 57208 327218 92652 327454
rect 92888 327218 92972 327454
rect 93208 327218 128652 327454
rect 128888 327218 128972 327454
rect 129208 327218 164652 327454
rect 164888 327218 164972 327454
rect 165208 327218 200652 327454
rect 200888 327218 200972 327454
rect 201208 327218 236652 327454
rect 236888 327218 236972 327454
rect 237208 327218 272652 327454
rect 272888 327218 272972 327454
rect 273208 327218 308652 327454
rect 308888 327218 308972 327454
rect 309208 327218 344652 327454
rect 344888 327218 344972 327454
rect 345208 327218 380652 327454
rect 380888 327218 380972 327454
rect 381208 327218 416652 327454
rect 416888 327218 416972 327454
rect 417208 327218 452652 327454
rect 452888 327218 452972 327454
rect 453208 327218 488652 327454
rect 488888 327218 488972 327454
rect 489208 327218 524652 327454
rect 524888 327218 524972 327454
rect 525208 327218 560652 327454
rect 560888 327218 560972 327454
rect 561208 327218 570292 327454
rect 570528 327218 570612 327454
rect 570848 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 607700 327454
rect -23776 327134 607700 327218
rect -23776 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 9116 327134
rect 9352 326898 9436 327134
rect 9672 326898 56652 327134
rect 56888 326898 56972 327134
rect 57208 326898 92652 327134
rect 92888 326898 92972 327134
rect 93208 326898 128652 327134
rect 128888 326898 128972 327134
rect 129208 326898 164652 327134
rect 164888 326898 164972 327134
rect 165208 326898 200652 327134
rect 200888 326898 200972 327134
rect 201208 326898 236652 327134
rect 236888 326898 236972 327134
rect 237208 326898 272652 327134
rect 272888 326898 272972 327134
rect 273208 326898 308652 327134
rect 308888 326898 308972 327134
rect 309208 326898 344652 327134
rect 344888 326898 344972 327134
rect 345208 326898 380652 327134
rect 380888 326898 380972 327134
rect 381208 326898 416652 327134
rect 416888 326898 416972 327134
rect 417208 326898 452652 327134
rect 452888 326898 452972 327134
rect 453208 326898 488652 327134
rect 488888 326898 488972 327134
rect 489208 326898 524652 327134
rect 524888 326898 524972 327134
rect 525208 326898 560652 327134
rect 560888 326898 560972 327134
rect 561208 326898 570292 327134
rect 570528 326898 570612 327134
rect 570848 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 607700 327134
rect -23776 326866 607700 326898
rect -23776 317494 607700 317526
rect -23776 317258 -23744 317494
rect -23508 317258 -23424 317494
rect -23188 317258 607112 317494
rect 607348 317258 607432 317494
rect 607668 317258 607700 317494
rect -23776 317174 607700 317258
rect -23776 316938 -23744 317174
rect -23508 316938 -23424 317174
rect -23188 316938 607112 317174
rect 607348 316938 607432 317174
rect 607668 316938 607700 317174
rect -23776 316906 607700 316938
rect -23776 313774 607700 313806
rect -23776 313538 -20634 313774
rect -20398 313538 -20314 313774
rect -20078 313538 604002 313774
rect 604238 313538 604322 313774
rect 604558 313538 607700 313774
rect -23776 313454 607700 313538
rect -23776 313218 -20634 313454
rect -20398 313218 -20314 313454
rect -20078 313218 604002 313454
rect 604238 313218 604322 313454
rect 604558 313218 607700 313454
rect -23776 313186 607700 313218
rect -23776 310054 607700 310086
rect -23776 309818 -17524 310054
rect -17288 309818 -17204 310054
rect -16968 309818 600892 310054
rect 601128 309818 601212 310054
rect 601448 309818 607700 310054
rect -23776 309734 607700 309818
rect -23776 309498 -17524 309734
rect -17288 309498 -17204 309734
rect -16968 309498 600892 309734
rect 601128 309498 601212 309734
rect 601448 309498 607700 309734
rect -23776 309466 607700 309498
rect -23776 306334 607700 306366
rect -23776 306098 -14414 306334
rect -14178 306098 -14094 306334
rect -13858 306098 597782 306334
rect 598018 306098 598102 306334
rect 598338 306098 607700 306334
rect -23776 306014 607700 306098
rect -23776 305778 -14414 306014
rect -14178 305778 -14094 306014
rect -13858 305778 597782 306014
rect 598018 305778 598102 306014
rect 598338 305778 607700 306014
rect -23776 305746 607700 305778
rect -23776 302614 607700 302646
rect -23776 302378 -11304 302614
rect -11068 302378 -10984 302614
rect -10748 302378 594672 302614
rect 594908 302378 594992 302614
rect 595228 302378 607700 302614
rect -23776 302294 607700 302378
rect -23776 302058 -11304 302294
rect -11068 302058 -10984 302294
rect -10748 302058 594672 302294
rect 594908 302058 594992 302294
rect 595228 302058 607700 302294
rect -23776 302026 607700 302058
rect -23776 298894 607700 298926
rect -23776 298658 -8194 298894
rect -7958 298658 -7874 298894
rect -7638 298658 591562 298894
rect 591798 298658 591882 298894
rect 592118 298658 607700 298894
rect -23776 298574 607700 298658
rect -23776 298338 -8194 298574
rect -7958 298338 -7874 298574
rect -7638 298338 591562 298574
rect 591798 298338 591882 298574
rect 592118 298338 607700 298574
rect -23776 298306 607700 298338
rect -23776 295174 607700 295206
rect -23776 294938 -5084 295174
rect -4848 294938 -4764 295174
rect -4528 294938 7876 295174
rect 8112 294938 8196 295174
rect 8432 294938 38032 295174
rect 38268 294938 38352 295174
rect 38588 294938 74032 295174
rect 74268 294938 74352 295174
rect 74588 294938 110032 295174
rect 110268 294938 110352 295174
rect 110588 294938 146032 295174
rect 146268 294938 146352 295174
rect 146588 294938 182032 295174
rect 182268 294938 182352 295174
rect 182588 294938 218032 295174
rect 218268 294938 218352 295174
rect 218588 294938 254032 295174
rect 254268 294938 254352 295174
rect 254588 294938 290032 295174
rect 290268 294938 290352 295174
rect 290588 294938 326032 295174
rect 326268 294938 326352 295174
rect 326588 294938 362032 295174
rect 362268 294938 362352 295174
rect 362588 294938 398032 295174
rect 398268 294938 398352 295174
rect 398588 294938 434032 295174
rect 434268 294938 434352 295174
rect 434588 294938 470032 295174
rect 470268 294938 470352 295174
rect 470588 294938 506032 295174
rect 506268 294938 506352 295174
rect 506588 294938 542032 295174
rect 542268 294938 542352 295174
rect 542588 294938 571532 295174
rect 571768 294938 571852 295174
rect 572088 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 588452 295174
rect 588688 294938 588772 295174
rect 589008 294938 607700 295174
rect -23776 294854 607700 294938
rect -23776 294618 -5084 294854
rect -4848 294618 -4764 294854
rect -4528 294618 7876 294854
rect 8112 294618 8196 294854
rect 8432 294618 38032 294854
rect 38268 294618 38352 294854
rect 38588 294618 74032 294854
rect 74268 294618 74352 294854
rect 74588 294618 110032 294854
rect 110268 294618 110352 294854
rect 110588 294618 146032 294854
rect 146268 294618 146352 294854
rect 146588 294618 182032 294854
rect 182268 294618 182352 294854
rect 182588 294618 218032 294854
rect 218268 294618 218352 294854
rect 218588 294618 254032 294854
rect 254268 294618 254352 294854
rect 254588 294618 290032 294854
rect 290268 294618 290352 294854
rect 290588 294618 326032 294854
rect 326268 294618 326352 294854
rect 326588 294618 362032 294854
rect 362268 294618 362352 294854
rect 362588 294618 398032 294854
rect 398268 294618 398352 294854
rect 398588 294618 434032 294854
rect 434268 294618 434352 294854
rect 434588 294618 470032 294854
rect 470268 294618 470352 294854
rect 470588 294618 506032 294854
rect 506268 294618 506352 294854
rect 506588 294618 542032 294854
rect 542268 294618 542352 294854
rect 542588 294618 571532 294854
rect 571768 294618 571852 294854
rect 572088 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 588452 294854
rect 588688 294618 588772 294854
rect 589008 294618 607700 294854
rect -23776 294586 607700 294618
rect -23776 291454 607700 291486
rect -23776 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 9116 291454
rect 9352 291218 9436 291454
rect 9672 291218 56652 291454
rect 56888 291218 56972 291454
rect 57208 291218 92652 291454
rect 92888 291218 92972 291454
rect 93208 291218 128652 291454
rect 128888 291218 128972 291454
rect 129208 291218 164652 291454
rect 164888 291218 164972 291454
rect 165208 291218 200652 291454
rect 200888 291218 200972 291454
rect 201208 291218 236652 291454
rect 236888 291218 236972 291454
rect 237208 291218 272652 291454
rect 272888 291218 272972 291454
rect 273208 291218 308652 291454
rect 308888 291218 308972 291454
rect 309208 291218 344652 291454
rect 344888 291218 344972 291454
rect 345208 291218 380652 291454
rect 380888 291218 380972 291454
rect 381208 291218 416652 291454
rect 416888 291218 416972 291454
rect 417208 291218 452652 291454
rect 452888 291218 452972 291454
rect 453208 291218 488652 291454
rect 488888 291218 488972 291454
rect 489208 291218 524652 291454
rect 524888 291218 524972 291454
rect 525208 291218 560652 291454
rect 560888 291218 560972 291454
rect 561208 291218 570292 291454
rect 570528 291218 570612 291454
rect 570848 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 607700 291454
rect -23776 291134 607700 291218
rect -23776 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 9116 291134
rect 9352 290898 9436 291134
rect 9672 290898 56652 291134
rect 56888 290898 56972 291134
rect 57208 290898 92652 291134
rect 92888 290898 92972 291134
rect 93208 290898 128652 291134
rect 128888 290898 128972 291134
rect 129208 290898 164652 291134
rect 164888 290898 164972 291134
rect 165208 290898 200652 291134
rect 200888 290898 200972 291134
rect 201208 290898 236652 291134
rect 236888 290898 236972 291134
rect 237208 290898 272652 291134
rect 272888 290898 272972 291134
rect 273208 290898 308652 291134
rect 308888 290898 308972 291134
rect 309208 290898 344652 291134
rect 344888 290898 344972 291134
rect 345208 290898 380652 291134
rect 380888 290898 380972 291134
rect 381208 290898 416652 291134
rect 416888 290898 416972 291134
rect 417208 290898 452652 291134
rect 452888 290898 452972 291134
rect 453208 290898 488652 291134
rect 488888 290898 488972 291134
rect 489208 290898 524652 291134
rect 524888 290898 524972 291134
rect 525208 290898 560652 291134
rect 560888 290898 560972 291134
rect 561208 290898 570292 291134
rect 570528 290898 570612 291134
rect 570848 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 607700 291134
rect -23776 290866 607700 290898
rect -23776 281494 607700 281526
rect -23776 281258 -23744 281494
rect -23508 281258 -23424 281494
rect -23188 281258 607112 281494
rect 607348 281258 607432 281494
rect 607668 281258 607700 281494
rect -23776 281174 607700 281258
rect -23776 280938 -23744 281174
rect -23508 280938 -23424 281174
rect -23188 280938 607112 281174
rect 607348 280938 607432 281174
rect 607668 280938 607700 281174
rect -23776 280906 607700 280938
rect -23776 277774 607700 277806
rect -23776 277538 -20634 277774
rect -20398 277538 -20314 277774
rect -20078 277538 604002 277774
rect 604238 277538 604322 277774
rect 604558 277538 607700 277774
rect -23776 277454 607700 277538
rect -23776 277218 -20634 277454
rect -20398 277218 -20314 277454
rect -20078 277218 604002 277454
rect 604238 277218 604322 277454
rect 604558 277218 607700 277454
rect -23776 277186 607700 277218
rect -23776 274054 607700 274086
rect -23776 273818 -17524 274054
rect -17288 273818 -17204 274054
rect -16968 273818 600892 274054
rect 601128 273818 601212 274054
rect 601448 273818 607700 274054
rect -23776 273734 607700 273818
rect -23776 273498 -17524 273734
rect -17288 273498 -17204 273734
rect -16968 273498 600892 273734
rect 601128 273498 601212 273734
rect 601448 273498 607700 273734
rect -23776 273466 607700 273498
rect -23776 270334 607700 270366
rect -23776 270098 -14414 270334
rect -14178 270098 -14094 270334
rect -13858 270098 597782 270334
rect 598018 270098 598102 270334
rect 598338 270098 607700 270334
rect -23776 270014 607700 270098
rect -23776 269778 -14414 270014
rect -14178 269778 -14094 270014
rect -13858 269778 597782 270014
rect 598018 269778 598102 270014
rect 598338 269778 607700 270014
rect -23776 269746 607700 269778
rect -23776 266614 607700 266646
rect -23776 266378 -11304 266614
rect -11068 266378 -10984 266614
rect -10748 266378 594672 266614
rect 594908 266378 594992 266614
rect 595228 266378 607700 266614
rect -23776 266294 607700 266378
rect -23776 266058 -11304 266294
rect -11068 266058 -10984 266294
rect -10748 266058 594672 266294
rect 594908 266058 594992 266294
rect 595228 266058 607700 266294
rect -23776 266026 607700 266058
rect -23776 262894 607700 262926
rect -23776 262658 -8194 262894
rect -7958 262658 -7874 262894
rect -7638 262658 591562 262894
rect 591798 262658 591882 262894
rect 592118 262658 607700 262894
rect -23776 262574 607700 262658
rect -23776 262338 -8194 262574
rect -7958 262338 -7874 262574
rect -7638 262338 591562 262574
rect 591798 262338 591882 262574
rect 592118 262338 607700 262574
rect -23776 262306 607700 262338
rect -23776 259174 607700 259206
rect -23776 258938 -5084 259174
rect -4848 258938 -4764 259174
rect -4528 258938 7876 259174
rect 8112 258938 8196 259174
rect 8432 258938 38032 259174
rect 38268 258938 38352 259174
rect 38588 258938 74032 259174
rect 74268 258938 74352 259174
rect 74588 258938 110032 259174
rect 110268 258938 110352 259174
rect 110588 258938 146032 259174
rect 146268 258938 146352 259174
rect 146588 258938 182032 259174
rect 182268 258938 182352 259174
rect 182588 258938 218032 259174
rect 218268 258938 218352 259174
rect 218588 258938 254032 259174
rect 254268 258938 254352 259174
rect 254588 258938 290032 259174
rect 290268 258938 290352 259174
rect 290588 258938 326032 259174
rect 326268 258938 326352 259174
rect 326588 258938 362032 259174
rect 362268 258938 362352 259174
rect 362588 258938 398032 259174
rect 398268 258938 398352 259174
rect 398588 258938 434032 259174
rect 434268 258938 434352 259174
rect 434588 258938 470032 259174
rect 470268 258938 470352 259174
rect 470588 258938 506032 259174
rect 506268 258938 506352 259174
rect 506588 258938 542032 259174
rect 542268 258938 542352 259174
rect 542588 258938 571532 259174
rect 571768 258938 571852 259174
rect 572088 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 588452 259174
rect 588688 258938 588772 259174
rect 589008 258938 607700 259174
rect -23776 258854 607700 258938
rect -23776 258618 -5084 258854
rect -4848 258618 -4764 258854
rect -4528 258618 7876 258854
rect 8112 258618 8196 258854
rect 8432 258618 38032 258854
rect 38268 258618 38352 258854
rect 38588 258618 74032 258854
rect 74268 258618 74352 258854
rect 74588 258618 110032 258854
rect 110268 258618 110352 258854
rect 110588 258618 146032 258854
rect 146268 258618 146352 258854
rect 146588 258618 182032 258854
rect 182268 258618 182352 258854
rect 182588 258618 218032 258854
rect 218268 258618 218352 258854
rect 218588 258618 254032 258854
rect 254268 258618 254352 258854
rect 254588 258618 290032 258854
rect 290268 258618 290352 258854
rect 290588 258618 326032 258854
rect 326268 258618 326352 258854
rect 326588 258618 362032 258854
rect 362268 258618 362352 258854
rect 362588 258618 398032 258854
rect 398268 258618 398352 258854
rect 398588 258618 434032 258854
rect 434268 258618 434352 258854
rect 434588 258618 470032 258854
rect 470268 258618 470352 258854
rect 470588 258618 506032 258854
rect 506268 258618 506352 258854
rect 506588 258618 542032 258854
rect 542268 258618 542352 258854
rect 542588 258618 571532 258854
rect 571768 258618 571852 258854
rect 572088 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 588452 258854
rect 588688 258618 588772 258854
rect 589008 258618 607700 258854
rect -23776 258586 607700 258618
rect -23776 255454 607700 255486
rect -23776 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 9116 255454
rect 9352 255218 9436 255454
rect 9672 255218 56652 255454
rect 56888 255218 56972 255454
rect 57208 255218 92652 255454
rect 92888 255218 92972 255454
rect 93208 255218 128652 255454
rect 128888 255218 128972 255454
rect 129208 255218 164652 255454
rect 164888 255218 164972 255454
rect 165208 255218 200652 255454
rect 200888 255218 200972 255454
rect 201208 255218 236652 255454
rect 236888 255218 236972 255454
rect 237208 255218 272652 255454
rect 272888 255218 272972 255454
rect 273208 255218 308652 255454
rect 308888 255218 308972 255454
rect 309208 255218 344652 255454
rect 344888 255218 344972 255454
rect 345208 255218 380652 255454
rect 380888 255218 380972 255454
rect 381208 255218 416652 255454
rect 416888 255218 416972 255454
rect 417208 255218 452652 255454
rect 452888 255218 452972 255454
rect 453208 255218 488652 255454
rect 488888 255218 488972 255454
rect 489208 255218 524652 255454
rect 524888 255218 524972 255454
rect 525208 255218 560652 255454
rect 560888 255218 560972 255454
rect 561208 255218 570292 255454
rect 570528 255218 570612 255454
rect 570848 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 607700 255454
rect -23776 255134 607700 255218
rect -23776 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 9116 255134
rect 9352 254898 9436 255134
rect 9672 254898 56652 255134
rect 56888 254898 56972 255134
rect 57208 254898 92652 255134
rect 92888 254898 92972 255134
rect 93208 254898 128652 255134
rect 128888 254898 128972 255134
rect 129208 254898 164652 255134
rect 164888 254898 164972 255134
rect 165208 254898 200652 255134
rect 200888 254898 200972 255134
rect 201208 254898 236652 255134
rect 236888 254898 236972 255134
rect 237208 254898 272652 255134
rect 272888 254898 272972 255134
rect 273208 254898 308652 255134
rect 308888 254898 308972 255134
rect 309208 254898 344652 255134
rect 344888 254898 344972 255134
rect 345208 254898 380652 255134
rect 380888 254898 380972 255134
rect 381208 254898 416652 255134
rect 416888 254898 416972 255134
rect 417208 254898 452652 255134
rect 452888 254898 452972 255134
rect 453208 254898 488652 255134
rect 488888 254898 488972 255134
rect 489208 254898 524652 255134
rect 524888 254898 524972 255134
rect 525208 254898 560652 255134
rect 560888 254898 560972 255134
rect 561208 254898 570292 255134
rect 570528 254898 570612 255134
rect 570848 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 607700 255134
rect -23776 254866 607700 254898
rect -23776 245494 607700 245526
rect -23776 245258 -23744 245494
rect -23508 245258 -23424 245494
rect -23188 245258 607112 245494
rect 607348 245258 607432 245494
rect 607668 245258 607700 245494
rect -23776 245174 607700 245258
rect -23776 244938 -23744 245174
rect -23508 244938 -23424 245174
rect -23188 244938 607112 245174
rect 607348 244938 607432 245174
rect 607668 244938 607700 245174
rect -23776 244906 607700 244938
rect -23776 241774 607700 241806
rect -23776 241538 -20634 241774
rect -20398 241538 -20314 241774
rect -20078 241538 604002 241774
rect 604238 241538 604322 241774
rect 604558 241538 607700 241774
rect -23776 241454 607700 241538
rect -23776 241218 -20634 241454
rect -20398 241218 -20314 241454
rect -20078 241218 604002 241454
rect 604238 241218 604322 241454
rect 604558 241218 607700 241454
rect -23776 241186 607700 241218
rect -23776 238054 607700 238086
rect -23776 237818 -17524 238054
rect -17288 237818 -17204 238054
rect -16968 237818 600892 238054
rect 601128 237818 601212 238054
rect 601448 237818 607700 238054
rect -23776 237734 607700 237818
rect -23776 237498 -17524 237734
rect -17288 237498 -17204 237734
rect -16968 237498 600892 237734
rect 601128 237498 601212 237734
rect 601448 237498 607700 237734
rect -23776 237466 607700 237498
rect -23776 234334 607700 234366
rect -23776 234098 -14414 234334
rect -14178 234098 -14094 234334
rect -13858 234098 597782 234334
rect 598018 234098 598102 234334
rect 598338 234098 607700 234334
rect -23776 234014 607700 234098
rect -23776 233778 -14414 234014
rect -14178 233778 -14094 234014
rect -13858 233778 597782 234014
rect 598018 233778 598102 234014
rect 598338 233778 607700 234014
rect -23776 233746 607700 233778
rect -23776 230614 607700 230646
rect -23776 230378 -11304 230614
rect -11068 230378 -10984 230614
rect -10748 230378 594672 230614
rect 594908 230378 594992 230614
rect 595228 230378 607700 230614
rect -23776 230294 607700 230378
rect -23776 230058 -11304 230294
rect -11068 230058 -10984 230294
rect -10748 230058 594672 230294
rect 594908 230058 594992 230294
rect 595228 230058 607700 230294
rect -23776 230026 607700 230058
rect -23776 226894 607700 226926
rect -23776 226658 -8194 226894
rect -7958 226658 -7874 226894
rect -7638 226658 591562 226894
rect 591798 226658 591882 226894
rect 592118 226658 607700 226894
rect -23776 226574 607700 226658
rect -23776 226338 -8194 226574
rect -7958 226338 -7874 226574
rect -7638 226338 591562 226574
rect 591798 226338 591882 226574
rect 592118 226338 607700 226574
rect -23776 226306 607700 226338
rect -23776 223174 607700 223206
rect -23776 222938 -5084 223174
rect -4848 222938 -4764 223174
rect -4528 222938 7876 223174
rect 8112 222938 8196 223174
rect 8432 222938 38032 223174
rect 38268 222938 38352 223174
rect 38588 222938 74032 223174
rect 74268 222938 74352 223174
rect 74588 222938 110032 223174
rect 110268 222938 110352 223174
rect 110588 222938 146032 223174
rect 146268 222938 146352 223174
rect 146588 222938 182032 223174
rect 182268 222938 182352 223174
rect 182588 222938 218032 223174
rect 218268 222938 218352 223174
rect 218588 222938 254032 223174
rect 254268 222938 254352 223174
rect 254588 222938 290032 223174
rect 290268 222938 290352 223174
rect 290588 222938 326032 223174
rect 326268 222938 326352 223174
rect 326588 222938 362032 223174
rect 362268 222938 362352 223174
rect 362588 222938 398032 223174
rect 398268 222938 398352 223174
rect 398588 222938 434032 223174
rect 434268 222938 434352 223174
rect 434588 222938 470032 223174
rect 470268 222938 470352 223174
rect 470588 222938 506032 223174
rect 506268 222938 506352 223174
rect 506588 222938 542032 223174
rect 542268 222938 542352 223174
rect 542588 222938 571532 223174
rect 571768 222938 571852 223174
rect 572088 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 588452 223174
rect 588688 222938 588772 223174
rect 589008 222938 607700 223174
rect -23776 222854 607700 222938
rect -23776 222618 -5084 222854
rect -4848 222618 -4764 222854
rect -4528 222618 7876 222854
rect 8112 222618 8196 222854
rect 8432 222618 38032 222854
rect 38268 222618 38352 222854
rect 38588 222618 74032 222854
rect 74268 222618 74352 222854
rect 74588 222618 110032 222854
rect 110268 222618 110352 222854
rect 110588 222618 146032 222854
rect 146268 222618 146352 222854
rect 146588 222618 182032 222854
rect 182268 222618 182352 222854
rect 182588 222618 218032 222854
rect 218268 222618 218352 222854
rect 218588 222618 254032 222854
rect 254268 222618 254352 222854
rect 254588 222618 290032 222854
rect 290268 222618 290352 222854
rect 290588 222618 326032 222854
rect 326268 222618 326352 222854
rect 326588 222618 362032 222854
rect 362268 222618 362352 222854
rect 362588 222618 398032 222854
rect 398268 222618 398352 222854
rect 398588 222618 434032 222854
rect 434268 222618 434352 222854
rect 434588 222618 470032 222854
rect 470268 222618 470352 222854
rect 470588 222618 506032 222854
rect 506268 222618 506352 222854
rect 506588 222618 542032 222854
rect 542268 222618 542352 222854
rect 542588 222618 571532 222854
rect 571768 222618 571852 222854
rect 572088 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 588452 222854
rect 588688 222618 588772 222854
rect 589008 222618 607700 222854
rect -23776 222586 607700 222618
rect -23776 219454 607700 219486
rect -23776 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 9116 219454
rect 9352 219218 9436 219454
rect 9672 219218 56652 219454
rect 56888 219218 56972 219454
rect 57208 219218 92652 219454
rect 92888 219218 92972 219454
rect 93208 219218 128652 219454
rect 128888 219218 128972 219454
rect 129208 219218 164652 219454
rect 164888 219218 164972 219454
rect 165208 219218 200652 219454
rect 200888 219218 200972 219454
rect 201208 219218 236652 219454
rect 236888 219218 236972 219454
rect 237208 219218 272652 219454
rect 272888 219218 272972 219454
rect 273208 219218 308652 219454
rect 308888 219218 308972 219454
rect 309208 219218 344652 219454
rect 344888 219218 344972 219454
rect 345208 219218 380652 219454
rect 380888 219218 380972 219454
rect 381208 219218 416652 219454
rect 416888 219218 416972 219454
rect 417208 219218 452652 219454
rect 452888 219218 452972 219454
rect 453208 219218 488652 219454
rect 488888 219218 488972 219454
rect 489208 219218 524652 219454
rect 524888 219218 524972 219454
rect 525208 219218 560652 219454
rect 560888 219218 560972 219454
rect 561208 219218 570292 219454
rect 570528 219218 570612 219454
rect 570848 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 607700 219454
rect -23776 219134 607700 219218
rect -23776 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 9116 219134
rect 9352 218898 9436 219134
rect 9672 218898 56652 219134
rect 56888 218898 56972 219134
rect 57208 218898 92652 219134
rect 92888 218898 92972 219134
rect 93208 218898 128652 219134
rect 128888 218898 128972 219134
rect 129208 218898 164652 219134
rect 164888 218898 164972 219134
rect 165208 218898 200652 219134
rect 200888 218898 200972 219134
rect 201208 218898 236652 219134
rect 236888 218898 236972 219134
rect 237208 218898 272652 219134
rect 272888 218898 272972 219134
rect 273208 218898 308652 219134
rect 308888 218898 308972 219134
rect 309208 218898 344652 219134
rect 344888 218898 344972 219134
rect 345208 218898 380652 219134
rect 380888 218898 380972 219134
rect 381208 218898 416652 219134
rect 416888 218898 416972 219134
rect 417208 218898 452652 219134
rect 452888 218898 452972 219134
rect 453208 218898 488652 219134
rect 488888 218898 488972 219134
rect 489208 218898 524652 219134
rect 524888 218898 524972 219134
rect 525208 218898 560652 219134
rect 560888 218898 560972 219134
rect 561208 218898 570292 219134
rect 570528 218898 570612 219134
rect 570848 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 607700 219134
rect -23776 218866 607700 218898
rect -23776 209494 607700 209526
rect -23776 209258 -23744 209494
rect -23508 209258 -23424 209494
rect -23188 209258 607112 209494
rect 607348 209258 607432 209494
rect 607668 209258 607700 209494
rect -23776 209174 607700 209258
rect -23776 208938 -23744 209174
rect -23508 208938 -23424 209174
rect -23188 208938 607112 209174
rect 607348 208938 607432 209174
rect 607668 208938 607700 209174
rect -23776 208906 607700 208938
rect -23776 205774 607700 205806
rect -23776 205538 -20634 205774
rect -20398 205538 -20314 205774
rect -20078 205538 604002 205774
rect 604238 205538 604322 205774
rect 604558 205538 607700 205774
rect -23776 205454 607700 205538
rect -23776 205218 -20634 205454
rect -20398 205218 -20314 205454
rect -20078 205218 604002 205454
rect 604238 205218 604322 205454
rect 604558 205218 607700 205454
rect -23776 205186 607700 205218
rect -23776 202054 607700 202086
rect -23776 201818 -17524 202054
rect -17288 201818 -17204 202054
rect -16968 201818 600892 202054
rect 601128 201818 601212 202054
rect 601448 201818 607700 202054
rect -23776 201734 607700 201818
rect -23776 201498 -17524 201734
rect -17288 201498 -17204 201734
rect -16968 201498 600892 201734
rect 601128 201498 601212 201734
rect 601448 201498 607700 201734
rect -23776 201466 607700 201498
rect -23776 198334 607700 198366
rect -23776 198098 -14414 198334
rect -14178 198098 -14094 198334
rect -13858 198098 597782 198334
rect 598018 198098 598102 198334
rect 598338 198098 607700 198334
rect -23776 198014 607700 198098
rect -23776 197778 -14414 198014
rect -14178 197778 -14094 198014
rect -13858 197778 597782 198014
rect 598018 197778 598102 198014
rect 598338 197778 607700 198014
rect -23776 197746 607700 197778
rect -23776 194614 607700 194646
rect -23776 194378 -11304 194614
rect -11068 194378 -10984 194614
rect -10748 194378 594672 194614
rect 594908 194378 594992 194614
rect 595228 194378 607700 194614
rect -23776 194294 607700 194378
rect -23776 194058 -11304 194294
rect -11068 194058 -10984 194294
rect -10748 194058 594672 194294
rect 594908 194058 594992 194294
rect 595228 194058 607700 194294
rect -23776 194026 607700 194058
rect -23776 190894 607700 190926
rect -23776 190658 -8194 190894
rect -7958 190658 -7874 190894
rect -7638 190658 591562 190894
rect 591798 190658 591882 190894
rect 592118 190658 607700 190894
rect -23776 190574 607700 190658
rect -23776 190338 -8194 190574
rect -7958 190338 -7874 190574
rect -7638 190338 591562 190574
rect 591798 190338 591882 190574
rect 592118 190338 607700 190574
rect -23776 190306 607700 190338
rect -23776 187174 607700 187206
rect -23776 186938 -5084 187174
rect -4848 186938 -4764 187174
rect -4528 186938 7876 187174
rect 8112 186938 8196 187174
rect 8432 186938 38032 187174
rect 38268 186938 38352 187174
rect 38588 186938 60622 187174
rect 60858 186938 159098 187174
rect 159334 186938 182032 187174
rect 182268 186938 182352 187174
rect 182588 186938 185622 187174
rect 185858 186938 284098 187174
rect 284334 186938 290032 187174
rect 290268 186938 290352 187174
rect 290588 186938 310622 187174
rect 310858 186938 409098 187174
rect 409334 186938 434032 187174
rect 434268 186938 434352 187174
rect 434588 186938 436622 187174
rect 436858 186938 535098 187174
rect 535334 186938 542032 187174
rect 542268 186938 542352 187174
rect 542588 186938 571532 187174
rect 571768 186938 571852 187174
rect 572088 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 588452 187174
rect 588688 186938 588772 187174
rect 589008 186938 607700 187174
rect -23776 186854 607700 186938
rect -23776 186618 -5084 186854
rect -4848 186618 -4764 186854
rect -4528 186618 7876 186854
rect 8112 186618 8196 186854
rect 8432 186618 38032 186854
rect 38268 186618 38352 186854
rect 38588 186618 60622 186854
rect 60858 186618 159098 186854
rect 159334 186618 182032 186854
rect 182268 186618 182352 186854
rect 182588 186618 185622 186854
rect 185858 186618 284098 186854
rect 284334 186618 290032 186854
rect 290268 186618 290352 186854
rect 290588 186618 310622 186854
rect 310858 186618 409098 186854
rect 409334 186618 434032 186854
rect 434268 186618 434352 186854
rect 434588 186618 436622 186854
rect 436858 186618 535098 186854
rect 535334 186618 542032 186854
rect 542268 186618 542352 186854
rect 542588 186618 571532 186854
rect 571768 186618 571852 186854
rect 572088 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 588452 186854
rect 588688 186618 588772 186854
rect 589008 186618 607700 186854
rect -23776 186586 607700 186618
rect -23776 183454 607700 183486
rect -23776 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 9116 183454
rect 9352 183218 9436 183454
rect 9672 183218 56652 183454
rect 56888 183218 56972 183454
rect 57208 183218 61342 183454
rect 61578 183218 158378 183454
rect 158614 183218 164652 183454
rect 164888 183218 164972 183454
rect 165208 183218 186342 183454
rect 186578 183218 283378 183454
rect 283614 183218 308652 183454
rect 308888 183218 308972 183454
rect 309208 183218 311342 183454
rect 311578 183218 408378 183454
rect 408614 183218 416652 183454
rect 416888 183218 416972 183454
rect 417208 183218 437342 183454
rect 437578 183218 534378 183454
rect 534614 183218 560652 183454
rect 560888 183218 560972 183454
rect 561208 183218 570292 183454
rect 570528 183218 570612 183454
rect 570848 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 607700 183454
rect -23776 183134 607700 183218
rect -23776 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 9116 183134
rect 9352 182898 9436 183134
rect 9672 182898 56652 183134
rect 56888 182898 56972 183134
rect 57208 182898 61342 183134
rect 61578 182898 158378 183134
rect 158614 182898 164652 183134
rect 164888 182898 164972 183134
rect 165208 182898 186342 183134
rect 186578 182898 283378 183134
rect 283614 182898 308652 183134
rect 308888 182898 308972 183134
rect 309208 182898 311342 183134
rect 311578 182898 408378 183134
rect 408614 182898 416652 183134
rect 416888 182898 416972 183134
rect 417208 182898 437342 183134
rect 437578 182898 534378 183134
rect 534614 182898 560652 183134
rect 560888 182898 560972 183134
rect 561208 182898 570292 183134
rect 570528 182898 570612 183134
rect 570848 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 607700 183134
rect -23776 182866 607700 182898
rect -23776 173494 607700 173526
rect -23776 173258 -23744 173494
rect -23508 173258 -23424 173494
rect -23188 173258 607112 173494
rect 607348 173258 607432 173494
rect 607668 173258 607700 173494
rect -23776 173174 607700 173258
rect -23776 172938 -23744 173174
rect -23508 172938 -23424 173174
rect -23188 172938 607112 173174
rect 607348 172938 607432 173174
rect 607668 172938 607700 173174
rect -23776 172906 607700 172938
rect -23776 169774 607700 169806
rect -23776 169538 -20634 169774
rect -20398 169538 -20314 169774
rect -20078 169538 604002 169774
rect 604238 169538 604322 169774
rect 604558 169538 607700 169774
rect -23776 169454 607700 169538
rect -23776 169218 -20634 169454
rect -20398 169218 -20314 169454
rect -20078 169218 604002 169454
rect 604238 169218 604322 169454
rect 604558 169218 607700 169454
rect -23776 169186 607700 169218
rect -23776 166054 607700 166086
rect -23776 165818 -17524 166054
rect -17288 165818 -17204 166054
rect -16968 165818 600892 166054
rect 601128 165818 601212 166054
rect 601448 165818 607700 166054
rect -23776 165734 607700 165818
rect -23776 165498 -17524 165734
rect -17288 165498 -17204 165734
rect -16968 165498 600892 165734
rect 601128 165498 601212 165734
rect 601448 165498 607700 165734
rect -23776 165466 607700 165498
rect -23776 162334 607700 162366
rect -23776 162098 -14414 162334
rect -14178 162098 -14094 162334
rect -13858 162098 597782 162334
rect 598018 162098 598102 162334
rect 598338 162098 607700 162334
rect -23776 162014 607700 162098
rect -23776 161778 -14414 162014
rect -14178 161778 -14094 162014
rect -13858 161778 597782 162014
rect 598018 161778 598102 162014
rect 598338 161778 607700 162014
rect -23776 161746 607700 161778
rect -23776 158614 607700 158646
rect -23776 158378 -11304 158614
rect -11068 158378 -10984 158614
rect -10748 158378 594672 158614
rect 594908 158378 594992 158614
rect 595228 158378 607700 158614
rect -23776 158294 607700 158378
rect -23776 158058 -11304 158294
rect -11068 158058 -10984 158294
rect -10748 158058 594672 158294
rect 594908 158058 594992 158294
rect 595228 158058 607700 158294
rect -23776 158026 607700 158058
rect -23776 154894 607700 154926
rect -23776 154658 -8194 154894
rect -7958 154658 -7874 154894
rect -7638 154658 591562 154894
rect 591798 154658 591882 154894
rect 592118 154658 607700 154894
rect -23776 154574 607700 154658
rect -23776 154338 -8194 154574
rect -7958 154338 -7874 154574
rect -7638 154338 591562 154574
rect 591798 154338 591882 154574
rect 592118 154338 607700 154574
rect -23776 154306 607700 154338
rect -23776 151174 607700 151206
rect -23776 150938 -5084 151174
rect -4848 150938 -4764 151174
rect -4528 150938 7876 151174
rect 8112 150938 8196 151174
rect 8432 150938 38032 151174
rect 38268 150938 38352 151174
rect 38588 150938 60622 151174
rect 60858 150938 159098 151174
rect 159334 150938 182032 151174
rect 182268 150938 182352 151174
rect 182588 150938 185622 151174
rect 185858 150938 284098 151174
rect 284334 150938 290032 151174
rect 290268 150938 290352 151174
rect 290588 150938 310622 151174
rect 310858 150938 409098 151174
rect 409334 150938 434032 151174
rect 434268 150938 434352 151174
rect 434588 150938 436622 151174
rect 436858 150938 535098 151174
rect 535334 150938 542032 151174
rect 542268 150938 542352 151174
rect 542588 150938 571532 151174
rect 571768 150938 571852 151174
rect 572088 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 588452 151174
rect 588688 150938 588772 151174
rect 589008 150938 607700 151174
rect -23776 150854 607700 150938
rect -23776 150618 -5084 150854
rect -4848 150618 -4764 150854
rect -4528 150618 7876 150854
rect 8112 150618 8196 150854
rect 8432 150618 38032 150854
rect 38268 150618 38352 150854
rect 38588 150618 60622 150854
rect 60858 150618 159098 150854
rect 159334 150618 182032 150854
rect 182268 150618 182352 150854
rect 182588 150618 185622 150854
rect 185858 150618 284098 150854
rect 284334 150618 290032 150854
rect 290268 150618 290352 150854
rect 290588 150618 310622 150854
rect 310858 150618 409098 150854
rect 409334 150618 434032 150854
rect 434268 150618 434352 150854
rect 434588 150618 436622 150854
rect 436858 150618 535098 150854
rect 535334 150618 542032 150854
rect 542268 150618 542352 150854
rect 542588 150618 571532 150854
rect 571768 150618 571852 150854
rect 572088 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 588452 150854
rect 588688 150618 588772 150854
rect 589008 150618 607700 150854
rect -23776 150586 607700 150618
rect -23776 147454 607700 147486
rect -23776 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 9116 147454
rect 9352 147218 9436 147454
rect 9672 147218 56652 147454
rect 56888 147218 56972 147454
rect 57208 147218 61342 147454
rect 61578 147218 158378 147454
rect 158614 147218 164652 147454
rect 164888 147218 164972 147454
rect 165208 147218 186342 147454
rect 186578 147218 283378 147454
rect 283614 147218 308652 147454
rect 308888 147218 308972 147454
rect 309208 147218 311342 147454
rect 311578 147218 408378 147454
rect 408614 147218 416652 147454
rect 416888 147218 416972 147454
rect 417208 147218 437342 147454
rect 437578 147218 534378 147454
rect 534614 147218 560652 147454
rect 560888 147218 560972 147454
rect 561208 147218 570292 147454
rect 570528 147218 570612 147454
rect 570848 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 607700 147454
rect -23776 147134 607700 147218
rect -23776 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 9116 147134
rect 9352 146898 9436 147134
rect 9672 146898 56652 147134
rect 56888 146898 56972 147134
rect 57208 146898 61342 147134
rect 61578 146898 158378 147134
rect 158614 146898 164652 147134
rect 164888 146898 164972 147134
rect 165208 146898 186342 147134
rect 186578 146898 283378 147134
rect 283614 146898 308652 147134
rect 308888 146898 308972 147134
rect 309208 146898 311342 147134
rect 311578 146898 408378 147134
rect 408614 146898 416652 147134
rect 416888 146898 416972 147134
rect 417208 146898 437342 147134
rect 437578 146898 534378 147134
rect 534614 146898 560652 147134
rect 560888 146898 560972 147134
rect 561208 146898 570292 147134
rect 570528 146898 570612 147134
rect 570848 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 607700 147134
rect -23776 146866 607700 146898
rect -23776 137494 607700 137526
rect -23776 137258 -23744 137494
rect -23508 137258 -23424 137494
rect -23188 137258 607112 137494
rect 607348 137258 607432 137494
rect 607668 137258 607700 137494
rect -23776 137174 607700 137258
rect -23776 136938 -23744 137174
rect -23508 136938 -23424 137174
rect -23188 136938 607112 137174
rect 607348 136938 607432 137174
rect 607668 136938 607700 137174
rect -23776 136906 607700 136938
rect -23776 133774 607700 133806
rect -23776 133538 -20634 133774
rect -20398 133538 -20314 133774
rect -20078 133538 604002 133774
rect 604238 133538 604322 133774
rect 604558 133538 607700 133774
rect -23776 133454 607700 133538
rect -23776 133218 -20634 133454
rect -20398 133218 -20314 133454
rect -20078 133218 604002 133454
rect 604238 133218 604322 133454
rect 604558 133218 607700 133454
rect -23776 133186 607700 133218
rect -23776 130054 607700 130086
rect -23776 129818 -17524 130054
rect -17288 129818 -17204 130054
rect -16968 129818 600892 130054
rect 601128 129818 601212 130054
rect 601448 129818 607700 130054
rect -23776 129734 607700 129818
rect -23776 129498 -17524 129734
rect -17288 129498 -17204 129734
rect -16968 129498 600892 129734
rect 601128 129498 601212 129734
rect 601448 129498 607700 129734
rect -23776 129466 607700 129498
rect -23776 126334 607700 126366
rect -23776 126098 -14414 126334
rect -14178 126098 -14094 126334
rect -13858 126098 597782 126334
rect 598018 126098 598102 126334
rect 598338 126098 607700 126334
rect -23776 126014 607700 126098
rect -23776 125778 -14414 126014
rect -14178 125778 -14094 126014
rect -13858 125778 597782 126014
rect 598018 125778 598102 126014
rect 598338 125778 607700 126014
rect -23776 125746 607700 125778
rect -23776 122614 607700 122646
rect -23776 122378 -11304 122614
rect -11068 122378 -10984 122614
rect -10748 122378 594672 122614
rect 594908 122378 594992 122614
rect 595228 122378 607700 122614
rect -23776 122294 607700 122378
rect -23776 122058 -11304 122294
rect -11068 122058 -10984 122294
rect -10748 122058 594672 122294
rect 594908 122058 594992 122294
rect 595228 122058 607700 122294
rect -23776 122026 607700 122058
rect 61280 121244 61640 121300
rect 61280 121008 61342 121244
rect 61578 121008 61640 121244
rect 61280 120952 61640 121008
rect 62952 121244 63300 121300
rect 62952 121008 63008 121244
rect 63244 121008 63300 121244
rect 62952 120952 63300 121008
rect 281656 121244 282004 121300
rect 281656 121008 281712 121244
rect 281948 121008 282004 121244
rect 281656 120952 282004 121008
rect 283316 121244 283676 121300
rect 283316 121008 283378 121244
rect 283614 121008 283676 121244
rect 283316 120952 283676 121008
rect 311280 121244 311640 121300
rect 311280 121008 311342 121244
rect 311578 121008 311640 121244
rect 311280 120952 311640 121008
rect 312952 121244 313300 121300
rect 312952 121008 313008 121244
rect 313244 121008 313300 121244
rect 312952 120952 313300 121008
rect 532656 121244 533004 121300
rect 532656 121008 532712 121244
rect 532948 121008 533004 121244
rect 532656 120952 533004 121008
rect 534316 121244 534676 121300
rect 534316 121008 534378 121244
rect 534614 121008 534676 121244
rect 534316 120952 534676 121008
rect 157336 120564 157684 120620
rect 157336 120328 157392 120564
rect 157628 120328 157684 120564
rect 157336 120272 157684 120328
rect 159036 120564 159396 120620
rect 159036 120328 159098 120564
rect 159334 120328 159396 120564
rect 159036 120272 159396 120328
rect 185560 120564 185920 120620
rect 185560 120328 185622 120564
rect 185858 120328 185920 120564
rect 185560 120272 185920 120328
rect 187272 120564 187620 120620
rect 187272 120328 187328 120564
rect 187564 120328 187620 120564
rect 187272 120272 187620 120328
rect 407336 120564 407684 120620
rect 407336 120328 407392 120564
rect 407628 120328 407684 120564
rect 407336 120272 407684 120328
rect 409036 120564 409396 120620
rect 409036 120328 409098 120564
rect 409334 120328 409396 120564
rect 409036 120272 409396 120328
rect 436560 120564 436920 120620
rect 436560 120328 436622 120564
rect 436858 120328 436920 120564
rect 436560 120272 436920 120328
rect 438272 120564 438620 120620
rect 438272 120328 438328 120564
rect 438564 120328 438620 120564
rect 438272 120272 438620 120328
rect -23776 118894 607700 118926
rect -23776 118658 -8194 118894
rect -7958 118658 -7874 118894
rect -7638 118658 591562 118894
rect 591798 118658 591882 118894
rect 592118 118658 607700 118894
rect -23776 118574 607700 118658
rect -23776 118338 -8194 118574
rect -7958 118338 -7874 118574
rect -7638 118338 591562 118574
rect 591798 118338 591882 118574
rect 592118 118338 607700 118574
rect -23776 118306 607700 118338
rect -23776 115174 607700 115206
rect -23776 114938 -5084 115174
rect -4848 114938 -4764 115174
rect -4528 114938 7876 115174
rect 8112 114938 8196 115174
rect 8432 114938 38032 115174
rect 38268 114938 38352 115174
rect 38588 114938 74032 115174
rect 74268 114938 74352 115174
rect 74588 114938 110032 115174
rect 110268 114938 110352 115174
rect 110588 114938 146032 115174
rect 146268 114938 146352 115174
rect 146588 114938 182032 115174
rect 182268 114938 182352 115174
rect 182588 114938 218032 115174
rect 218268 114938 218352 115174
rect 218588 114938 254032 115174
rect 254268 114938 254352 115174
rect 254588 114938 290032 115174
rect 290268 114938 290352 115174
rect 290588 114938 326032 115174
rect 326268 114938 326352 115174
rect 326588 114938 362032 115174
rect 362268 114938 362352 115174
rect 362588 114938 398032 115174
rect 398268 114938 398352 115174
rect 398588 114938 434032 115174
rect 434268 114938 434352 115174
rect 434588 114938 470032 115174
rect 470268 114938 470352 115174
rect 470588 114938 506032 115174
rect 506268 114938 506352 115174
rect 506588 114938 542032 115174
rect 542268 114938 542352 115174
rect 542588 114938 571532 115174
rect 571768 114938 571852 115174
rect 572088 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 588452 115174
rect 588688 114938 588772 115174
rect 589008 114938 607700 115174
rect -23776 114854 607700 114938
rect -23776 114618 -5084 114854
rect -4848 114618 -4764 114854
rect -4528 114618 7876 114854
rect 8112 114618 8196 114854
rect 8432 114618 38032 114854
rect 38268 114618 38352 114854
rect 38588 114618 74032 114854
rect 74268 114618 74352 114854
rect 74588 114618 110032 114854
rect 110268 114618 110352 114854
rect 110588 114618 146032 114854
rect 146268 114618 146352 114854
rect 146588 114618 182032 114854
rect 182268 114618 182352 114854
rect 182588 114618 218032 114854
rect 218268 114618 218352 114854
rect 218588 114618 254032 114854
rect 254268 114618 254352 114854
rect 254588 114618 290032 114854
rect 290268 114618 290352 114854
rect 290588 114618 326032 114854
rect 326268 114618 326352 114854
rect 326588 114618 362032 114854
rect 362268 114618 362352 114854
rect 362588 114618 398032 114854
rect 398268 114618 398352 114854
rect 398588 114618 434032 114854
rect 434268 114618 434352 114854
rect 434588 114618 470032 114854
rect 470268 114618 470352 114854
rect 470588 114618 506032 114854
rect 506268 114618 506352 114854
rect 506588 114618 542032 114854
rect 542268 114618 542352 114854
rect 542588 114618 571532 114854
rect 571768 114618 571852 114854
rect 572088 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 588452 114854
rect 588688 114618 588772 114854
rect 589008 114618 607700 114854
rect -23776 114586 607700 114618
rect -23776 111454 607700 111486
rect -23776 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 9116 111454
rect 9352 111218 9436 111454
rect 9672 111218 56652 111454
rect 56888 111218 56972 111454
rect 57208 111218 92652 111454
rect 92888 111218 92972 111454
rect 93208 111218 128652 111454
rect 128888 111218 128972 111454
rect 129208 111218 164652 111454
rect 164888 111218 164972 111454
rect 165208 111218 200652 111454
rect 200888 111218 200972 111454
rect 201208 111218 236652 111454
rect 236888 111218 236972 111454
rect 237208 111218 272652 111454
rect 272888 111218 272972 111454
rect 273208 111218 308652 111454
rect 308888 111218 308972 111454
rect 309208 111218 344652 111454
rect 344888 111218 344972 111454
rect 345208 111218 380652 111454
rect 380888 111218 380972 111454
rect 381208 111218 416652 111454
rect 416888 111218 416972 111454
rect 417208 111218 452652 111454
rect 452888 111218 452972 111454
rect 453208 111218 488652 111454
rect 488888 111218 488972 111454
rect 489208 111218 524652 111454
rect 524888 111218 524972 111454
rect 525208 111218 560652 111454
rect 560888 111218 560972 111454
rect 561208 111218 570292 111454
rect 570528 111218 570612 111454
rect 570848 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 607700 111454
rect -23776 111134 607700 111218
rect -23776 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 9116 111134
rect 9352 110898 9436 111134
rect 9672 110898 56652 111134
rect 56888 110898 56972 111134
rect 57208 110898 92652 111134
rect 92888 110898 92972 111134
rect 93208 110898 128652 111134
rect 128888 110898 128972 111134
rect 129208 110898 164652 111134
rect 164888 110898 164972 111134
rect 165208 110898 200652 111134
rect 200888 110898 200972 111134
rect 201208 110898 236652 111134
rect 236888 110898 236972 111134
rect 237208 110898 272652 111134
rect 272888 110898 272972 111134
rect 273208 110898 308652 111134
rect 308888 110898 308972 111134
rect 309208 110898 344652 111134
rect 344888 110898 344972 111134
rect 345208 110898 380652 111134
rect 380888 110898 380972 111134
rect 381208 110898 416652 111134
rect 416888 110898 416972 111134
rect 417208 110898 452652 111134
rect 452888 110898 452972 111134
rect 453208 110898 488652 111134
rect 488888 110898 488972 111134
rect 489208 110898 524652 111134
rect 524888 110898 524972 111134
rect 525208 110898 560652 111134
rect 560888 110898 560972 111134
rect 561208 110898 570292 111134
rect 570528 110898 570612 111134
rect 570848 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 607700 111134
rect -23776 110866 607700 110898
rect -23776 101494 607700 101526
rect -23776 101258 -23744 101494
rect -23508 101258 -23424 101494
rect -23188 101258 607112 101494
rect 607348 101258 607432 101494
rect 607668 101258 607700 101494
rect -23776 101174 607700 101258
rect -23776 100938 -23744 101174
rect -23508 100938 -23424 101174
rect -23188 100938 607112 101174
rect 607348 100938 607432 101174
rect 607668 100938 607700 101174
rect -23776 100906 607700 100938
rect -23776 97774 607700 97806
rect -23776 97538 -20634 97774
rect -20398 97538 -20314 97774
rect -20078 97538 604002 97774
rect 604238 97538 604322 97774
rect 604558 97538 607700 97774
rect -23776 97454 607700 97538
rect -23776 97218 -20634 97454
rect -20398 97218 -20314 97454
rect -20078 97218 604002 97454
rect 604238 97218 604322 97454
rect 604558 97218 607700 97454
rect -23776 97186 607700 97218
rect -23776 94054 607700 94086
rect -23776 93818 -17524 94054
rect -17288 93818 -17204 94054
rect -16968 93818 600892 94054
rect 601128 93818 601212 94054
rect 601448 93818 607700 94054
rect -23776 93734 607700 93818
rect -23776 93498 -17524 93734
rect -17288 93498 -17204 93734
rect -16968 93498 600892 93734
rect 601128 93498 601212 93734
rect 601448 93498 607700 93734
rect -23776 93466 607700 93498
rect -23776 90334 607700 90366
rect -23776 90098 -14414 90334
rect -14178 90098 -14094 90334
rect -13858 90098 597782 90334
rect 598018 90098 598102 90334
rect 598338 90098 607700 90334
rect -23776 90014 607700 90098
rect -23776 89778 -14414 90014
rect -14178 89778 -14094 90014
rect -13858 89778 597782 90014
rect 598018 89778 598102 90014
rect 598338 89778 607700 90014
rect -23776 89746 607700 89778
rect -23776 86614 607700 86646
rect -23776 86378 -11304 86614
rect -11068 86378 -10984 86614
rect -10748 86378 594672 86614
rect 594908 86378 594992 86614
rect 595228 86378 607700 86614
rect -23776 86294 607700 86378
rect -23776 86058 -11304 86294
rect -11068 86058 -10984 86294
rect -10748 86058 594672 86294
rect 594908 86058 594992 86294
rect 595228 86058 607700 86294
rect -23776 86026 607700 86058
rect -23776 82894 607700 82926
rect -23776 82658 -8194 82894
rect -7958 82658 -7874 82894
rect -7638 82658 591562 82894
rect 591798 82658 591882 82894
rect 592118 82658 607700 82894
rect -23776 82574 607700 82658
rect -23776 82338 -8194 82574
rect -7958 82338 -7874 82574
rect -7638 82338 591562 82574
rect 591798 82338 591882 82574
rect 592118 82338 607700 82574
rect -23776 82306 607700 82338
rect -23776 79174 607700 79206
rect -23776 78938 -5084 79174
rect -4848 78938 -4764 79174
rect -4528 78938 7876 79174
rect 8112 78938 8196 79174
rect 8432 78938 38032 79174
rect 38268 78938 38352 79174
rect 38588 78938 60622 79174
rect 60858 78938 159098 79174
rect 159334 78938 182032 79174
rect 182268 78938 182352 79174
rect 182588 78938 185622 79174
rect 185858 78938 284098 79174
rect 284334 78938 290032 79174
rect 290268 78938 290352 79174
rect 290588 78938 310622 79174
rect 310858 78938 409098 79174
rect 409334 78938 434032 79174
rect 434268 78938 434352 79174
rect 434588 78938 436622 79174
rect 436858 78938 535098 79174
rect 535334 78938 542032 79174
rect 542268 78938 542352 79174
rect 542588 78938 571532 79174
rect 571768 78938 571852 79174
rect 572088 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 588452 79174
rect 588688 78938 588772 79174
rect 589008 78938 607700 79174
rect -23776 78854 607700 78938
rect -23776 78618 -5084 78854
rect -4848 78618 -4764 78854
rect -4528 78618 7876 78854
rect 8112 78618 8196 78854
rect 8432 78618 38032 78854
rect 38268 78618 38352 78854
rect 38588 78618 60622 78854
rect 60858 78618 159098 78854
rect 159334 78618 182032 78854
rect 182268 78618 182352 78854
rect 182588 78618 185622 78854
rect 185858 78618 284098 78854
rect 284334 78618 290032 78854
rect 290268 78618 290352 78854
rect 290588 78618 310622 78854
rect 310858 78618 409098 78854
rect 409334 78618 434032 78854
rect 434268 78618 434352 78854
rect 434588 78618 436622 78854
rect 436858 78618 535098 78854
rect 535334 78618 542032 78854
rect 542268 78618 542352 78854
rect 542588 78618 571532 78854
rect 571768 78618 571852 78854
rect 572088 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 588452 78854
rect 588688 78618 588772 78854
rect 589008 78618 607700 78854
rect -23776 78586 607700 78618
rect -23776 75454 607700 75486
rect -23776 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 9116 75454
rect 9352 75218 9436 75454
rect 9672 75218 56652 75454
rect 56888 75218 56972 75454
rect 57208 75218 61342 75454
rect 61578 75218 158378 75454
rect 158614 75218 164652 75454
rect 164888 75218 164972 75454
rect 165208 75218 186342 75454
rect 186578 75218 283378 75454
rect 283614 75218 308652 75454
rect 308888 75218 308972 75454
rect 309208 75218 311342 75454
rect 311578 75218 408378 75454
rect 408614 75218 416652 75454
rect 416888 75218 416972 75454
rect 417208 75218 437342 75454
rect 437578 75218 534378 75454
rect 534614 75218 560652 75454
rect 560888 75218 560972 75454
rect 561208 75218 570292 75454
rect 570528 75218 570612 75454
rect 570848 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 607700 75454
rect -23776 75134 607700 75218
rect -23776 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 9116 75134
rect 9352 74898 9436 75134
rect 9672 74898 56652 75134
rect 56888 74898 56972 75134
rect 57208 74898 61342 75134
rect 61578 74898 158378 75134
rect 158614 74898 164652 75134
rect 164888 74898 164972 75134
rect 165208 74898 186342 75134
rect 186578 74898 283378 75134
rect 283614 74898 308652 75134
rect 308888 74898 308972 75134
rect 309208 74898 311342 75134
rect 311578 74898 408378 75134
rect 408614 74898 416652 75134
rect 416888 74898 416972 75134
rect 417208 74898 437342 75134
rect 437578 74898 534378 75134
rect 534614 74898 560652 75134
rect 560888 74898 560972 75134
rect 561208 74898 570292 75134
rect 570528 74898 570612 75134
rect 570848 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 607700 75134
rect -23776 74866 607700 74898
rect -23776 65494 607700 65526
rect -23776 65258 -23744 65494
rect -23508 65258 -23424 65494
rect -23188 65258 607112 65494
rect 607348 65258 607432 65494
rect 607668 65258 607700 65494
rect -23776 65174 607700 65258
rect -23776 64938 -23744 65174
rect -23508 64938 -23424 65174
rect -23188 64938 607112 65174
rect 607348 64938 607432 65174
rect 607668 64938 607700 65174
rect -23776 64906 607700 64938
rect -23776 61774 607700 61806
rect -23776 61538 -20634 61774
rect -20398 61538 -20314 61774
rect -20078 61538 604002 61774
rect 604238 61538 604322 61774
rect 604558 61538 607700 61774
rect -23776 61454 607700 61538
rect -23776 61218 -20634 61454
rect -20398 61218 -20314 61454
rect -20078 61218 604002 61454
rect 604238 61218 604322 61454
rect 604558 61218 607700 61454
rect -23776 61186 607700 61218
rect -23776 58054 607700 58086
rect -23776 57818 -17524 58054
rect -17288 57818 -17204 58054
rect -16968 57818 600892 58054
rect 601128 57818 601212 58054
rect 601448 57818 607700 58054
rect -23776 57734 607700 57818
rect -23776 57498 -17524 57734
rect -17288 57498 -17204 57734
rect -16968 57498 600892 57734
rect 601128 57498 601212 57734
rect 601448 57498 607700 57734
rect -23776 57466 607700 57498
rect -23776 54334 607700 54366
rect -23776 54098 -14414 54334
rect -14178 54098 -14094 54334
rect -13858 54098 597782 54334
rect 598018 54098 598102 54334
rect 598338 54098 607700 54334
rect -23776 54014 607700 54098
rect -23776 53778 -14414 54014
rect -14178 53778 -14094 54014
rect -13858 53778 597782 54014
rect 598018 53778 598102 54014
rect 598338 53778 607700 54014
rect -23776 53746 607700 53778
rect -23776 50614 607700 50646
rect -23776 50378 -11304 50614
rect -11068 50378 -10984 50614
rect -10748 50378 594672 50614
rect 594908 50378 594992 50614
rect 595228 50378 607700 50614
rect -23776 50294 607700 50378
rect -23776 50058 -11304 50294
rect -11068 50058 -10984 50294
rect -10748 50058 594672 50294
rect 594908 50058 594992 50294
rect 595228 50058 607700 50294
rect -23776 50026 607700 50058
rect -23776 46894 607700 46926
rect -23776 46658 -8194 46894
rect -7958 46658 -7874 46894
rect -7638 46658 591562 46894
rect 591798 46658 591882 46894
rect 592118 46658 607700 46894
rect -23776 46574 607700 46658
rect -23776 46338 -8194 46574
rect -7958 46338 -7874 46574
rect -7638 46338 591562 46574
rect 591798 46338 591882 46574
rect 592118 46338 607700 46574
rect -23776 46306 607700 46338
rect -23776 43174 607700 43206
rect -23776 42938 -5084 43174
rect -4848 42938 -4764 43174
rect -4528 42938 7876 43174
rect 8112 42938 8196 43174
rect 8432 42938 38032 43174
rect 38268 42938 38352 43174
rect 38588 42938 60622 43174
rect 60858 42938 159098 43174
rect 159334 42938 182032 43174
rect 182268 42938 182352 43174
rect 182588 42938 185622 43174
rect 185858 42938 284098 43174
rect 284334 42938 290032 43174
rect 290268 42938 290352 43174
rect 290588 42938 310622 43174
rect 310858 42938 409098 43174
rect 409334 42938 434032 43174
rect 434268 42938 434352 43174
rect 434588 42938 436622 43174
rect 436858 42938 535098 43174
rect 535334 42938 542032 43174
rect 542268 42938 542352 43174
rect 542588 42938 571532 43174
rect 571768 42938 571852 43174
rect 572088 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 588452 43174
rect 588688 42938 588772 43174
rect 589008 42938 607700 43174
rect -23776 42854 607700 42938
rect -23776 42618 -5084 42854
rect -4848 42618 -4764 42854
rect -4528 42618 7876 42854
rect 8112 42618 8196 42854
rect 8432 42618 38032 42854
rect 38268 42618 38352 42854
rect 38588 42618 60622 42854
rect 60858 42618 159098 42854
rect 159334 42618 182032 42854
rect 182268 42618 182352 42854
rect 182588 42618 185622 42854
rect 185858 42618 284098 42854
rect 284334 42618 290032 42854
rect 290268 42618 290352 42854
rect 290588 42618 310622 42854
rect 310858 42618 409098 42854
rect 409334 42618 434032 42854
rect 434268 42618 434352 42854
rect 434588 42618 436622 42854
rect 436858 42618 535098 42854
rect 535334 42618 542032 42854
rect 542268 42618 542352 42854
rect 542588 42618 571532 42854
rect 571768 42618 571852 42854
rect 572088 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 588452 42854
rect 588688 42618 588772 42854
rect 589008 42618 607700 42854
rect -23776 42586 607700 42618
rect -23776 39454 607700 39486
rect -23776 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 9116 39454
rect 9352 39218 9436 39454
rect 9672 39218 56652 39454
rect 56888 39218 56972 39454
rect 57208 39218 61342 39454
rect 61578 39218 158378 39454
rect 158614 39218 164652 39454
rect 164888 39218 164972 39454
rect 165208 39218 186342 39454
rect 186578 39218 283378 39454
rect 283614 39218 308652 39454
rect 308888 39218 308972 39454
rect 309208 39218 311342 39454
rect 311578 39218 408378 39454
rect 408614 39218 416652 39454
rect 416888 39218 416972 39454
rect 417208 39218 437342 39454
rect 437578 39218 534378 39454
rect 534614 39218 560652 39454
rect 560888 39218 560972 39454
rect 561208 39218 570292 39454
rect 570528 39218 570612 39454
rect 570848 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 607700 39454
rect -23776 39134 607700 39218
rect -23776 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 9116 39134
rect 9352 38898 9436 39134
rect 9672 38898 56652 39134
rect 56888 38898 56972 39134
rect 57208 38898 61342 39134
rect 61578 38898 158378 39134
rect 158614 38898 164652 39134
rect 164888 38898 164972 39134
rect 165208 38898 186342 39134
rect 186578 38898 283378 39134
rect 283614 38898 308652 39134
rect 308888 38898 308972 39134
rect 309208 38898 311342 39134
rect 311578 38898 408378 39134
rect 408614 38898 416652 39134
rect 416888 38898 416972 39134
rect 417208 38898 437342 39134
rect 437578 38898 534378 39134
rect 534614 38898 560652 39134
rect 560888 38898 560972 39134
rect 561208 38898 570292 39134
rect 570528 38898 570612 39134
rect 570848 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 607700 39134
rect -23776 38866 607700 38898
rect -23776 29494 607700 29526
rect -23776 29258 -23744 29494
rect -23508 29258 -23424 29494
rect -23188 29258 607112 29494
rect 607348 29258 607432 29494
rect 607668 29258 607700 29494
rect -23776 29174 607700 29258
rect -23776 28938 -23744 29174
rect -23508 28938 -23424 29174
rect -23188 28938 607112 29174
rect 607348 28938 607432 29174
rect 607668 28938 607700 29174
rect -23776 28906 607700 28938
rect -23776 25774 607700 25806
rect -23776 25538 -20634 25774
rect -20398 25538 -20314 25774
rect -20078 25538 604002 25774
rect 604238 25538 604322 25774
rect 604558 25538 607700 25774
rect -23776 25454 607700 25538
rect -23776 25218 -20634 25454
rect -20398 25218 -20314 25454
rect -20078 25218 604002 25454
rect 604238 25218 604322 25454
rect 604558 25218 607700 25454
rect -23776 25186 607700 25218
rect 61280 21244 61640 21300
rect 61280 21008 61342 21244
rect 61578 21008 61640 21244
rect 61280 20952 61640 21008
rect 62952 21244 63300 21300
rect 62952 21008 63008 21244
rect 63244 21008 63300 21244
rect 62952 20952 63300 21008
rect 187952 21244 188300 21300
rect 187952 21008 188008 21244
rect 188244 21008 188300 21244
rect 187952 20952 188300 21008
rect 311280 21244 311640 21300
rect 311280 21008 311342 21244
rect 311578 21008 311640 21244
rect 311280 20952 311640 21008
rect 312952 21244 313300 21300
rect 312952 21008 313008 21244
rect 313244 21008 313300 21244
rect 312952 20952 313300 21008
rect 438952 21244 439300 21300
rect 438952 21008 439008 21244
rect 439244 21008 439300 21244
rect 438952 20952 439300 21008
rect 62272 20564 62620 20620
rect 62272 20328 62328 20564
rect 62564 20328 62620 20564
rect 62272 20272 62620 20328
rect 185560 20564 185920 20620
rect 185560 20328 185622 20564
rect 185858 20328 185920 20564
rect 185560 20272 185920 20328
rect 187272 20564 187620 20620
rect 187272 20328 187328 20564
rect 187564 20328 187620 20564
rect 187272 20272 187620 20328
rect 312272 20564 312620 20620
rect 312272 20328 312328 20564
rect 312564 20328 312620 20564
rect 312272 20272 312620 20328
rect 436560 20564 436920 20620
rect 436560 20328 436622 20564
rect 436858 20328 436920 20564
rect 436560 20272 436920 20328
rect 438272 20564 438620 20620
rect 438272 20328 438328 20564
rect 438564 20328 438620 20564
rect 438272 20272 438620 20328
rect 62272 19834 62620 19858
rect 62272 19598 62328 19834
rect 62564 19598 62620 19834
rect 312272 19834 312620 19858
rect 62272 19574 62620 19598
rect 187952 19578 188300 19640
rect 187952 19342 188008 19578
rect 188244 19342 188300 19578
rect 312272 19598 312328 19834
rect 312564 19598 312620 19834
rect 312272 19574 312620 19598
rect 438952 19578 439300 19640
rect 187952 19280 188300 19342
rect 438952 19342 439008 19578
rect 439244 19342 439300 19578
rect 438952 19280 439300 19342
rect -23776 18334 607700 18366
rect -23776 18098 -14414 18334
rect -14178 18098 -14094 18334
rect -13858 18098 597782 18334
rect 598018 18098 598102 18334
rect 598338 18098 607700 18334
rect -23776 18014 607700 18098
rect -23776 17778 -14414 18014
rect -14178 17778 -14094 18014
rect -13858 17778 597782 18014
rect 598018 17778 598102 18014
rect 598338 17778 607700 18014
rect -23776 17746 607700 17778
rect -23776 14614 607700 14646
rect -23776 14378 -11304 14614
rect -11068 14378 -10984 14614
rect -10748 14378 594672 14614
rect 594908 14378 594992 14614
rect 595228 14378 607700 14614
rect -23776 14294 607700 14378
rect -23776 14058 -11304 14294
rect -11068 14058 -10984 14294
rect -10748 14058 594672 14294
rect 594908 14058 594992 14294
rect 595228 14058 607700 14294
rect -23776 14026 607700 14058
rect -23776 10894 607700 10926
rect -23776 10658 -8194 10894
rect -7958 10658 -7874 10894
rect -7638 10658 591562 10894
rect 591798 10658 591882 10894
rect 592118 10658 607700 10894
rect -23776 10574 607700 10658
rect -23776 10338 -8194 10574
rect -7958 10338 -7874 10574
rect -7638 10338 591562 10574
rect 591798 10338 591882 10574
rect 592118 10338 607700 10574
rect -23776 10306 607700 10338
rect 9092 9680 9696 9712
rect 9092 9444 9116 9680
rect 9352 9444 9436 9680
rect 9672 9444 9696 9680
rect 9092 9360 9696 9444
rect 9092 9124 9116 9360
rect 9352 9124 9436 9360
rect 9672 9124 9696 9360
rect 9092 9092 9696 9124
rect 56628 9680 57232 9712
rect 56628 9444 56652 9680
rect 56888 9444 56972 9680
rect 57208 9444 57232 9680
rect 56628 9360 57232 9444
rect 56628 9124 56652 9360
rect 56888 9124 56972 9360
rect 57208 9124 57232 9360
rect 56628 9092 57232 9124
rect 92628 9680 93232 9712
rect 92628 9444 92652 9680
rect 92888 9444 92972 9680
rect 93208 9444 93232 9680
rect 92628 9360 93232 9444
rect 92628 9124 92652 9360
rect 92888 9124 92972 9360
rect 93208 9124 93232 9360
rect 92628 9092 93232 9124
rect 128628 9680 129232 9712
rect 128628 9444 128652 9680
rect 128888 9444 128972 9680
rect 129208 9444 129232 9680
rect 128628 9360 129232 9444
rect 128628 9124 128652 9360
rect 128888 9124 128972 9360
rect 129208 9124 129232 9360
rect 128628 9092 129232 9124
rect 164628 9680 165232 9712
rect 164628 9444 164652 9680
rect 164888 9444 164972 9680
rect 165208 9444 165232 9680
rect 164628 9360 165232 9444
rect 164628 9124 164652 9360
rect 164888 9124 164972 9360
rect 165208 9124 165232 9360
rect 164628 9092 165232 9124
rect 200628 9680 201232 9712
rect 200628 9444 200652 9680
rect 200888 9444 200972 9680
rect 201208 9444 201232 9680
rect 200628 9360 201232 9444
rect 200628 9124 200652 9360
rect 200888 9124 200972 9360
rect 201208 9124 201232 9360
rect 200628 9092 201232 9124
rect 236628 9680 237232 9712
rect 236628 9444 236652 9680
rect 236888 9444 236972 9680
rect 237208 9444 237232 9680
rect 236628 9360 237232 9444
rect 236628 9124 236652 9360
rect 236888 9124 236972 9360
rect 237208 9124 237232 9360
rect 236628 9092 237232 9124
rect 272628 9680 273232 9712
rect 272628 9444 272652 9680
rect 272888 9444 272972 9680
rect 273208 9444 273232 9680
rect 272628 9360 273232 9444
rect 272628 9124 272652 9360
rect 272888 9124 272972 9360
rect 273208 9124 273232 9360
rect 272628 9092 273232 9124
rect 308628 9680 309232 9712
rect 308628 9444 308652 9680
rect 308888 9444 308972 9680
rect 309208 9444 309232 9680
rect 308628 9360 309232 9444
rect 308628 9124 308652 9360
rect 308888 9124 308972 9360
rect 309208 9124 309232 9360
rect 308628 9092 309232 9124
rect 344628 9680 345232 9712
rect 344628 9444 344652 9680
rect 344888 9444 344972 9680
rect 345208 9444 345232 9680
rect 344628 9360 345232 9444
rect 344628 9124 344652 9360
rect 344888 9124 344972 9360
rect 345208 9124 345232 9360
rect 344628 9092 345232 9124
rect 380628 9680 381232 9712
rect 380628 9444 380652 9680
rect 380888 9444 380972 9680
rect 381208 9444 381232 9680
rect 380628 9360 381232 9444
rect 380628 9124 380652 9360
rect 380888 9124 380972 9360
rect 381208 9124 381232 9360
rect 380628 9092 381232 9124
rect 416628 9680 417232 9712
rect 416628 9444 416652 9680
rect 416888 9444 416972 9680
rect 417208 9444 417232 9680
rect 416628 9360 417232 9444
rect 416628 9124 416652 9360
rect 416888 9124 416972 9360
rect 417208 9124 417232 9360
rect 416628 9092 417232 9124
rect 452628 9680 453232 9712
rect 452628 9444 452652 9680
rect 452888 9444 452972 9680
rect 453208 9444 453232 9680
rect 452628 9360 453232 9444
rect 452628 9124 452652 9360
rect 452888 9124 452972 9360
rect 453208 9124 453232 9360
rect 452628 9092 453232 9124
rect 488628 9680 489232 9712
rect 488628 9444 488652 9680
rect 488888 9444 488972 9680
rect 489208 9444 489232 9680
rect 488628 9360 489232 9444
rect 488628 9124 488652 9360
rect 488888 9124 488972 9360
rect 489208 9124 489232 9360
rect 488628 9092 489232 9124
rect 524628 9680 525232 9712
rect 524628 9444 524652 9680
rect 524888 9444 524972 9680
rect 525208 9444 525232 9680
rect 524628 9360 525232 9444
rect 524628 9124 524652 9360
rect 524888 9124 524972 9360
rect 525208 9124 525232 9360
rect 524628 9092 525232 9124
rect 560628 9680 561232 9712
rect 560628 9444 560652 9680
rect 560888 9444 560972 9680
rect 561208 9444 561232 9680
rect 560628 9360 561232 9444
rect 560628 9124 560652 9360
rect 560888 9124 560972 9360
rect 561208 9124 561232 9360
rect 560628 9092 561232 9124
rect 570268 9680 570872 9712
rect 570268 9444 570292 9680
rect 570528 9444 570612 9680
rect 570848 9444 570872 9680
rect 570268 9360 570872 9444
rect 570268 9124 570292 9360
rect 570528 9124 570612 9360
rect 570848 9124 570872 9360
rect 570268 9092 570872 9124
rect 7852 8440 8456 8472
rect 7852 8204 7876 8440
rect 8112 8204 8196 8440
rect 8432 8204 8456 8440
rect 7852 8120 8456 8204
rect 7852 7884 7876 8120
rect 8112 7884 8196 8120
rect 8432 7884 8456 8120
rect 7852 7852 8456 7884
rect 38008 8440 38612 8472
rect 38008 8204 38032 8440
rect 38268 8204 38352 8440
rect 38588 8204 38612 8440
rect 38008 8120 38612 8204
rect 38008 7884 38032 8120
rect 38268 7884 38352 8120
rect 38588 7884 38612 8120
rect 38008 7852 38612 7884
rect 74008 8440 74612 8472
rect 74008 8204 74032 8440
rect 74268 8204 74352 8440
rect 74588 8204 74612 8440
rect 74008 8120 74612 8204
rect 74008 7884 74032 8120
rect 74268 7884 74352 8120
rect 74588 7884 74612 8120
rect 74008 7852 74612 7884
rect 110008 8440 110612 8472
rect 110008 8204 110032 8440
rect 110268 8204 110352 8440
rect 110588 8204 110612 8440
rect 110008 8120 110612 8204
rect 110008 7884 110032 8120
rect 110268 7884 110352 8120
rect 110588 7884 110612 8120
rect 110008 7852 110612 7884
rect 146008 8440 146612 8472
rect 146008 8204 146032 8440
rect 146268 8204 146352 8440
rect 146588 8204 146612 8440
rect 146008 8120 146612 8204
rect 146008 7884 146032 8120
rect 146268 7884 146352 8120
rect 146588 7884 146612 8120
rect 146008 7852 146612 7884
rect 182008 8440 182612 8472
rect 182008 8204 182032 8440
rect 182268 8204 182352 8440
rect 182588 8204 182612 8440
rect 182008 8120 182612 8204
rect 182008 7884 182032 8120
rect 182268 7884 182352 8120
rect 182588 7884 182612 8120
rect 182008 7852 182612 7884
rect 218008 8440 218612 8472
rect 218008 8204 218032 8440
rect 218268 8204 218352 8440
rect 218588 8204 218612 8440
rect 218008 8120 218612 8204
rect 218008 7884 218032 8120
rect 218268 7884 218352 8120
rect 218588 7884 218612 8120
rect 218008 7852 218612 7884
rect 254008 8440 254612 8472
rect 254008 8204 254032 8440
rect 254268 8204 254352 8440
rect 254588 8204 254612 8440
rect 254008 8120 254612 8204
rect 254008 7884 254032 8120
rect 254268 7884 254352 8120
rect 254588 7884 254612 8120
rect 254008 7852 254612 7884
rect 290008 8440 290612 8472
rect 290008 8204 290032 8440
rect 290268 8204 290352 8440
rect 290588 8204 290612 8440
rect 290008 8120 290612 8204
rect 290008 7884 290032 8120
rect 290268 7884 290352 8120
rect 290588 7884 290612 8120
rect 290008 7852 290612 7884
rect 326008 8440 326612 8472
rect 326008 8204 326032 8440
rect 326268 8204 326352 8440
rect 326588 8204 326612 8440
rect 326008 8120 326612 8204
rect 326008 7884 326032 8120
rect 326268 7884 326352 8120
rect 326588 7884 326612 8120
rect 326008 7852 326612 7884
rect 362008 8440 362612 8472
rect 362008 8204 362032 8440
rect 362268 8204 362352 8440
rect 362588 8204 362612 8440
rect 362008 8120 362612 8204
rect 362008 7884 362032 8120
rect 362268 7884 362352 8120
rect 362588 7884 362612 8120
rect 362008 7852 362612 7884
rect 398008 8440 398612 8472
rect 398008 8204 398032 8440
rect 398268 8204 398352 8440
rect 398588 8204 398612 8440
rect 398008 8120 398612 8204
rect 398008 7884 398032 8120
rect 398268 7884 398352 8120
rect 398588 7884 398612 8120
rect 398008 7852 398612 7884
rect 434008 8440 434612 8472
rect 434008 8204 434032 8440
rect 434268 8204 434352 8440
rect 434588 8204 434612 8440
rect 434008 8120 434612 8204
rect 434008 7884 434032 8120
rect 434268 7884 434352 8120
rect 434588 7884 434612 8120
rect 434008 7852 434612 7884
rect 470008 8440 470612 8472
rect 470008 8204 470032 8440
rect 470268 8204 470352 8440
rect 470588 8204 470612 8440
rect 470008 8120 470612 8204
rect 470008 7884 470032 8120
rect 470268 7884 470352 8120
rect 470588 7884 470612 8120
rect 470008 7852 470612 7884
rect 506008 8440 506612 8472
rect 506008 8204 506032 8440
rect 506268 8204 506352 8440
rect 506588 8204 506612 8440
rect 506008 8120 506612 8204
rect 506008 7884 506032 8120
rect 506268 7884 506352 8120
rect 506588 7884 506612 8120
rect 506008 7852 506612 7884
rect 542008 8440 542612 8472
rect 542008 8204 542032 8440
rect 542268 8204 542352 8440
rect 542588 8204 542612 8440
rect 542008 8120 542612 8204
rect 542008 7884 542032 8120
rect 542268 7884 542352 8120
rect 542588 7884 542612 8120
rect 542008 7852 542612 7884
rect 571508 8440 572112 8472
rect 571508 8204 571532 8440
rect 571768 8204 571852 8440
rect 572088 8204 572112 8440
rect 571508 8120 572112 8204
rect 571508 7884 571532 8120
rect 571768 7884 571852 8120
rect 572088 7884 572112 8120
rect 571508 7852 572112 7884
rect -23776 7174 607700 7206
rect -23776 6938 -5084 7174
rect -4848 6938 -4764 7174
rect -4528 6938 7876 7174
rect 8112 6938 8196 7174
rect 8432 6938 571532 7174
rect 571768 6938 571852 7174
rect 572088 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 588452 7174
rect 588688 6938 588772 7174
rect 589008 6938 607700 7174
rect -23776 6854 607700 6938
rect -23776 6618 -5084 6854
rect -4848 6618 -4764 6854
rect -4528 6618 7876 6854
rect 8112 6618 8196 6854
rect 8432 6618 571532 6854
rect 571768 6618 571852 6854
rect 572088 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 588452 6854
rect 588688 6618 588772 6854
rect 589008 6618 607700 6854
rect -23776 6586 607700 6618
rect -23776 3454 607700 3486
rect -23776 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 607700 3454
rect -23776 3134 607700 3218
rect -23776 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 607700 3134
rect -23776 2866 607700 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -5116 -3456 589040 -3424
rect -5116 -3692 -5084 -3456
rect -4848 -3692 -4764 -3456
rect -4528 -3692 581546 -3456
rect 581782 -3692 581866 -3456
rect 582102 -3692 588452 -3456
rect 588688 -3692 588772 -3456
rect 589008 -3692 589040 -3456
rect -5116 -3776 589040 -3692
rect -5116 -4012 -5084 -3776
rect -4848 -4012 -4764 -3776
rect -4528 -4012 581546 -3776
rect 581782 -4012 581866 -3776
rect 582102 -4012 588452 -3776
rect 588688 -4012 588772 -3776
rect 589008 -4012 589040 -3776
rect -5116 -4044 589040 -4012
rect -8226 -6566 592150 -6534
rect -8226 -6802 -8194 -6566
rect -7958 -6802 -7874 -6566
rect -7638 -6802 591562 -6566
rect 591798 -6802 591882 -6566
rect 592118 -6802 592150 -6566
rect -8226 -6886 592150 -6802
rect -8226 -7122 -8194 -6886
rect -7958 -7122 -7874 -6886
rect -7638 -7122 591562 -6886
rect 591798 -7122 591882 -6886
rect 592118 -7122 592150 -6886
rect -8226 -7154 592150 -7122
rect -11336 -9676 595260 -9644
rect -11336 -9912 -11304 -9676
rect -11068 -9912 -10984 -9676
rect -10748 -9912 594672 -9676
rect 594908 -9912 594992 -9676
rect 595228 -9912 595260 -9676
rect -11336 -9996 595260 -9912
rect -11336 -10232 -11304 -9996
rect -11068 -10232 -10984 -9996
rect -10748 -10232 594672 -9996
rect 594908 -10232 594992 -9996
rect 595228 -10232 595260 -9996
rect -11336 -10264 595260 -10232
rect -14446 -12786 598370 -12754
rect -14446 -13022 -14414 -12786
rect -14178 -13022 -14094 -12786
rect -13858 -13022 597782 -12786
rect 598018 -13022 598102 -12786
rect 598338 -13022 598370 -12786
rect -14446 -13106 598370 -13022
rect -14446 -13342 -14414 -13106
rect -14178 -13342 -14094 -13106
rect -13858 -13342 597782 -13106
rect 598018 -13342 598102 -13106
rect 598338 -13342 598370 -13106
rect -14446 -13374 598370 -13342
rect -17556 -15896 601480 -15864
rect -17556 -16132 -17524 -15896
rect -17288 -16132 -17204 -15896
rect -16968 -16132 600892 -15896
rect 601128 -16132 601212 -15896
rect 601448 -16132 601480 -15896
rect -17556 -16216 601480 -16132
rect -17556 -16452 -17524 -16216
rect -17288 -16452 -17204 -16216
rect -16968 -16452 600892 -16216
rect 601128 -16452 601212 -16216
rect 601448 -16452 601480 -16216
rect -17556 -16484 601480 -16452
rect -20666 -19006 604590 -18974
rect -20666 -19242 -20634 -19006
rect -20398 -19242 -20314 -19006
rect -20078 -19242 604002 -19006
rect 604238 -19242 604322 -19006
rect 604558 -19242 604590 -19006
rect -20666 -19326 604590 -19242
rect -20666 -19562 -20634 -19326
rect -20398 -19562 -20314 -19326
rect -20078 -19562 604002 -19326
rect 604238 -19562 604322 -19326
rect 604558 -19562 604590 -19326
rect -20666 -19594 604590 -19562
rect -23776 -22116 607700 -22084
rect -23776 -22352 -23744 -22116
rect -23508 -22352 -23424 -22116
rect -23188 -22352 607112 -22116
rect 607348 -22352 607432 -22116
rect 607668 -22352 607700 -22116
rect -23776 -22436 607700 -22352
rect -23776 -22672 -23744 -22436
rect -23508 -22672 -23424 -22436
rect -23188 -22672 607112 -22436
rect 607348 -22672 607432 -22436
rect 607668 -22672 607700 -22436
rect -23776 -22704 607700 -22672
use user_proj_example  mprj
timestamp 0
transform 1 0 4000 0 1 4000
box 0 0 571964 694008
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 2866 607700 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 38866 607700 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 74866 607700 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 110866 607700 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 146866 607700 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 182866 607700 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 218866 607700 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 254866 607700 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 290866 607700 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 326866 607700 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 362866 607700 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 398866 607700 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 434866 607700 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 470866 607700 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 506866 607700 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 542866 607700 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 578866 607700 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 614866 607700 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 650866 607700 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -23776 686866 607700 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -8226 -7154 -7606 711090 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8226 -7154 592150 -6534 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8226 710470 592150 711090 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 591530 -7154 592150 711090 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 10306 607700 10926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 46306 607700 46926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 82306 607700 82926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 118306 607700 118926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 154306 607700 154926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 190306 607700 190926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 226306 607700 226926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 262306 607700 262926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 298306 607700 298926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 334306 607700 334926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 370306 607700 370926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 406306 607700 406926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 442306 607700 442926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 478306 607700 478926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 514306 607700 514926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 550306 607700 550926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 586306 607700 586926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 622306 607700 622926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 658306 607700 658926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -23776 694306 607700 694926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -14446 -13374 -13826 717310 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -14446 -13374 598370 -12754 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -14446 716690 598370 717310 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 597750 -13374 598370 717310 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 17746 607700 18366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 53746 607700 54366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 89746 607700 90366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 125746 607700 126366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 161746 607700 162366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 197746 607700 198366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 233746 607700 234366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 269746 607700 270366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 305746 607700 306366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 341746 607700 342366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 377746 607700 378366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 413746 607700 414366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 449746 607700 450366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 485746 607700 486366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 521746 607700 522366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 557746 607700 558366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 593746 607700 594366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 629746 607700 630366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -23776 665746 607700 666366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -20666 -19594 -20046 723530 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -20666 -19594 604590 -18974 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -20666 722910 604590 723530 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 603970 -19594 604590 723530 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 25186 607700 25806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 61186 607700 61806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 97186 607700 97806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 133186 607700 133806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 169186 607700 169806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 205186 607700 205806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 241186 607700 241806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 277186 607700 277806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 313186 607700 313806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 349186 607700 349806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 385186 607700 385806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 421186 607700 421806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 457186 607700 457806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 493186 607700 493806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 529186 607700 529806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 565186 607700 565806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 601186 607700 601806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 637186 607700 637806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -23776 673186 607700 673806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -17556 -16484 -16936 720420 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -17556 -16484 601480 -15864 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -17556 719800 601480 720420 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 600860 -16484 601480 720420 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 57466 607700 58086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 93466 607700 94086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 129466 607700 130086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 165466 607700 166086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 201466 607700 202086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 237466 607700 238086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 273466 607700 274086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 309466 607700 310086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 345466 607700 346086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 381466 607700 382086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 417466 607700 418086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 453466 607700 454086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 489466 607700 490086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 525466 607700 526086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 561466 607700 562086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 597466 607700 598086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 633466 607700 634086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -23776 669466 607700 670086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -23776 -22704 -23156 726640 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 -22704 607700 -22084 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 726020 607700 726640 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 607080 -22704 607700 726640 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 28906 607700 29526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 64906 607700 65526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 100906 607700 101526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 136906 607700 137526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 172906 607700 173526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 208906 607700 209526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 244906 607700 245526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 280906 607700 281526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 316906 607700 317526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 352906 607700 353526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 388906 607700 389526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 424906 607700 425526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 460906 607700 461526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 496906 607700 497526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 532906 607700 533526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 568906 607700 569526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 604906 607700 605526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 640906 607700 641526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -23776 676906 607700 677526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -5116 -4044 -4496 707980 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -5116 -4044 589040 -3424 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -5116 707360 589040 707980 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 588420 -4044 589040 707980 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 581514 -22704 582134 726640 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 6586 607700 7206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 42586 607700 43206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 78586 607700 79206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 114586 607700 115206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 150586 607700 151206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 186586 607700 187206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 222586 607700 223206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 258586 607700 259206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 294586 607700 295206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 330586 607700 331206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 366586 607700 367206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 402586 607700 403206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 438586 607700 439206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 474586 607700 475206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 510586 607700 511206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 546586 607700 547206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 582586 607700 583206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 618586 607700 619206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 654586 607700 655206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -23776 690586 607700 691206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -11336 -10264 -10716 714200 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -11336 -10264 595260 -9644 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -11336 713580 595260 714200 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 594640 -10264 595260 714200 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 14026 607700 14646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 50026 607700 50646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 86026 607700 86646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 122026 607700 122646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 158026 607700 158646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 194026 607700 194646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 230026 607700 230646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 266026 607700 266646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 302026 607700 302646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 338026 607700 338646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 374026 607700 374646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 410026 607700 410646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 446026 607700 446646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 482026 607700 482646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 518026 607700 518646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 554026 607700 554646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 590026 607700 590646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 626026 607700 626646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 662026 607700 662646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -23776 698026 607700 698646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
rlabel via4 570730 692358 570730 692358 0 vccd1
rlabel metal5 291962 694616 291962 694616 0 vccd2
rlabel metal5 291962 666056 291962 666056 0 vdda1
rlabel metal5 291962 673496 291962 673496 0 vdda2
rlabel metal5 291962 669776 291962 669776 0 vssa1
rlabel metal5 291962 677216 291962 677216 0 vssa2
rlabel via4 571970 693598 571970 693598 0 vssd1
rlabel metal5 291962 698336 291962 698336 0 vssd2
rlabel metal2 580198 284920 580198 284920 0 analog_io[0]
rlabel metal2 445186 698064 445186 698064 0 analog_io[10]
rlabel metal2 379774 698064 379774 698064 0 analog_io[11]
rlabel metal2 314454 698064 314454 698064 0 analog_io[12]
rlabel metal2 249042 698064 249042 698064 0 analog_io[13]
rlabel metal2 183722 698064 183722 698064 0 analog_io[14]
rlabel metal2 118402 698064 118402 698064 0 analog_io[15]
rlabel metal2 56810 702076 56810 702076 0 analog_io[16]
rlabel metal3 3780 697948 3780 697948 0 analog_io[17]
rlabel metal3 3711 645488 3711 645488 0 analog_io[18]
rlabel metal3 3711 593150 3711 593150 0 analog_io[19]
rlabel metal2 579600 337892 579600 337892 0 analog_io[1]
rlabel metal3 3711 540812 3711 540812 0 analog_io[20]
rlabel metal3 3711 488474 3711 488474 0 analog_io[21]
rlabel metal3 3734 436014 3734 436014 0 analog_io[22]
rlabel metal3 3734 383676 3734 383676 0 analog_io[23]
rlabel metal3 3734 331338 3734 331338 0 analog_io[24]
rlabel metal3 3734 279000 3734 279000 0 analog_io[25]
rlabel metal3 3734 226662 3734 226662 0 analog_io[26]
rlabel metal3 3734 174202 3734 174202 0 analog_io[27]
rlabel metal3 3734 121864 3734 121864 0 analog_io[28]
rlabel metal3 583556 391408 583556 391408 0 analog_io[2]
rlabel metal3 580183 444788 580183 444788 0 analog_io[3]
rlabel metal3 576165 497868 576165 497868 0 analog_io[4]
rlabel metal3 576165 551182 576165 551182 0 analog_io[5]
rlabel metal3 579692 604316 579692 604316 0 analog_io[6]
rlabel metal3 583556 657696 583556 657696 0 analog_io[7]
rlabel metal2 575918 698064 575918 698064 0 analog_io[8]
rlabel metal2 510506 698064 510506 698064 0 analog_io[9]
rlabel metal2 576886 4845 576886 4845 0 io_in[0]
rlabel metal3 580183 458116 580183 458116 0 io_in[10]
rlabel metal3 576165 511166 576165 511166 0 io_in[11]
rlabel metal3 579692 564400 579692 564400 0 io_in[12]
rlabel metal3 583556 617780 583556 617780 0 io_in[13]
rlabel metal3 583556 671092 583556 671092 0 io_in[14]
rlabel metal2 559542 698064 559542 698064 0 io_in[15]
rlabel metal2 494222 698064 494222 698064 0 io_in[16]
rlabel metal2 428810 698064 428810 698064 0 io_in[17]
rlabel metal2 365010 701974 365010 701974 0 io_in[18]
rlabel metal2 298078 698064 298078 698064 0 io_in[19]
rlabel metal2 578358 44625 578358 44625 0 io_in[1]
rlabel metal2 232758 698064 232758 698064 0 io_in[20]
rlabel metal2 167346 698064 167346 698064 0 io_in[21]
rlabel metal2 102026 698064 102026 698064 0 io_in[22]
rlabel metal2 36706 698064 36706 698064 0 io_in[23]
rlabel metal3 3711 684772 3711 684772 0 io_in[24]
rlabel metal3 3711 632434 3711 632434 0 io_in[25]
rlabel metal3 3711 580096 3711 580096 0 io_in[26]
rlabel metal3 3711 527758 3711 527758 0 io_in[27]
rlabel metal3 3711 475298 3711 475298 0 io_in[28]
rlabel metal3 3734 422960 3734 422960 0 io_in[29]
rlabel metal2 579600 84252 579600 84252 0 io_in[2]
rlabel metal3 3734 370622 3734 370622 0 io_in[30]
rlabel metal3 3734 318284 3734 318284 0 io_in[31]
rlabel metal3 3734 265946 3734 265946 0 io_in[32]
rlabel metal3 3734 213486 3734 213486 0 io_in[33]
rlabel metal3 3711 161148 3711 161148 0 io_in[34]
rlabel metal3 3711 108810 3711 108810 0 io_in[35]
rlabel metal3 3734 69526 3734 69526 0 io_in[36]
rlabel metal3 3711 30242 3711 30242 0 io_in[37]
rlabel metal2 579600 124372 579600 124372 0 io_in[3]
rlabel metal2 579600 164356 579600 164356 0 io_in[4]
rlabel metal2 579600 204340 579600 204340 0 io_in[5]
rlabel metal2 580198 245004 580198 245004 0 io_in[6]
rlabel metal2 579600 297772 579600 297772 0 io_in[7]
rlabel metal2 579554 351492 579554 351492 0 io_in[8]
rlabel metal3 583556 404668 583556 404668 0 io_in[9]
rlabel metal2 579600 30940 579600 30940 0 io_oeb[0]
rlabel metal3 576165 484570 576165 484570 0 io_oeb[10]
rlabel metal3 576165 537884 576165 537884 0 io_oeb[11]
rlabel metal3 580183 590988 580183 590988 0 io_oeb[12]
rlabel metal3 582230 644028 582230 644028 0 io_oeb[13]
rlabel metal2 580198 697731 580198 697731 0 io_oeb[14]
rlabel metal2 526882 698064 526882 698064 0 io_oeb[15]
rlabel metal2 461470 698064 461470 698064 0 io_oeb[16]
rlabel metal2 396150 698064 396150 698064 0 io_oeb[17]
rlabel metal2 330738 698064 330738 698064 0 io_oeb[18]
rlabel metal2 265418 698064 265418 698064 0 io_oeb[19]
rlabel metal2 579600 70924 579600 70924 0 io_oeb[1]
rlabel metal2 200098 698064 200098 698064 0 io_oeb[20]
rlabel metal2 134686 698064 134686 698064 0 io_oeb[21]
rlabel metal2 69366 698064 69366 698064 0 io_oeb[22]
rlabel metal2 4046 698081 4046 698081 0 io_oeb[23]
rlabel metal3 3711 658664 3711 658664 0 io_oeb[24]
rlabel metal3 3711 606204 3711 606204 0 io_oeb[25]
rlabel metal3 3711 553866 3711 553866 0 io_oeb[26]
rlabel metal3 3711 501528 3711 501528 0 io_oeb[27]
rlabel metal3 3711 449190 3711 449190 0 io_oeb[28]
rlabel metal3 3734 396852 3734 396852 0 io_oeb[29]
rlabel metal2 579600 110908 579600 110908 0 io_oeb[2]
rlabel metal3 1878 345372 1878 345372 0 io_oeb[30]
rlabel metal3 3734 292054 3734 292054 0 io_oeb[31]
rlabel metal3 3734 239716 3734 239716 0 io_oeb[32]
rlabel metal3 3826 187378 3826 187378 0 io_oeb[33]
rlabel metal3 3711 135040 3711 135040 0 io_oeb[34]
rlabel metal3 3711 82580 3711 82580 0 io_oeb[35]
rlabel metal3 3734 43296 3734 43296 0 io_oeb[36]
rlabel metal3 3895 4134 3895 4134 0 io_oeb[37]
rlabel metal3 582230 152660 582230 152660 0 io_oeb[3]
rlabel metal2 579600 191012 579600 191012 0 io_oeb[4]
rlabel metal2 579600 231132 579600 231132 0 io_oeb[5]
rlabel metal2 579600 271116 579600 271116 0 io_oeb[6]
rlabel metal2 580198 324836 580198 324836 0 io_oeb[7]
rlabel metal3 579508 378012 579508 378012 0 io_oeb[8]
rlabel metal3 583556 431324 583556 431324 0 io_oeb[9]
rlabel metal2 579600 17612 579600 17612 0 io_out[0]
rlabel metal3 580183 471444 580183 471444 0 io_out[10]
rlabel metal3 576165 524586 576165 524586 0 io_out[11]
rlabel metal3 580183 577660 580183 577660 0 io_out[12]
rlabel metal3 583556 631108 583556 631108 0 io_out[13]
rlabel metal2 579600 684692 579600 684692 0 io_out[14]
rlabel metal2 543166 698064 543166 698064 0 io_out[15]
rlabel metal2 477846 698064 477846 698064 0 io_out[16]
rlabel metal2 412434 698064 412434 698064 0 io_out[17]
rlabel metal2 347114 698064 347114 698064 0 io_out[18]
rlabel metal2 281794 698064 281794 698064 0 io_out[19]
rlabel metal2 579600 57596 579600 57596 0 io_out[1]
rlabel metal2 216382 698064 216382 698064 0 io_out[20]
rlabel metal2 154146 702076 154146 702076 0 io_out[21]
rlabel metal2 85742 698064 85742 698064 0 io_out[22]
rlabel metal2 20330 698064 20330 698064 0 io_out[23]
rlabel metal3 3711 671718 3711 671718 0 io_out[24]
rlabel metal3 3711 619380 3711 619380 0 io_out[25]
rlabel metal3 3711 566920 3711 566920 0 io_out[26]
rlabel metal3 3711 514582 3711 514582 0 io_out[27]
rlabel metal3 3711 462244 3711 462244 0 io_out[28]
rlabel metal3 3734 409906 3734 409906 0 io_out[29]
rlabel metal2 579600 97580 579600 97580 0 io_out[2]
rlabel metal3 3734 357568 3734 357568 0 io_out[30]
rlabel metal3 3734 305108 3734 305108 0 io_out[31]
rlabel metal3 3734 252770 3734 252770 0 io_out[32]
rlabel metal3 3734 200432 3734 200432 0 io_out[33]
rlabel metal3 3734 148094 3734 148094 0 io_out[34]
rlabel metal3 3734 95756 3734 95756 0 io_out[35]
rlabel metal3 3711 56472 3711 56472 0 io_out[36]
rlabel metal3 3711 17188 3711 17188 0 io_out[37]
rlabel metal2 579600 137564 579600 137564 0 io_out[3]
rlabel metal2 579600 177684 579600 177684 0 io_out[4]
rlabel metal2 579600 217668 579600 217668 0 io_out[5]
rlabel metal2 578910 257737 578910 257737 0 io_out[6]
rlabel metal2 579600 311100 579600 311100 0 io_out[7]
rlabel metal3 583556 364684 583556 364684 0 io_out[8]
rlabel metal3 579692 418200 579692 418200 0 io_out[9]
rlabel metal2 125902 840 125902 840 0 la_data_in[0]
rlabel metal2 480562 772 480562 772 0 la_data_in[100]
rlabel metal2 484058 1588 484058 1588 0 la_data_in[101]
rlabel metal2 487455 340 487455 340 0 la_data_in[102]
rlabel metal2 485530 2397 485530 2397 0 la_data_in[103]
rlabel metal2 489026 2499 489026 2499 0 la_data_in[104]
rlabel metal2 498226 772 498226 772 0 la_data_in[105]
rlabel metal2 501814 670 501814 670 0 la_data_in[106]
rlabel via1 505586 51 505586 51 0 la_data_in[107]
rlabel metal2 508898 670 508898 670 0 la_data_in[108]
rlabel metal2 506322 1887 506322 1887 0 la_data_in[109]
rlabel metal2 161598 2040 161598 2040 0 la_data_in[10]
rlabel metal2 515883 340 515883 340 0 la_data_in[110]
rlabel metal2 519570 772 519570 772 0 la_data_in[111]
rlabel via1 523250 51 523250 51 0 la_data_in[112]
rlabel metal2 526654 670 526654 670 0 la_data_in[113]
rlabel metal2 523802 2431 523802 2431 0 la_data_in[114]
rlabel metal2 527298 2499 527298 2499 0 la_data_in[115]
rlabel metal2 537234 738 537234 738 0 la_data_in[116]
rlabel metal2 540631 340 540631 340 0 la_data_in[117]
rlabel via1 544594 323 544594 323 0 la_data_in[118]
rlabel metal2 541190 2227 541190 2227 0 la_data_in[119]
rlabel metal2 164910 2047 164910 2047 0 la_data_in[11]
rlabel metal2 544686 2091 544686 2091 0 la_data_in[120]
rlabel metal2 554990 772 554990 772 0 la_data_in[121]
rlabel metal2 558578 840 558578 840 0 la_data_in[122]
rlabel via1 562258 85 562258 85 0 la_data_in[123]
rlabel metal2 565662 772 565662 772 0 la_data_in[124]
rlabel metal2 562074 2499 562074 2499 0 la_data_in[125]
rlabel metal2 565478 1921 565478 1921 0 la_data_in[126]
rlabel metal2 576334 772 576334 772 0 la_data_in[127]
rlabel metal2 168406 2047 168406 2047 0 la_data_in[12]
rlabel metal2 172139 340 172139 340 0 la_data_in[13]
rlabel metal2 175635 340 175635 340 0 la_data_in[14]
rlabel metal2 179078 2047 179078 2047 0 la_data_in[15]
rlabel metal2 182574 2047 182574 2047 0 la_data_in[16]
rlabel metal2 186162 2047 186162 2047 0 la_data_in[17]
rlabel metal2 189750 2047 189750 2047 0 la_data_in[18]
rlabel metal2 193246 2047 193246 2047 0 la_data_in[19]
rlabel metal2 129398 840 129398 840 0 la_data_in[1]
rlabel metal2 196834 2047 196834 2047 0 la_data_in[20]
rlabel metal2 200098 3869 200098 3869 0 la_data_in[21]
rlabel metal2 203773 340 203773 340 0 la_data_in[22]
rlabel metal2 207269 340 207269 340 0 la_data_in[23]
rlabel metal2 211002 2047 211002 2047 0 la_data_in[24]
rlabel metal2 214498 2047 214498 2047 0 la_data_in[25]
rlabel metal2 217849 340 217849 340 0 la_data_in[26]
rlabel metal2 221345 340 221345 340 0 la_data_in[27]
rlabel metal2 225170 2064 225170 2064 0 la_data_in[28]
rlabel metal2 228521 340 228521 340 0 la_data_in[29]
rlabel metal2 132986 840 132986 840 0 la_data_in[2]
rlabel metal2 232254 2064 232254 2064 0 la_data_in[30]
rlabel metal2 235842 2047 235842 2047 0 la_data_in[31]
rlabel metal2 238370 3886 238370 3886 0 la_data_in[32]
rlabel metal2 242926 2064 242926 2064 0 la_data_in[33]
rlabel metal2 246422 2064 246422 2064 0 la_data_in[34]
rlabel metal2 250010 1588 250010 1588 0 la_data_in[35]
rlabel metal2 253506 2064 253506 2064 0 la_data_in[36]
rlabel metal2 257094 2064 257094 2064 0 la_data_in[37]
rlabel metal2 260682 2098 260682 2098 0 la_data_in[38]
rlabel metal2 264178 2064 264178 2064 0 la_data_in[39]
rlabel metal2 136482 806 136482 806 0 la_data_in[3]
rlabel metal2 267766 840 267766 840 0 la_data_in[40]
rlabel metal2 271262 2064 271262 2064 0 la_data_in[41]
rlabel metal2 274850 840 274850 840 0 la_data_in[42]
rlabel metal2 276734 3886 276734 3886 0 la_data_in[43]
rlabel metal2 281934 840 281934 840 0 la_data_in[44]
rlabel metal2 285430 2064 285430 2064 0 la_data_in[45]
rlabel metal2 289018 2064 289018 2064 0 la_data_in[46]
rlabel metal2 292606 466 292606 466 0 la_data_in[47]
rlabel metal2 296102 2064 296102 2064 0 la_data_in[48]
rlabel metal2 299690 840 299690 840 0 la_data_in[49]
rlabel metal2 140070 806 140070 806 0 la_data_in[4]
rlabel metal2 303186 2064 303186 2064 0 la_data_in[50]
rlabel metal2 306774 466 306774 466 0 la_data_in[51]
rlabel metal2 310270 2064 310270 2064 0 la_data_in[52]
rlabel metal2 313858 772 313858 772 0 la_data_in[53]
rlabel metal2 315054 3281 315054 3281 0 la_data_in[54]
rlabel metal2 320942 806 320942 806 0 la_data_in[55]
rlabel metal2 324438 840 324438 840 0 la_data_in[56]
rlabel metal2 328026 840 328026 840 0 la_data_in[57]
rlabel metal2 331614 840 331614 840 0 la_data_in[58]
rlabel metal2 335110 840 335110 840 0 la_data_in[59]
rlabel metal2 143566 2047 143566 2047 0 la_data_in[5]
rlabel metal2 338698 840 338698 840 0 la_data_in[60]
rlabel metal2 342194 840 342194 840 0 la_data_in[61]
rlabel metal2 345782 534 345782 534 0 la_data_in[62]
rlabel metal2 349278 534 349278 534 0 la_data_in[63]
rlabel metal2 352866 840 352866 840 0 la_data_in[64]
rlabel metal2 353234 2533 353234 2533 0 la_data_in[65]
rlabel metal2 359950 840 359950 840 0 la_data_in[66]
rlabel metal2 363538 738 363538 738 0 la_data_in[67]
rlabel metal2 367034 806 367034 806 0 la_data_in[68]
rlabel metal2 370622 840 370622 840 0 la_data_in[69]
rlabel metal2 147391 340 147391 340 0 la_data_in[6]
rlabel metal2 370714 2533 370714 2533 0 la_data_in[70]
rlabel metal2 377706 670 377706 670 0 la_data_in[71]
rlabel metal2 381202 806 381202 806 0 la_data_in[72]
rlabel metal2 384790 772 384790 772 0 la_data_in[73]
rlabel metal2 388286 602 388286 602 0 la_data_in[74]
rlabel metal2 391874 806 391874 806 0 la_data_in[75]
rlabel metal2 391598 2295 391598 2295 0 la_data_in[76]
rlabel metal2 398958 840 398958 840 0 la_data_in[77]
rlabel metal2 402546 806 402546 806 0 la_data_in[78]
rlabel via1 406226 51 406226 51 0 la_data_in[79]
rlabel metal2 150887 340 150887 340 0 la_data_in[7]
rlabel metal2 409630 840 409630 840 0 la_data_in[80]
rlabel metal2 408986 2431 408986 2431 0 la_data_in[81]
rlabel metal2 412482 1989 412482 1989 0 la_data_in[82]
rlabel metal2 420210 840 420210 840 0 la_data_in[83]
rlabel metal2 423607 340 423607 340 0 la_data_in[84]
rlabel metal2 427294 670 427294 670 0 la_data_in[85]
rlabel metal2 430882 772 430882 772 0 la_data_in[86]
rlabel metal2 429870 2295 429870 2295 0 la_data_in[87]
rlabel metal2 437966 551 437966 551 0 la_data_in[88]
rlabel metal2 441554 738 441554 738 0 la_data_in[89]
rlabel metal2 154238 840 154238 840 0 la_data_in[8]
rlabel metal2 445050 1588 445050 1588 0 la_data_in[90]
rlabel metal2 448447 340 448447 340 0 la_data_in[91]
rlabel metal2 447258 2397 447258 2397 0 la_data_in[92]
rlabel metal2 450754 2499 450754 2499 0 la_data_in[93]
rlabel metal2 459218 738 459218 738 0 la_data_in[94]
rlabel metal2 462615 340 462615 340 0 la_data_in[95]
rlabel metal2 466302 738 466302 738 0 la_data_in[96]
rlabel metal2 469890 670 469890 670 0 la_data_in[97]
rlabel metal2 468142 2533 468142 2533 0 la_data_in[98]
rlabel metal2 476783 340 476783 340 0 la_data_in[99]
rlabel metal2 158063 340 158063 340 0 la_data_in[9]
rlabel metal2 127006 755 127006 755 0 la_data_out[0]
rlabel metal2 481567 340 481567 340 0 la_data_out[100]
rlabel metal2 485063 340 485063 340 0 la_data_out[101]
rlabel metal2 488842 636 488842 636 0 la_data_out[102]
rlabel metal2 486726 2431 486726 2431 0 la_data_out[103]
rlabel metal2 495735 340 495735 340 0 la_data_out[104]
rlabel metal2 499422 738 499422 738 0 la_data_out[105]
rlabel metal2 503010 840 503010 840 0 la_data_out[106]
rlabel metal2 506506 738 506506 738 0 la_data_out[107]
rlabel metal2 504114 2533 504114 2533 0 la_data_out[108]
rlabel metal2 507518 2091 507518 2091 0 la_data_out[109]
rlabel metal2 162518 840 162518 840 0 la_data_out[10]
rlabel metal2 517178 806 517178 806 0 la_data_out[110]
rlabel metal2 520766 704 520766 704 0 la_data_out[111]
rlabel metal2 524071 340 524071 340 0 la_data_out[112]
rlabel metal2 527850 704 527850 704 0 la_data_out[113]
rlabel metal2 524998 1921 524998 1921 0 la_data_out[114]
rlabel metal2 528494 1989 528494 1989 0 la_data_out[115]
rlabel metal2 538430 772 538430 772 0 la_data_out[116]
rlabel metal2 542117 340 542117 340 0 la_data_out[117]
rlabel metal2 545514 738 545514 738 0 la_data_out[118]
rlabel metal2 542294 2533 542294 2533 0 la_data_out[119]
rlabel metal2 166297 340 166297 340 0 la_data_out[11]
rlabel metal2 545882 2023 545882 2023 0 la_data_out[120]
rlabel metal2 556186 704 556186 704 0 la_data_out[121]
rlabel metal2 559774 738 559774 738 0 la_data_out[122]
rlabel metal2 563270 466 563270 466 0 la_data_out[123]
rlabel metal2 566858 704 566858 704 0 la_data_out[124]
rlabel metal2 563178 2193 563178 2193 0 la_data_out[125]
rlabel metal2 566674 2091 566674 2091 0 la_data_out[126]
rlabel metal2 577438 806 577438 806 0 la_data_out[127]
rlabel metal2 169793 340 169793 340 0 la_data_out[12]
rlabel metal2 173190 2047 173190 2047 0 la_data_out[13]
rlabel metal2 176686 2047 176686 2047 0 la_data_out[14]
rlabel metal2 180373 204 180373 204 0 la_data_out[15]
rlabel metal2 183869 204 183869 204 0 la_data_out[16]
rlabel metal2 187358 2047 187358 2047 0 la_data_out[17]
rlabel metal2 190854 2047 190854 2047 0 la_data_out[18]
rlabel metal2 194442 2047 194442 2047 0 la_data_out[19]
rlabel metal2 130594 840 130594 840 0 la_data_out[1]
rlabel metal2 197938 2047 197938 2047 0 la_data_out[20]
rlabel metal2 201427 340 201427 340 0 la_data_out[21]
rlabel metal2 205114 2047 205114 2047 0 la_data_out[22]
rlabel metal2 208610 2047 208610 2047 0 la_data_out[23]
rlabel metal2 211961 340 211961 340 0 la_data_out[24]
rlabel metal2 215457 340 215457 340 0 la_data_out[25]
rlabel metal2 219282 2047 219282 2047 0 la_data_out[26]
rlabel metal2 222778 2064 222778 2064 0 la_data_out[27]
rlabel metal2 226129 340 226129 340 0 la_data_out[28]
rlabel metal2 229625 340 229625 340 0 la_data_out[29]
rlabel metal2 134182 2047 134182 2047 0 la_data_out[2]
rlabel metal2 233450 2064 233450 2064 0 la_data_out[30]
rlabel metal2 236801 340 236801 340 0 la_data_out[31]
rlabel metal2 240534 2064 240534 2064 0 la_data_out[32]
rlabel metal2 244122 2047 244122 2047 0 la_data_out[33]
rlabel metal2 247618 2064 247618 2064 0 la_data_out[34]
rlabel metal2 251206 2064 251206 2064 0 la_data_out[35]
rlabel metal2 254702 1622 254702 1622 0 la_data_out[36]
rlabel metal2 256954 3920 256954 3920 0 la_data_out[37]
rlabel metal2 261786 2064 261786 2064 0 la_data_out[38]
rlabel metal2 265374 2098 265374 2098 0 la_data_out[39]
rlabel metal2 137678 840 137678 840 0 la_data_out[3]
rlabel metal2 268870 2064 268870 2064 0 la_data_out[40]
rlabel metal2 272458 2098 272458 2098 0 la_data_out[41]
rlabel metal2 276046 534 276046 534 0 la_data_out[42]
rlabel metal2 279542 2098 279542 2098 0 la_data_out[43]
rlabel metal2 283130 806 283130 806 0 la_data_out[44]
rlabel metal2 286626 2098 286626 2098 0 la_data_out[45]
rlabel metal2 290214 840 290214 840 0 la_data_out[46]
rlabel metal2 293710 2064 293710 2064 0 la_data_out[47]
rlabel metal2 295274 2533 295274 2533 0 la_data_out[48]
rlabel metal2 300794 2064 300794 2064 0 la_data_out[49]
rlabel metal2 141503 340 141503 340 0 la_data_out[4]
rlabel metal2 304382 840 304382 840 0 la_data_out[50]
rlabel metal2 307970 840 307970 840 0 la_data_out[51]
rlabel metal2 311466 1588 311466 1588 0 la_data_out[52]
rlabel metal2 315054 806 315054 806 0 la_data_out[53]
rlabel metal2 318550 2064 318550 2064 0 la_data_out[54]
rlabel metal2 322138 772 322138 772 0 la_data_out[55]
rlabel metal2 325634 2064 325634 2064 0 la_data_out[56]
rlabel metal2 329222 772 329222 772 0 la_data_out[57]
rlabel metal2 332718 806 332718 806 0 la_data_out[58]
rlabel metal2 333546 2227 333546 2227 0 la_data_out[59]
rlabel metal2 144762 840 144762 840 0 la_data_out[5]
rlabel metal2 339894 772 339894 772 0 la_data_out[60]
rlabel metal2 343390 806 343390 806 0 la_data_out[61]
rlabel metal2 346978 806 346978 806 0 la_data_out[62]
rlabel metal2 350474 602 350474 602 0 la_data_out[63]
rlabel metal2 354062 534 354062 534 0 la_data_out[64]
rlabel metal2 354430 1887 354430 1887 0 la_data_out[65]
rlabel metal2 361146 772 361146 772 0 la_data_out[66]
rlabel metal2 364642 602 364642 602 0 la_data_out[67]
rlabel metal2 368230 772 368230 772 0 la_data_out[68]
rlabel metal2 371726 602 371726 602 0 la_data_out[69]
rlabel metal2 148350 840 148350 840 0 la_data_out[6]
rlabel metal2 371818 2295 371818 2295 0 la_data_out[70]
rlabel metal2 378902 772 378902 772 0 la_data_out[71]
rlabel metal2 382398 704 382398 704 0 la_data_out[72]
rlabel metal2 385986 738 385986 738 0 la_data_out[73]
rlabel metal2 389482 840 389482 840 0 la_data_out[74]
rlabel metal2 393070 738 393070 738 0 la_data_out[75]
rlabel metal2 392702 1989 392702 1989 0 la_data_out[76]
rlabel metal2 400154 602 400154 602 0 la_data_out[77]
rlabel metal2 403650 840 403650 840 0 la_data_out[78]
rlabel metal2 407238 806 407238 806 0 la_data_out[79]
rlabel metal2 151846 2047 151846 2047 0 la_data_out[7]
rlabel metal2 410826 602 410826 602 0 la_data_out[80]
rlabel metal2 410090 2499 410090 2499 0 la_data_out[81]
rlabel metal2 417910 772 417910 772 0 la_data_out[82]
rlabel metal2 421406 602 421406 602 0 la_data_out[83]
rlabel metal2 424994 738 424994 738 0 la_data_out[84]
rlabel metal2 428490 806 428490 806 0 la_data_out[85]
rlabel metal2 431894 833 431894 833 0 la_data_out[86]
rlabel metal2 431066 1921 431066 1921 0 la_data_out[87]
rlabel metal2 439162 568 439162 568 0 la_data_out[88]
rlabel metal2 442658 636 442658 636 0 la_data_out[89]
rlabel metal2 155671 340 155671 340 0 la_data_out[8]
rlabel metal2 446055 340 446055 340 0 la_data_out[90]
rlabel metal2 449834 806 449834 806 0 la_data_out[91]
rlabel metal2 448454 2533 448454 2533 0 la_data_out[92]
rlabel metal2 456727 340 456727 340 0 la_data_out[93]
rlabel metal2 460269 340 460269 340 0 la_data_out[94]
rlabel metal2 464002 840 464002 840 0 la_data_out[95]
rlabel metal2 467498 806 467498 806 0 la_data_out[96]
rlabel metal2 465842 2465 465842 2465 0 la_data_out[97]
rlabel metal2 469338 1989 469338 1989 0 la_data_out[98]
rlabel metal2 478170 738 478170 738 0 la_data_out[99]
rlabel metal2 159167 340 159167 340 0 la_data_out[9]
rlabel metal2 128202 806 128202 806 0 la_oenb[0]
rlabel metal2 482671 340 482671 340 0 la_oenb[100]
rlabel metal2 486450 840 486450 840 0 la_oenb[101]
rlabel metal2 484334 2363 484334 2363 0 la_oenb[102]
rlabel metal2 487830 2533 487830 2533 0 la_oenb[103]
rlabel metal2 497122 636 497122 636 0 la_oenb[104]
rlabel metal2 500618 704 500618 704 0 la_oenb[105]
rlabel metal2 504015 340 504015 340 0 la_oenb[106]
rlabel metal2 507511 340 507511 340 0 la_oenb[107]
rlabel metal2 505218 2465 505218 2465 0 la_oenb[108]
rlabel metal2 508714 1989 508714 1989 0 la_oenb[109]
rlabel metal2 163905 340 163905 340 0 la_oenb[10]
rlabel metal2 518183 340 518183 340 0 la_oenb[110]
rlabel via1 521686 85 521686 85 0 la_oenb[111]
rlabel metal2 525458 840 525458 840 0 la_oenb[112]
rlabel metal2 522698 2465 522698 2465 0 la_oenb[113]
rlabel metal2 526102 2533 526102 2533 0 la_oenb[114]
rlabel metal2 536130 704 536130 704 0 la_oenb[115]
rlabel metal2 539626 670 539626 670 0 la_oenb[116]
rlabel metal2 543023 340 543023 340 0 la_oenb[117]
rlabel metal2 546710 772 546710 772 0 la_oenb[118]
rlabel metal2 543490 2499 543490 2499 0 la_oenb[119]
rlabel metal2 167401 340 167401 340 0 la_oenb[11]
rlabel metal2 546986 2057 546986 2057 0 la_oenb[120]
rlabel metal2 557382 806 557382 806 0 la_oenb[121]
rlabel metal2 560878 466 560878 466 0 la_oenb[122]
rlabel metal2 564466 534 564466 534 0 la_oenb[123]
rlabel metal2 560970 2533 560970 2533 0 la_oenb[124]
rlabel metal2 564282 1955 564282 1955 0 la_oenb[125]
rlabel metal2 575138 738 575138 738 0 la_oenb[126]
rlabel metal2 578634 840 578634 840 0 la_oenb[127]
rlabel metal2 170798 2047 170798 2047 0 la_oenb[12]
rlabel metal2 174294 2047 174294 2047 0 la_oenb[13]
rlabel metal2 177981 340 177981 340 0 la_oenb[14]
rlabel metal2 181470 2047 181470 2047 0 la_oenb[15]
rlabel metal2 184966 2047 184966 2047 0 la_oenb[16]
rlabel metal2 188554 2047 188554 2047 0 la_oenb[17]
rlabel metal2 192050 2047 192050 2047 0 la_oenb[18]
rlabel metal2 195539 204 195539 204 0 la_oenb[19]
rlabel metal2 132802 2533 132802 2533 0 la_oenb[1]
rlabel metal2 199035 204 199035 204 0 la_oenb[20]
rlabel metal2 202722 2047 202722 2047 0 la_oenb[21]
rlabel metal2 206218 2047 206218 2047 0 la_oenb[22]
rlabel metal2 209776 340 209776 340 0 la_oenb[23]
rlabel metal2 213394 2047 213394 2047 0 la_oenb[24]
rlabel metal2 216890 2064 216890 2064 0 la_oenb[25]
rlabel metal2 220241 340 220241 340 0 la_oenb[26]
rlabel metal2 223737 340 223737 340 0 la_oenb[27]
rlabel metal2 227562 2047 227562 2047 0 la_oenb[28]
rlabel metal2 231058 2064 231058 2064 0 la_oenb[29]
rlabel metal2 135286 2047 135286 2047 0 la_oenb[2]
rlabel metal2 234646 2064 234646 2064 0 la_oenb[30]
rlabel metal2 238142 2064 238142 2064 0 la_oenb[31]
rlabel metal2 241730 2064 241730 2064 0 la_oenb[32]
rlabel metal2 245226 2098 245226 2098 0 la_oenb[33]
rlabel metal2 248715 340 248715 340 0 la_oenb[34]
rlabel metal2 252402 1588 252402 1588 0 la_oenb[35]
rlabel metal2 255898 1588 255898 1588 0 la_oenb[36]
rlabel metal2 259486 2064 259486 2064 0 la_oenb[37]
rlabel metal2 262982 2098 262982 2098 0 la_oenb[38]
rlabel metal2 266570 2064 266570 2064 0 la_oenb[39]
rlabel metal2 138874 806 138874 806 0 la_oenb[3]
rlabel metal2 270066 2098 270066 2098 0 la_oenb[40]
rlabel metal2 273654 2064 273654 2064 0 la_oenb[41]
rlabel metal2 277150 2098 277150 2098 0 la_oenb[42]
rlabel metal2 280738 2064 280738 2064 0 la_oenb[43]
rlabel metal2 284326 840 284326 840 0 la_oenb[44]
rlabel metal2 287822 2132 287822 2132 0 la_oenb[45]
rlabel metal2 291410 806 291410 806 0 la_oenb[46]
rlabel metal2 294906 2098 294906 2098 0 la_oenb[47]
rlabel metal2 296470 2499 296470 2499 0 la_oenb[48]
rlabel metal2 301990 2098 301990 2098 0 la_oenb[49]
rlabel metal2 142462 2047 142462 2047 0 la_oenb[4]
rlabel metal2 305578 806 305578 806 0 la_oenb[50]
rlabel metal2 309074 2098 309074 2098 0 la_oenb[51]
rlabel metal2 312662 840 312662 840 0 la_oenb[52]
rlabel metal2 313858 2533 313858 2533 0 la_oenb[53]
rlabel metal2 319746 840 319746 840 0 la_oenb[54]
rlabel metal2 323334 738 323334 738 0 la_oenb[55]
rlabel metal2 326830 806 326830 806 0 la_oenb[56]
rlabel metal2 330418 738 330418 738 0 la_oenb[57]
rlabel metal2 333914 772 333914 772 0 la_oenb[58]
rlabel metal2 334742 2499 334742 2499 0 la_oenb[59]
rlabel metal2 145958 840 145958 840 0 la_oenb[5]
rlabel metal2 340998 534 340998 534 0 la_oenb[60]
rlabel metal2 344586 772 344586 772 0 la_oenb[61]
rlabel metal2 348082 840 348082 840 0 la_oenb[62]
rlabel metal2 351670 806 351670 806 0 la_oenb[63]
rlabel metal2 352130 2499 352130 2499 0 la_oenb[64]
rlabel metal2 358754 806 358754 806 0 la_oenb[65]
rlabel metal2 362342 806 362342 806 0 la_oenb[66]
rlabel metal2 365838 840 365838 840 0 la_oenb[67]
rlabel metal2 369426 534 369426 534 0 la_oenb[68]
rlabel metal2 372922 534 372922 534 0 la_oenb[69]
rlabel metal2 149783 340 149783 340 0 la_oenb[6]
rlabel metal2 373014 2499 373014 2499 0 la_oenb[70]
rlabel metal2 380006 840 380006 840 0 la_oenb[71]
rlabel metal2 383594 670 383594 670 0 la_oenb[72]
rlabel metal2 386991 340 386991 340 0 la_oenb[73]
rlabel metal2 390678 704 390678 704 0 la_oenb[74]
rlabel metal2 390402 2465 390402 2465 0 la_oenb[75]
rlabel metal2 397762 806 397762 806 0 la_oenb[76]
rlabel metal2 401350 738 401350 738 0 la_oenb[77]
rlabel metal2 404846 772 404846 772 0 la_oenb[78]
rlabel metal2 408434 738 408434 738 0 la_oenb[79]
rlabel metal2 153279 340 153279 340 0 la_oenb[7]
rlabel metal2 411930 772 411930 772 0 la_oenb[80]
rlabel metal2 411194 3281 411194 3281 0 la_oenb[81]
rlabel metal2 419014 670 419014 670 0 la_oenb[82]
rlabel metal2 422602 806 422602 806 0 la_oenb[83]
rlabel via1 425822 221 425822 221 0 la_oenb[84]
rlabel metal2 429686 704 429686 704 0 la_oenb[85]
rlabel metal2 428674 2431 428674 2431 0 la_oenb[86]
rlabel metal2 436770 670 436770 670 0 la_oenb[87]
rlabel metal2 440167 340 440167 340 0 la_oenb[88]
rlabel metal2 443854 704 443854 704 0 la_oenb[89]
rlabel metal2 156630 2047 156630 2047 0 la_oenb[8]
rlabel metal2 447442 840 447442 840 0 la_oenb[90]
rlabel metal2 450938 772 450938 772 0 la_oenb[91]
rlabel metal2 449558 3281 449558 3281 0 la_oenb[92]
rlabel metal2 458114 670 458114 670 0 la_oenb[93]
rlabel metal2 461610 806 461610 806 0 la_oenb[94]
rlabel via1 465014 85 465014 85 0 la_oenb[95]
rlabel metal2 468694 602 468694 602 0 la_oenb[96]
rlabel metal2 466946 2397 466946 2397 0 la_oenb[97]
rlabel metal2 470442 1921 470442 1921 0 la_oenb[98]
rlabel metal2 479366 670 479366 670 0 la_oenb[99]
rlabel metal2 160126 2047 160126 2047 0 la_oenb[9]
rlabel via1 579646 51 579646 51 0 user_clock2
rlabel via1 581210 323 581210 323 0 user_irq[0]
rlabel via1 581854 187 581854 187 0 user_irq[1]
rlabel via1 583602 85 583602 85 0 user_irq[2]
rlabel metal2 598 2064 598 2064 0 wb_clk_i
rlabel metal2 1702 2098 1702 2098 0 wb_rst_i
rlabel metal2 3089 340 3089 340 0 wbs_ack_o
rlabel metal2 7682 2064 7682 2064 0 wbs_adr_i[0]
rlabel metal2 47886 2064 47886 2064 0 wbs_adr_i[10]
rlabel metal2 51382 2064 51382 2064 0 wbs_adr_i[11]
rlabel metal2 57406 3886 57406 3886 0 wbs_adr_i[12]
rlabel metal2 58466 2064 58466 2064 0 wbs_adr_i[13]
rlabel metal2 62054 1588 62054 1588 0 wbs_adr_i[14]
rlabel metal2 65550 1588 65550 1588 0 wbs_adr_i[15]
rlabel metal2 69138 466 69138 466 0 wbs_adr_i[16]
rlabel metal2 74886 3954 74886 3954 0 wbs_adr_i[17]
rlabel metal2 76222 840 76222 840 0 wbs_adr_i[18]
rlabel metal2 79718 2064 79718 2064 0 wbs_adr_i[19]
rlabel metal2 12374 2064 12374 2064 0 wbs_adr_i[1]
rlabel metal2 83306 840 83306 840 0 wbs_adr_i[20]
rlabel metal2 86894 2064 86894 2064 0 wbs_adr_i[21]
rlabel metal2 90390 806 90390 806 0 wbs_adr_i[22]
rlabel metal2 93978 840 93978 840 0 wbs_adr_i[23]
rlabel metal2 97474 840 97474 840 0 wbs_adr_i[24]
rlabel metal2 101062 840 101062 840 0 wbs_adr_i[25]
rlabel metal2 104558 840 104558 840 0 wbs_adr_i[26]
rlabel metal2 108146 806 108146 806 0 wbs_adr_i[27]
rlabel metal2 111642 738 111642 738 0 wbs_adr_i[28]
rlabel metal2 115230 806 115230 806 0 wbs_adr_i[29]
rlabel metal2 17066 1588 17066 1588 0 wbs_adr_i[2]
rlabel metal2 119055 340 119055 340 0 wbs_adr_i[30]
rlabel metal2 122314 806 122314 806 0 wbs_adr_i[31]
rlabel metal2 21850 2064 21850 2064 0 wbs_adr_i[3]
rlabel metal2 26542 2098 26542 2098 0 wbs_adr_i[4]
rlabel metal2 30130 2098 30130 2098 0 wbs_adr_i[5]
rlabel metal2 36614 3920 36614 3920 0 wbs_adr_i[6]
rlabel metal2 37214 2098 37214 2098 0 wbs_adr_i[7]
rlabel metal2 40710 2064 40710 2064 0 wbs_adr_i[8]
rlabel metal2 44298 2064 44298 2064 0 wbs_adr_i[9]
rlabel metal2 4094 1588 4094 1588 0 wbs_cyc_i
rlabel metal2 8786 636 8786 636 0 wbs_dat_i[0]
rlabel metal2 48990 2098 48990 2098 0 wbs_dat_i[10]
rlabel metal2 52578 534 52578 534 0 wbs_dat_i[11]
rlabel metal2 56074 2132 56074 2132 0 wbs_dat_i[12]
rlabel metal2 59662 534 59662 534 0 wbs_dat_i[13]
rlabel metal2 63250 1690 63250 1690 0 wbs_dat_i[14]
rlabel metal2 66937 340 66937 340 0 wbs_dat_i[15]
rlabel metal2 70334 2064 70334 2064 0 wbs_dat_i[16]
rlabel metal2 75990 3886 75990 3886 0 wbs_dat_i[17]
rlabel metal2 77418 806 77418 806 0 wbs_dat_i[18]
rlabel metal2 80914 2098 80914 2098 0 wbs_dat_i[19]
rlabel metal2 16834 3920 16834 3920 0 wbs_dat_i[1]
rlabel metal2 84502 806 84502 806 0 wbs_dat_i[20]
rlabel metal2 87998 2098 87998 2098 0 wbs_dat_i[21]
rlabel metal2 91586 840 91586 840 0 wbs_dat_i[22]
rlabel metal2 95174 2064 95174 2064 0 wbs_dat_i[23]
rlabel metal2 98670 806 98670 806 0 wbs_dat_i[24]
rlabel metal2 102258 806 102258 806 0 wbs_dat_i[25]
rlabel metal2 105754 534 105754 534 0 wbs_dat_i[26]
rlabel metal2 109342 840 109342 840 0 wbs_dat_i[27]
rlabel metal2 114218 2533 114218 2533 0 wbs_dat_i[28]
rlabel metal2 116426 840 116426 840 0 wbs_dat_i[29]
rlabel metal2 18262 1622 18262 1622 0 wbs_dat_i[2]
rlabel metal2 119922 840 119922 840 0 wbs_dat_i[30]
rlabel metal2 123510 738 123510 738 0 wbs_dat_i[31]
rlabel metal2 23046 2098 23046 2098 0 wbs_dat_i[3]
rlabel metal2 27738 2132 27738 2132 0 wbs_dat_i[4]
rlabel metal2 31326 2064 31326 2064 0 wbs_dat_i[5]
rlabel metal2 37718 3886 37718 3886 0 wbs_dat_i[6]
rlabel metal2 38410 2132 38410 2132 0 wbs_dat_i[7]
rlabel metal2 41906 2098 41906 2098 0 wbs_dat_i[8]
rlabel metal2 45494 2098 45494 2098 0 wbs_dat_i[9]
rlabel metal2 9982 1588 9982 1588 0 wbs_dat_o[0]
rlabel metal2 50186 2132 50186 2132 0 wbs_dat_o[10]
rlabel metal2 56302 3920 56302 3920 0 wbs_dat_o[11]
rlabel metal2 57270 2098 57270 2098 0 wbs_dat_o[12]
rlabel metal2 60858 840 60858 840 0 wbs_dat_o[13]
rlabel metal2 64354 2064 64354 2064 0 wbs_dat_o[14]
rlabel metal2 67942 840 67942 840 0 wbs_dat_o[15]
rlabel metal2 71530 2098 71530 2098 0 wbs_dat_o[16]
rlabel metal2 75026 806 75026 806 0 wbs_dat_o[17]
rlabel metal2 78614 2098 78614 2098 0 wbs_dat_o[18]
rlabel metal2 82110 806 82110 806 0 wbs_dat_o[19]
rlabel metal2 18030 3954 18030 3954 0 wbs_dat_o[1]
rlabel metal2 85698 840 85698 840 0 wbs_dat_o[20]
rlabel metal2 89194 840 89194 840 0 wbs_dat_o[21]
rlabel metal2 94530 2499 94530 2499 0 wbs_dat_o[22]
rlabel metal2 96278 2098 96278 2098 0 wbs_dat_o[23]
rlabel metal2 99866 772 99866 772 0 wbs_dat_o[24]
rlabel metal2 103362 2064 103362 2064 0 wbs_dat_o[25]
rlabel metal2 106950 840 106950 840 0 wbs_dat_o[26]
rlabel metal2 110538 806 110538 806 0 wbs_dat_o[27]
rlabel metal2 114034 772 114034 772 0 wbs_dat_o[28]
rlabel metal2 117622 806 117622 806 0 wbs_dat_o[29]
rlabel metal2 19458 2098 19458 2098 0 wbs_dat_o[2]
rlabel metal2 121118 636 121118 636 0 wbs_dat_o[30]
rlabel metal2 124706 806 124706 806 0 wbs_dat_o[31]
rlabel metal2 24242 2132 24242 2132 0 wbs_dat_o[3]
rlabel metal2 28934 1588 28934 1588 0 wbs_dat_o[4]
rlabel metal2 32430 2132 32430 2132 0 wbs_dat_o[5]
rlabel metal2 36018 1588 36018 1588 0 wbs_dat_o[6]
rlabel metal2 39606 1588 39606 1588 0 wbs_dat_o[7]
rlabel metal2 43102 2132 43102 2132 0 wbs_dat_o[8]
rlabel metal2 46690 2132 46690 2132 0 wbs_dat_o[9]
rlabel metal2 11178 2132 11178 2132 0 wbs_sel_i[0]
rlabel metal2 19134 3886 19134 3886 0 wbs_sel_i[1]
rlabel metal2 20654 2132 20654 2132 0 wbs_sel_i[2]
rlabel metal2 25346 2064 25346 2064 0 wbs_sel_i[3]
rlabel metal2 5481 340 5481 340 0 wbs_stb_i
rlabel metal2 6486 1690 6486 1690 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
