* NGSPICE file created from user_proj_example.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
.ends

.subckt sky130_fd_sc_hd__inv_2 A Y VPWR VGND VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__ha_2 VGND VPWR A COUT SUM B VNB VPB
X0 VPWR A a_342_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_766_47# B a_342_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND B a_389_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 COUT a_342_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND A a_766_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_342_199# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 a_468_369# B a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 a_79_21# a_342_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_389_47# a_342_199# a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_389_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 COUT a_342_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR a_342_199# COUT VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND a_79_21# SUM VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR a_79_21# SUM VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND a_342_199# COUT VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 SUM a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR A a_468_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 SUM a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2b_4 B X A_N VGND VPWR VNB VPB
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_33_199# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_33_199# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_47# a_33_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_109_47# a_33_199# a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR X A VNB VPB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
.ends

.subckt sky130_fd_sc_hd__sdlclkp_4 SCE CLK GCLK GATE VGND VPWR VNB VPB
X0 a_257_147# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_109_369# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_465_315# a_287_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_1045_47# GCLK VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_287_413# a_257_147# a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X5 VPWR a_257_147# a_257_243# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 GCLK a_1045_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_257_147# a_257_243# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND a_1045_47# GCLK VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR a_465_315# a_383_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR a_1045_47# GCLK VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_1127_47# a_465_315# a_1045_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_27_47# GATE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 GCLK a_1045_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_287_413# a_257_243# a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_383_413# a_257_147# a_287_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VGND CLK a_1127_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_257_147# CLK VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 GCLK a_1045_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 GCLK a_1045_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_27_47# GATE a_109_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 VPWR CLK a_1045_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1045_47# a_465_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_395_47# a_257_243# a_287_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24 VGND a_1045_47# GCLK VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VGND a_465_315# a_395_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND SCE a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_465_315# a_287_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_1 B Y A VGND VPWR VNB VPB
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_1 Y A VGND VPWR VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22oi_1 B1 A1 B2 A2 Y VPWR VGND VNB VPB
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_381_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_12 A X VGND VPWR VNB VPB
X0 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__xnor2_1 VGND VPWR B Y A VNB VPB
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_4 A Y VPWR VGND VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_16 Y A VGND VPWR VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_1 VGND VPWR A2 A1 B1 Y VNB VPB
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__xor2_1 B X A VPWR VGND VNB VPB
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a222oi_1 VPWR VGND C2 C1 B1 A2 A1 Y B2 VNB VPB
X0 Y B1 a_393_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 VGND A2 a_561_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VGND C2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 Y C2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A1 a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_311_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_311_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_297# B2 a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_109_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_393_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_109_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 a_561_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 Q CLK D VPWR VGND VNB VPB
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X18 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2_0 VPWR VGND X B A VNB VPB
X0 VPWR B a_40_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_40_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VGND B a_123_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_40_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_123_47# A a_40_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_40_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2_0 A X B VGND VPWR VNB VPB
X0 VGND A a_68_355# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_150_355# B a_68_355# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_68_355# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_68_355# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR A a_150_355# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X a_68_355# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a211o_1 VGND VPWR X A2 B1 A1 C1 VNB VPB
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_1 Y B A VGND VPWR VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux2_2 VGND VPWR A1 A0 S X VNB VPB
X0 VPWR S a_591_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_591_369# A0 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_79_21# A1 a_306_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND S a_578_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_306_369# a_257_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 a_79_21# A0 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_288_47# a_257_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_257_199# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_578_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_257_199# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__conb_1 LO HI VPB VNB VGND VPWR
R0 HI VPWR sky130_fd_pr__res_generic_po w=480000u l=45000u
R1 VGND LO sky130_fd_pr__res_generic_po w=480000u l=45000u
.ends

.subckt sky130_fd_sc_hd__fa_2 COUT SUM A B CIN VGND VPWR VNB VPB
X0 a_1171_369# CIN a_1086_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 VGND CIN a_829_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_1086_47# SUM VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 COUT a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_829_369# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 VPWR CIN a_829_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 a_473_371# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X7 a_294_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR A a_473_371# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X9 a_829_369# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_829_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_829_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_473_371# CIN a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X13 a_473_47# CIN a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_473_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VPWR a_1086_47# SUM VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND a_80_21# COUT VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 COUT a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 SUM a_1086_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_80_21# B a_289_371# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X20 a_80_21# B a_294_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND A a_473_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 SUM a_1086_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VPWR a_80_21# COUT VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_289_371# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X25 a_1194_47# CIN a_1086_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_1086_47# a_80_21# a_829_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 VGND A a_1266_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_1266_371# B a_1171_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X29 VPWR A a_1266_371# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X30 a_1266_47# B a_1194_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 a_1086_47# a_80_21# a_829_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_4 Y A VPWR VGND VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_8 A B Y VGND VPWR VNB VPB
X0 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2b_1 B_N Y A VGND VPWR VNB VPB
X0 Y a_74_47# a_265_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR B_N a_74_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_265_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND B_N a_74_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND a_74_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND X A VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or3_1 A X B C VPWR VGND VNB VPB
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21oi_1 A1 B1 Y A2 VPWR VGND VNB VPB
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_6 VPWR VGND X A VNB VPB
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR VPB VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=5.36e+06u area=4.347e+11p
.ends

.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 Y C1 B1 VGND VPWR VNB VPB
X0 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_326_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y C1 a_326_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_2 B1 Y A2 A1 VGND VPWR VNB VPB
X0 VGND A2 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A1 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_29_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A2 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_112_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_112_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_29_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_29_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_8 X A VGND VPWR VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_8 Y A VGND VPWR VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_bd_sram__openram_dff QN D Q clk vdd gnd VSUBS
X0 vdd a_28_102# a_389_712# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1 a_47_611# clk a_197_712# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X2 a_239_76# clk vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3 a_197_712# D vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X4 QN clk a_547_102# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 gnd Q a_739_102# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Q QN gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_389_712# a_239_76# a_47_611# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X8 vdd a_47_611# a_28_102# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X9 a_547_712# a_28_102# vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X10 a_739_712# clk QN vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X11 gnd a_28_102# a_389_102# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_47_611# a_239_76# a_197_102# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_239_76# clk gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_197_102# D gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_389_102# clk a_47_611# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 gnd a_47_611# a_28_102# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_547_102# a_28_102# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_739_102# a_239_76# QN gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 vdd Q a_739_712# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X20 QN a_239_76# a_547_712# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X21 Q QN vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_wmask_dff clk dout_0 din_1 dout_1 din_2
+ dout_2 din_3 dout_3 gnd vdd din_0
Xsky130_fd_bd_sram__openram_dff_0 sky130_fd_bd_sram__openram_dff_0/QN din_3 dout_3
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_1 sky130_fd_bd_sram__openram_dff_1/QN din_2 dout_2
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_2 sky130_fd_bd_sram__openram_dff_2/QN din_1 dout_1
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_3 sky130_fd_bd_sram__openram_dff_3/QN din_0 dout_0
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m3_w1_680_sli_dli_da_p S D G S_uq0
+ VSUBS
X0 D G S VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X1 D G S_uq0 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X2 S_uq0 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m3_w1_680_sli_dli_da_p S D G S_uq0
+ w_n59_84#
X0 D G S w_n59_84# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X1 D G S_uq0 w_n59_84# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X2 S_uq0 G D w_n59_84# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pinv_2 A Z gnd vdd VSUBS
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m3_w1_680_sli_dli_da_p_0 gnd Z A gnd gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m3_w1_680_sli_dli_da_p
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m3_w1_680_sli_dli_da_p_0 vdd Z A vdd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m3_w1_680_sli_dli_da_p
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_360_sli_dli_da_p S D G VSUBS
X0 D G S VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli_da_p S D G w_n59_28#
X0 D G S w_n59_28# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pinv_0 A Z gnd vdd VSUBS
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_360_sli_dli_da_p_0 gnd Z A gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_360_sli_dli_da_p
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli_da_p_0 vdd Z A vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli_da_p
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m2_w0_740_sli_dli_da_p S D G S_uq0
+ VSUBS
X0 D G S VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 S_uq0 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m2_w1_260_sli_dli_da_p S D G S_uq0
+ w_n59_42#
X0 D G S w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X1 S_uq0 G D w_n59_42# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pinv_1 A Z gnd vdd VSUBS
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m2_w0_740_sli_dli_da_p_0 gnd Z A gnd gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m2_w0_740_sli_dli_da_p
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m2_w1_260_sli_dli_da_p_0 vdd Z A vdd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m2_w1_260_sli_dli_da_p
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pinvbuf gnd Z Zb A gnd_uq0 vdd
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_2_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_2_0/A
+ Z gnd vdd VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_pinv_2
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_2_1 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_2_1/A
+ Zb gnd_uq0 vdd VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_pinv_2
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_0_0 A sky130_sram_1kbyte_1rw1r_32x256_8_pinv_2_0/A
+ gnd_uq0 vdd VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_pinv_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_1_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_2_0/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_2_1/A gnd_uq0 vdd VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_pinv_1
.ends

.subckt sky130_fd_bd_sram__openram_dp_nand3_dec A B C Z vdd gnd
X0 Z B vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 vdd C Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 a_198_136# A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 gnd C a_198_208# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 a_198_208# B a_198_136# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec gnd vdd A Z VSUBS
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_360_sli_dli_da_p_0 gnd Z A gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_360_sli_dli_da_p
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli_da_p_0 vdd Z A vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli_da_p
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec vdd_uq0 vdd Z C B A gnd
Xsky130_fd_bd_sram__openram_dp_nand3_dec_0 A B C sky130_fd_bd_sram__openram_dp_nand3_dec_0/Z
+ vdd gnd sky130_fd_bd_sram__openram_dp_nand3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_0 gnd vdd_uq0 sky130_fd_bd_sram__openram_dp_nand3_dec_0/Z
+ Z sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_0/VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_predecode3x8 in_0 in_1 in_2
+ out_0 out_1 out_2 out_3 out_6 out_7 vdd_uq0 vdd vdd_uq2 out_4 out_5 gnd_uq1 gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_0 vdd_uq0 vdd out_7 in_2 in_1 in_0 gnd
+ sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_1 vdd_uq0 vdd out_6 in_2 in_1 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_2/Z
+ gnd sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_2 vdd_uq0 vdd out_5 in_2 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_1/Z
+ in_0 gnd sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_3 vdd_uq0 vdd out_4 in_2 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_1/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_2/Z gnd sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_4 vdd_uq0 vdd out_3 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_0/Z
+ in_1 in_0 gnd sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_5 vdd_uq0 vdd out_2 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_0/Z
+ in_1 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_2/Z gnd sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_6 vdd_uq0 vdd out_1 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_0/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_1/Z in_0 gnd sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_0 gnd_uq1 vdd_uq2 in_2 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_0/Z
+ gnd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_7 vdd_uq0 vdd out_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_0/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_1/Z sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_2/Z
+ gnd sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_1 gnd_uq1 vdd_uq2 in_1 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_1/Z
+ gnd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_2 gnd_uq1 vdd_uq2 in_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_2/Z
+ gnd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec
.ends

.subckt sky130_fd_bd_sram__openram_dp_nand2_dec A B Z vdd gnd VSUBS
X0 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 vdd B Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 a_196_224# B gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 Z A a_196_224# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_and2_dec gnd A B vdd_uq0 gnd_uq0 Z vdd
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_0 gnd_uq0 vdd_uq0 sky130_fd_bd_sram__openram_dp_nand2_dec_0/Z
+ Z VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec
Xsky130_fd_bd_sram__openram_dp_nand2_dec_0 A B sky130_fd_bd_sram__openram_dp_nand2_dec_0/Z
+ vdd gnd VSUBS sky130_fd_bd_sram__openram_dp_nand2_dec
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_predecode2x4 in_0 in_1 out_0
+ out_3 vdd_uq0 vdd_uq1 gnd_uq0 gnd_uq1 out_1 out_2 vdd gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_and2_dec_0 gnd in_0 in_1 vdd_uq0 gnd_uq0 out_3
+ vdd sky130_sram_1kbyte_1rw1r_32x256_8_and2_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and2_dec_2 gnd in_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_0/Z
+ vdd_uq0 gnd_uq0 out_1 vdd sky130_sram_1kbyte_1rw1r_32x256_8_and2_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and2_dec_1 gnd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_1/Z
+ in_1 vdd_uq0 gnd_uq0 out_2 vdd sky130_sram_1kbyte_1rw1r_32x256_8_and2_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and2_dec_3 gnd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_1/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_0/Z vdd_uq0 gnd_uq0 out_0 vdd sky130_sram_1kbyte_1rw1r_32x256_8_and2_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_1 gnd_uq1 vdd_uq1 in_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_1/Z
+ VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_0 gnd_uq1 vdd_uq1 in_1 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_0/Z
+ VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder addr_0 addr_1 addr_2
+ addr_3 addr_4 addr_5 addr_6 predecode_0 predecode_1 predecode_2 predecode_3 predecode_4
+ predecode_5 predecode_6 predecode_7 predecode_8 predecode_9 predecode_10 predecode_11
+ predecode_12 predecode_13 predecode_14 predecode_15 decode_64 decode_65 decode_66
+ decode_67 decode_68 decode_69 decode_70 decode_71 decode_72 decode_73 decode_74
+ decode_75 decode_76 decode_77 decode_78 decode_79 decode_80 decode_81 decode_82
+ decode_83 decode_84 decode_85 decode_86 decode_87 decode_88 decode_89 decode_90
+ decode_91 decode_92 decode_93 decode_94 decode_95 decode_96 decode_97 decode_98
+ decode_99 decode_100 decode_101 decode_102 decode_103 decode_104 decode_105 decode_106
+ decode_107 decode_108 decode_109 decode_110 decode_111 decode_112 decode_113 decode_114
+ decode_115 decode_116 decode_117 decode_118 decode_119 decode_120 decode_121 decode_122
+ decode_123 decode_124 decode_125 decode_126 decode_0 decode_1 decode_2 decode_3
+ decode_4 decode_5 decode_6 decode_7 decode_8 decode_9 decode_10 decode_11 decode_12
+ decode_13 decode_14 decode_15 decode_16 decode_17 decode_18 decode_19 decode_20
+ decode_21 decode_22 decode_23 decode_24 decode_25 decode_26 decode_27 decode_28
+ decode_29 decode_30 decode_31 decode_32 decode_33 decode_34 decode_35 decode_36
+ decode_37 decode_38 decode_39 decode_40 decode_41 decode_42 decode_43 decode_44
+ decode_45 decode_46 decode_47 decode_48 decode_49 decode_50 decode_51 decode_52
+ decode_53 decode_54 decode_55 decode_56 decode_57 decode_58 decode_59 decode_60
+ decode_61 decode_62 decode_63 vdd_uq2 vdd vdd_uq7 vdd_uq8 vdd_uq6 vdd_uq9 vdd_uq22
+ gnd_uq2 gnd_uq1 gnd gnd_uq7 gnd_uq8 gnd_uq6 decode_127 vdd_uq21 vdd_uq12 vdd_uq1
+ gnd_uq11 vdd_uq24 VSUBS
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_108 vdd_uq22 vdd_uq24 decode_118 predecode_15
+ predecode_5 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_119 vdd_uq22 vdd_uq24 decode_107 predecode_14
+ predecode_6 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_predecode3x8_0 addr_4 addr_5 addr_6
+ predecode_8 predecode_9 predecode_10 predecode_11 predecode_14 predecode_15 vdd_uq9
+ vdd_uq21 vdd_uq12 predecode_12 predecode_13 gnd_uq11 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_predecode3x8
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_109 vdd_uq22 vdd_uq24 decode_117 predecode_15
+ predecode_5 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_90 vdd_uq22 vdd_uq24 decode_86 predecode_13
+ predecode_5 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_80 vdd_uq22 vdd_uq24 decode_74 predecode_12
+ predecode_6 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_91 vdd_uq22 vdd_uq24 decode_85 predecode_13
+ predecode_5 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_70 vdd_uq22 vdd_uq24 decode_65 predecode_12
+ predecode_4 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_81 vdd_uq22 vdd_uq24 decode_73 predecode_12
+ predecode_6 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_92 vdd_uq22 vdd_uq24 decode_84 predecode_13
+ predecode_5 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_93 vdd_uq22 vdd_uq24 decode_102 predecode_14
+ predecode_5 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_82 vdd_uq22 vdd_uq24 decode_94 predecode_13
+ predecode_7 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_60 vdd_uq22 vdd_uq24 decode_62 predecode_11
+ predecode_7 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_71 vdd_uq22 vdd_uq24 decode_83 predecode_13
+ predecode_4 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_94 vdd_uq22 vdd_uq24 decode_101 predecode_14
+ predecode_5 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_83 vdd_uq22 vdd_uq24 decode_93 predecode_13
+ predecode_7 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_61 vdd_uq22 vdd_uq24 decode_32 predecode_10
+ predecode_4 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_50 vdd_uq22 vdd_uq24 decode_42 predecode_10
+ predecode_6 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_72 vdd_uq22 vdd_uq24 decode_82 predecode_13
+ predecode_4 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_95 vdd_uq22 vdd_uq24 decode_100 predecode_14
+ predecode_5 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_84 vdd_uq22 vdd_uq24 decode_92 predecode_13
+ predecode_7 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_62 vdd_uq22 vdd_uq24 decode_31 predecode_9
+ predecode_7 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_51 vdd_uq22 vdd_uq24 decode_41 predecode_10
+ predecode_6 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_40 vdd_uq22 vdd_uq24 decode_52 predecode_11
+ predecode_5 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_73 vdd_uq22 vdd_uq24 decode_81 predecode_13
+ predecode_4 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_96 vdd_uq22 vdd_uq24 decode_99 predecode_14
+ predecode_4 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_30 vdd_uq22 vdd_uq24 decode_13 predecode_8
+ predecode_7 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_52 vdd_uq22 vdd_uq24 decode_40 predecode_10
+ predecode_6 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_41 vdd_uq22 vdd_uq24 decode_51 predecode_11
+ predecode_4 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_63 vdd_uq22 vdd_uq24 decode_72 predecode_12
+ predecode_6 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_74 vdd_uq22 vdd_uq24 decode_80 predecode_13
+ predecode_4 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_85 vdd_uq22 vdd_uq24 decode_91 predecode_13
+ predecode_6 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_predecode2x4_0 addr_2 addr_3 predecode_4
+ predecode_7 vdd_uq7 vdd_uq6 gnd_uq7 gnd_uq6 predecode_5 predecode_6 vdd_uq8 gnd_uq8
+ sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_predecode2x4
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_97 vdd_uq22 vdd_uq24 decode_98 predecode_14
+ predecode_4 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_20 vdd_uq22 vdd_uq24 decode_23 predecode_9
+ predecode_5 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_53 vdd_uq22 vdd_uq24 decode_39 predecode_10
+ predecode_5 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_42 vdd_uq22 vdd_uq24 decode_50 predecode_11
+ predecode_4 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_31 vdd_uq22 vdd_uq24 decode_61 predecode_11
+ predecode_7 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_64 vdd_uq22 vdd_uq24 decode_71 predecode_12
+ predecode_5 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_75 vdd_uq22 vdd_uq24 decode_79 predecode_12
+ predecode_7 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_86 vdd_uq22 vdd_uq24 decode_90 predecode_13
+ predecode_6 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_predecode2x4_1 addr_0 addr_1 predecode_0
+ predecode_3 vdd_uq2 vdd_uq1 gnd_uq2 gnd_uq1 predecode_1 predecode_2 vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_predecode2x4
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_98 vdd_uq22 vdd_uq24 decode_97 predecode_14
+ predecode_4 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_10 vdd_uq22 vdd_uq24 decode_2 predecode_8
+ predecode_4 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_21 vdd_uq22 vdd_uq24 decode_22 predecode_9
+ predecode_5 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_54 vdd_uq22 vdd_uq24 decode_38 predecode_10
+ predecode_5 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_43 vdd_uq22 vdd_uq24 decode_49 predecode_11
+ predecode_4 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_32 vdd_uq22 vdd_uq24 decode_60 predecode_11
+ predecode_7 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_65 vdd_uq22 vdd_uq24 decode_70 predecode_12
+ predecode_5 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_76 vdd_uq22 vdd_uq24 decode_78 predecode_12
+ predecode_7 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_87 vdd_uq22 vdd_uq24 decode_89 predecode_13
+ predecode_6 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_99 vdd_uq22 vdd_uq24 decode_127 predecode_15
+ predecode_7 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_11 vdd_uq22 vdd_uq24 decode_1 predecode_8
+ predecode_4 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_0 vdd_uq22 vdd_uq24 decode_12 predecode_8
+ predecode_7 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_22 vdd_uq22 vdd_uq24 decode_21 predecode_9
+ predecode_5 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_55 vdd_uq22 vdd_uq24 decode_37 predecode_10
+ predecode_5 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_44 vdd_uq22 vdd_uq24 decode_48 predecode_11
+ predecode_4 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_33 vdd_uq22 vdd_uq24 decode_59 predecode_11
+ predecode_6 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_66 vdd_uq22 vdd_uq24 decode_69 predecode_12
+ predecode_5 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_77 vdd_uq22 vdd_uq24 decode_77 predecode_12
+ predecode_7 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_88 vdd_uq22 vdd_uq24 decode_88 predecode_13
+ predecode_6 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_12 vdd_uq22 vdd_uq24 decode_0 predecode_8
+ predecode_4 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_23 vdd_uq22 vdd_uq24 decode_20 predecode_9
+ predecode_5 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_56 vdd_uq22 vdd_uq24 decode_36 predecode_10
+ predecode_5 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_45 vdd_uq22 vdd_uq24 decode_47 predecode_10
+ predecode_7 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_34 vdd_uq22 vdd_uq24 decode_58 predecode_11
+ predecode_6 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_67 vdd_uq22 vdd_uq24 decode_68 predecode_12
+ predecode_5 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_78 vdd_uq22 vdd_uq24 decode_76 predecode_12
+ predecode_7 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_89 vdd_uq22 vdd_uq24 decode_87 predecode_13
+ predecode_5 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_1 vdd_uq22 vdd_uq24 decode_11 predecode_8
+ predecode_6 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_24 vdd_uq22 vdd_uq24 decode_19 predecode_9
+ predecode_4 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_13 vdd_uq22 vdd_uq24 decode_30 predecode_9
+ predecode_7 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_57 vdd_uq22 vdd_uq24 decode_35 predecode_10
+ predecode_4 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_46 vdd_uq22 vdd_uq24 decode_46 predecode_10
+ predecode_7 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_35 vdd_uq22 vdd_uq24 decode_57 predecode_11
+ predecode_6 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_68 vdd_uq22 vdd_uq24 decode_67 predecode_12
+ predecode_4 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_79 vdd_uq22 vdd_uq24 decode_75 predecode_12
+ predecode_6 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_2 vdd_uq22 vdd_uq24 decode_10 predecode_8
+ predecode_6 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_25 vdd_uq22 vdd_uq24 decode_18 predecode_9
+ predecode_4 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_14 vdd_uq22 vdd_uq24 decode_29 predecode_9
+ predecode_7 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_58 vdd_uq22 vdd_uq24 decode_34 predecode_10
+ predecode_4 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_47 vdd_uq22 vdd_uq24 decode_45 predecode_10
+ predecode_7 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_36 vdd_uq22 vdd_uq24 decode_56 predecode_11
+ predecode_6 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_69 vdd_uq22 vdd_uq24 decode_66 predecode_12
+ predecode_4 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_3 vdd_uq22 vdd_uq24 decode_9 predecode_8
+ predecode_6 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_26 vdd_uq22 vdd_uq24 decode_17 predecode_9
+ predecode_4 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_59 vdd_uq22 vdd_uq24 decode_33 predecode_10
+ predecode_4 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_15 vdd_uq22 vdd_uq24 decode_28 predecode_9
+ predecode_7 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_48 vdd_uq22 vdd_uq24 decode_44 predecode_10
+ predecode_7 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_37 vdd_uq22 vdd_uq24 decode_55 predecode_11
+ predecode_5 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_4 vdd_uq22 vdd_uq24 decode_8 predecode_8
+ predecode_6 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_5 vdd_uq22 vdd_uq24 decode_7 predecode_8
+ predecode_5 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_27 vdd_uq22 vdd_uq24 decode_16 predecode_9
+ predecode_4 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_16 vdd_uq22 vdd_uq24 decode_27 predecode_9
+ predecode_6 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_49 vdd_uq22 vdd_uq24 decode_43 predecode_10
+ predecode_6 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_38 vdd_uq22 vdd_uq24 decode_54 predecode_11
+ predecode_5 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_28 vdd_uq22 vdd_uq24 decode_15 predecode_8
+ predecode_7 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_17 vdd_uq22 vdd_uq24 decode_26 predecode_9
+ predecode_6 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_39 vdd_uq22 vdd_uq24 decode_53 predecode_11
+ predecode_5 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_120 vdd_uq22 vdd_uq24 decode_106 predecode_14
+ predecode_6 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_6 vdd_uq22 vdd_uq24 decode_6 predecode_8
+ predecode_5 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_110 vdd_uq22 vdd_uq24 decode_116 predecode_15
+ predecode_5 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_121 vdd_uq22 vdd_uq24 decode_105 predecode_14
+ predecode_6 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_7 vdd_uq22 vdd_uq24 decode_5 predecode_8
+ predecode_5 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_29 vdd_uq22 vdd_uq24 decode_14 predecode_8
+ predecode_7 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_18 vdd_uq22 vdd_uq24 decode_25 predecode_9
+ predecode_6 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_19 vdd_uq22 vdd_uq24 decode_24 predecode_9
+ predecode_6 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_100 vdd_uq22 vdd_uq24 decode_126 predecode_15
+ predecode_7 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_111 vdd_uq22 vdd_uq24 decode_115 predecode_15
+ predecode_4 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_122 vdd_uq22 vdd_uq24 decode_104 predecode_14
+ predecode_6 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_8 vdd_uq22 vdd_uq24 decode_4 predecode_8
+ predecode_5 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_101 vdd_uq22 vdd_uq24 decode_125 predecode_15
+ predecode_7 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_112 vdd_uq22 vdd_uq24 decode_114 predecode_15
+ predecode_4 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_123 vdd_uq22 vdd_uq24 decode_103 predecode_14
+ predecode_5 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_9 vdd_uq22 vdd_uq24 decode_3 predecode_8
+ predecode_4 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_102 vdd_uq22 vdd_uq24 decode_124 predecode_15
+ predecode_7 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_113 vdd_uq22 vdd_uq24 decode_113 predecode_15
+ predecode_4 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_124 vdd_uq22 vdd_uq24 decode_96 predecode_14
+ predecode_4 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_103 vdd_uq22 vdd_uq24 decode_123 predecode_15
+ predecode_6 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_114 vdd_uq22 vdd_uq24 decode_112 predecode_15
+ predecode_4 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_125 vdd_uq22 vdd_uq24 decode_95 predecode_13
+ predecode_7 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_104 vdd_uq22 vdd_uq24 decode_122 predecode_15
+ predecode_6 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_115 vdd_uq22 vdd_uq24 decode_111 predecode_14
+ predecode_7 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_126 vdd_uq22 vdd_uq24 decode_64 predecode_12
+ predecode_4 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_105 vdd_uq22 vdd_uq24 decode_121 predecode_15
+ predecode_6 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_116 vdd_uq22 vdd_uq24 decode_110 predecode_14
+ predecode_7 predecode_2 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_127 vdd_uq22 vdd_uq24 decode_63 predecode_11
+ predecode_7 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_106 vdd_uq22 vdd_uq24 decode_120 predecode_15
+ predecode_6 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_117 vdd_uq22 vdd_uq24 decode_109 predecode_14
+ predecode_7 predecode_1 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_107 vdd_uq22 vdd_uq24 decode_119 predecode_15
+ predecode_5 predecode_3 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
Xsky130_sram_1kbyte_1rw1r_32x256_8_and3_dec_118 vdd_uq22 vdd_uq24 decode_108 predecode_14
+ predecode_7 predecode_0 VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_and3_dec
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w7_000_sli_dli_da_p S D G w_n59_616#
X0 D G S w_n59_616# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w7_000_sli_dli_da_p S D G VSUBS
X0 D G S VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_0 A gnd vdd Z VSUBS
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w7_000_sli_dli_da_p_0 vdd Z A vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w7_000_sli_dli_da_p
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w7_000_sli_dli_da_p_0 gnd Z A gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w7_000_sli_dli_da_p
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_and2_dec_0 A B vdd_uq0 vdd gnd Z
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_0_0 sky130_fd_bd_sram__openram_dp_nand2_dec_0/Z
+ gnd vdd_uq0 Z sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_0_0/VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_0
Xsky130_fd_bd_sram__openram_dp_nand2_dec_0 A B sky130_fd_bd_sram__openram_dp_nand2_dec_0/Z
+ vdd gnd sky130_fd_bd_sram__openram_dp_nand2_dec_0/VSUBS sky130_fd_bd_sram__openram_dp_nand2_dec
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver vdd_uq0 gnd_uq0 B A vdd
+ gnd Z
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_0_0 sky130_fd_bd_sram__openram_dp_nand2_dec_0/Z
+ gnd_uq0 vdd_uq0 Z VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_pinv_dec_0
Xsky130_fd_bd_sram__openram_dp_nand2_dec_0 A B sky130_fd_bd_sram__openram_dp_nand2_dec_0/Z
+ vdd gnd VSUBS sky130_fd_bd_sram__openram_dp_nand2_dec
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array en wl_64 wl_65 wl_66
+ wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80
+ wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94
+ wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107
+ wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119
+ wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 in_96 in_80 in_97 in_98
+ in_81 in_99 in_100 in_82 in_101 in_102 in_83 in_103 in_104 in_84 in_105 in_74 in_85
+ in_86 in_75 in_110 in_87 in_65 in_88 in_76 in_90 in_77 in_91 in_92 in_121 in_78
+ in_93 in_79 in_95 in_64 in_6 in_7 in_8 in_9 in_10 in_11 in_12 in_13 in_14 in_15
+ in_16 in_20 in_34 in_35 in_36 in_37 in_38 in_39 in_40 in_41 in_42 in_43 in_44 in_45
+ in_46 in_47 in_50 in_51 in_62 wl_0 wl_32 wl_16 wl_33 wl_8 wl_34 wl_17 wl_35 wl_4
+ wl_36 wl_18 wl_37 wl_9 wl_38 wl_19 wl_39 wl_2 wl_40 wl_20 wl_41 wl_10 wl_42 wl_21
+ wl_43 wl_5 wl_44 wl_22 wl_45 wl_11 wl_46 wl_23 wl_47 wl_1 wl_48 wl_24 wl_49 wl_12
+ wl_50 wl_25 wl_51 wl_6 wl_52 wl_26 wl_53 wl_13 wl_54 wl_27 wl_55 wl_3 wl_56 wl_28
+ wl_57 wl_14 wl_58 wl_29 wl_59 wl_7 wl_60 wl_30 wl_61 wl_15 wl_62 wl_31 wl_63 in_106
+ in_17 in_107 in_18 in_108 in_48 in_19 in_109 in_49 in_27 in_89 in_111 in_28 in_21
+ in_122 in_112 in_29 in_22 in_123 in_113 in_52 in_30 in_23 in_124 in_114 in_53 in_2
+ in_24 in_125 in_54 in_115 in_3 in_25 in_126 in_94 in_55 in_116 in_4 in_26 in_127
+ in_56 in_117 in_0 in_68 in_66 in_57 in_118 in_1 in_69 in_67 in_58 in_119 in_5 in_70
+ in_31 in_59 in_71 in_120 in_63 in_32 in_60 in_72 vdd in_33 vdd_uq0 in_61 gnd_uq0
+ in_73 gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_24 vdd_uq0 gnd_uq0 en in_12 vdd
+ gnd wl_12 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_13 vdd_uq0 gnd_uq0 en in_23 vdd
+ gnd wl_23 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_57 vdd_uq0 gnd_uq0 en in_36 vdd
+ gnd wl_36 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_46 vdd_uq0 gnd_uq0 en in_47 vdd
+ gnd wl_47 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_35 vdd_uq0 gnd_uq0 en in_58 vdd
+ gnd wl_58 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_79 vdd_uq0 gnd_uq0 en in_81 vdd
+ gnd wl_81 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_68 vdd_uq0 gnd_uq0 en in_92 vdd
+ gnd wl_92 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_25 vdd_uq0 gnd_uq0 en in_11 vdd
+ gnd wl_11 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_14 vdd_uq0 gnd_uq0 en in_22 vdd
+ gnd wl_22 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_58 vdd_uq0 gnd_uq0 en in_35 vdd
+ gnd wl_35 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_47 vdd_uq0 gnd_uq0 en in_46 vdd
+ gnd wl_46 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_36 vdd_uq0 gnd_uq0 en in_57 vdd
+ gnd wl_57 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_69 vdd_uq0 gnd_uq0 en in_91 vdd
+ gnd wl_91 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_26 vdd_uq0 gnd_uq0 en in_10 vdd
+ gnd wl_10 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_15 vdd_uq0 gnd_uq0 en in_21 vdd
+ gnd wl_21 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_59 vdd_uq0 gnd_uq0 en in_34 vdd
+ gnd wl_34 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_48 vdd_uq0 gnd_uq0 en in_45 vdd
+ gnd wl_45 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_37 vdd_uq0 gnd_uq0 en in_56 vdd
+ gnd wl_56 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_27 vdd_uq0 gnd_uq0 en in_9 vdd
+ gnd wl_9 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_16 vdd_uq0 gnd_uq0 en in_20 vdd
+ gnd wl_20 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_49 vdd_uq0 gnd_uq0 en in_44 vdd
+ gnd wl_44 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_38 vdd_uq0 gnd_uq0 en in_55 vdd
+ gnd wl_55 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_0 vdd_uq0 gnd_uq0 en in_5 vdd gnd
+ wl_5 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_28 vdd_uq0 gnd_uq0 en in_8 vdd
+ gnd wl_8 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_17 vdd_uq0 gnd_uq0 en in_19 vdd
+ gnd wl_19 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_39 vdd_uq0 gnd_uq0 en in_54 vdd
+ gnd wl_54 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_1 vdd_uq0 gnd_uq0 en in_1 vdd gnd
+ wl_1 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_29 vdd_uq0 gnd_uq0 en in_7 vdd
+ gnd wl_7 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_18 vdd_uq0 gnd_uq0 en in_18 vdd
+ gnd wl_18 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_2 vdd_uq0 gnd_uq0 en in_0 vdd gnd
+ wl_0 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_19 vdd_uq0 gnd_uq0 en in_17 vdd
+ gnd wl_17 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_3 vdd_uq0 gnd_uq0 en in_4 vdd gnd
+ wl_4 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_4 vdd_uq0 gnd_uq0 en in_3 vdd gnd
+ wl_3 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_5 vdd_uq0 gnd_uq0 en in_2 vdd gnd
+ wl_2 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_6 vdd_uq0 gnd_uq0 en in_30 vdd
+ gnd wl_30 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_7 vdd_uq0 gnd_uq0 en in_29 vdd
+ gnd wl_29 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_8 vdd_uq0 gnd_uq0 en in_28 vdd
+ gnd wl_28 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_9 vdd_uq0 gnd_uq0 en in_27 vdd
+ gnd wl_27 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_120 vdd_uq0 gnd_uq0 en in_100 vdd
+ gnd wl_100 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_110 vdd_uq0 gnd_uq0 en in_110 vdd
+ gnd wl_110 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_121 vdd_uq0 gnd_uq0 en in_99 vdd
+ gnd wl_99 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_100 vdd_uq0 gnd_uq0 en in_120 vdd
+ gnd wl_120 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_111 vdd_uq0 gnd_uq0 en in_109 vdd
+ gnd wl_109 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_122 vdd_uq0 gnd_uq0 en in_98 vdd
+ gnd wl_98 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_101 vdd_uq0 gnd_uq0 en in_119 vdd
+ gnd wl_119 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_112 vdd_uq0 gnd_uq0 en in_108 vdd
+ gnd wl_108 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_123 vdd_uq0 gnd_uq0 en in_97 vdd
+ gnd wl_97 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_102 vdd_uq0 gnd_uq0 en in_118 vdd
+ gnd wl_118 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_113 vdd_uq0 gnd_uq0 en in_107 vdd
+ gnd wl_107 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_124 vdd_uq0 gnd_uq0 en in_96 vdd
+ gnd wl_96 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_103 vdd_uq0 gnd_uq0 en in_117 vdd
+ gnd wl_117 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_114 vdd_uq0 gnd_uq0 en in_106 vdd
+ gnd wl_106 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_125 vdd_uq0 gnd_uq0 en in_95 vdd
+ gnd wl_95 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_104 vdd_uq0 gnd_uq0 en in_116 vdd
+ gnd wl_116 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_115 vdd_uq0 gnd_uq0 en in_105 vdd
+ gnd wl_105 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_126 vdd_uq0 gnd_uq0 en in_64 vdd
+ gnd wl_64 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_105 vdd_uq0 gnd_uq0 en in_115 vdd
+ gnd wl_115 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_116 vdd_uq0 gnd_uq0 en in_104 vdd
+ gnd wl_104 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_127 vdd_uq0 gnd_uq0 en in_63 vdd
+ gnd wl_63 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_106 vdd_uq0 gnd_uq0 en in_114 vdd
+ gnd wl_114 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_117 vdd_uq0 gnd_uq0 en in_103 vdd
+ gnd wl_103 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_107 vdd_uq0 gnd_uq0 en in_113 vdd
+ gnd wl_113 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_118 vdd_uq0 gnd_uq0 en in_102 vdd
+ gnd wl_102 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_108 vdd_uq0 gnd_uq0 en in_112 vdd
+ gnd wl_112 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_119 vdd_uq0 gnd_uq0 en in_101 vdd
+ gnd wl_101 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_109 vdd_uq0 gnd_uq0 en in_111 vdd
+ gnd wl_111 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_90 vdd_uq0 gnd_uq0 en in_70 vdd
+ gnd wl_70 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_91 vdd_uq0 gnd_uq0 en in_69 vdd
+ gnd wl_69 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_80 vdd_uq0 gnd_uq0 en in_80 vdd
+ gnd wl_80 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_92 vdd_uq0 gnd_uq0 en in_68 vdd
+ gnd wl_68 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_81 vdd_uq0 gnd_uq0 en in_79 vdd
+ gnd wl_79 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_70 vdd_uq0 gnd_uq0 en in_90 vdd
+ gnd wl_90 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_93 vdd_uq0 gnd_uq0 en in_127 vdd
+ gnd wl_127 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_60 vdd_uq0 gnd_uq0 en in_33 vdd
+ gnd wl_33 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_82 vdd_uq0 gnd_uq0 en in_78 vdd
+ gnd wl_78 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_71 vdd_uq0 gnd_uq0 en in_89 vdd
+ gnd wl_89 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_94 vdd_uq0 gnd_uq0 en in_126 vdd
+ gnd wl_126 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_61 vdd_uq0 gnd_uq0 en in_32 vdd
+ gnd wl_32 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_50 vdd_uq0 gnd_uq0 en in_43 vdd
+ gnd wl_43 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_83 vdd_uq0 gnd_uq0 en in_77 vdd
+ gnd wl_77 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_72 vdd_uq0 gnd_uq0 en in_88 vdd
+ gnd wl_88 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_95 vdd_uq0 gnd_uq0 en in_125 vdd
+ gnd wl_125 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_62 vdd_uq0 gnd_uq0 en in_31 vdd
+ gnd wl_31 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_51 vdd_uq0 gnd_uq0 en in_42 vdd
+ gnd wl_42 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_40 vdd_uq0 gnd_uq0 en in_53 vdd
+ gnd wl_53 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_84 vdd_uq0 gnd_uq0 en in_76 vdd
+ gnd wl_76 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_73 vdd_uq0 gnd_uq0 en in_87 vdd
+ gnd wl_87 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_96 vdd_uq0 gnd_uq0 en in_124 vdd
+ gnd wl_124 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_30 vdd_uq0 gnd_uq0 en in_6 vdd
+ gnd wl_6 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_52 vdd_uq0 gnd_uq0 en in_41 vdd
+ gnd wl_41 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_41 vdd_uq0 gnd_uq0 en in_52 vdd
+ gnd wl_52 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_63 vdd_uq0 gnd_uq0 en in_67 vdd
+ gnd wl_67 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_85 vdd_uq0 gnd_uq0 en in_75 vdd
+ gnd wl_75 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_74 vdd_uq0 gnd_uq0 en in_86 vdd
+ gnd wl_86 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_97 vdd_uq0 gnd_uq0 en in_123 vdd
+ gnd wl_123 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_20 vdd_uq0 gnd_uq0 en in_16 vdd
+ gnd wl_16 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_53 vdd_uq0 gnd_uq0 en in_40 vdd
+ gnd wl_40 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_42 vdd_uq0 gnd_uq0 en in_51 vdd
+ gnd wl_51 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_31 vdd_uq0 gnd_uq0 en in_62 vdd
+ gnd wl_62 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_64 vdd_uq0 gnd_uq0 en in_66 vdd
+ gnd wl_66 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_86 vdd_uq0 gnd_uq0 en in_74 vdd
+ gnd wl_74 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_75 vdd_uq0 gnd_uq0 en in_85 vdd
+ gnd wl_85 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_98 vdd_uq0 gnd_uq0 en in_122 vdd
+ gnd wl_122 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_21 vdd_uq0 gnd_uq0 en in_15 vdd
+ gnd wl_15 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_10 vdd_uq0 gnd_uq0 en in_26 vdd
+ gnd wl_26 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_54 vdd_uq0 gnd_uq0 en in_39 vdd
+ gnd wl_39 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_43 vdd_uq0 gnd_uq0 en in_50 vdd
+ gnd wl_50 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_32 vdd_uq0 gnd_uq0 en in_61 vdd
+ gnd wl_61 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_65 vdd_uq0 gnd_uq0 en in_65 vdd
+ gnd wl_65 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_87 vdd_uq0 gnd_uq0 en in_73 vdd
+ gnd wl_73 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_76 vdd_uq0 gnd_uq0 en in_84 vdd
+ gnd wl_84 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_99 vdd_uq0 gnd_uq0 en in_121 vdd
+ gnd wl_121 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_22 vdd_uq0 gnd_uq0 en in_14 vdd
+ gnd wl_14 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_11 vdd_uq0 gnd_uq0 en in_25 vdd
+ gnd wl_25 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_55 vdd_uq0 gnd_uq0 en in_38 vdd
+ gnd wl_38 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_44 vdd_uq0 gnd_uq0 en in_49 vdd
+ gnd wl_49 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_33 vdd_uq0 gnd_uq0 en in_60 vdd
+ gnd wl_60 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_88 vdd_uq0 gnd_uq0 en in_72 vdd
+ gnd wl_72 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_77 vdd_uq0 gnd_uq0 en in_83 vdd
+ gnd wl_83 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_66 vdd_uq0 gnd_uq0 en in_94 vdd
+ gnd wl_94 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_23 vdd_uq0 gnd_uq0 en in_13 vdd
+ gnd wl_13 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_12 vdd_uq0 gnd_uq0 en in_24 vdd
+ gnd wl_24 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_56 vdd_uq0 gnd_uq0 en in_37 vdd
+ gnd wl_37 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_45 vdd_uq0 gnd_uq0 en in_48 vdd
+ gnd wl_48 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_34 vdd_uq0 gnd_uq0 en in_59 vdd
+ gnd wl_59 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_89 vdd_uq0 gnd_uq0 en in_71 vdd
+ gnd wl_71 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_78 vdd_uq0 gnd_uq0 en in_82 vdd
+ gnd wl_82 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_67 vdd_uq0 gnd_uq0 en in_93 vdd
+ gnd wl_93 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0 wl_en addr_0 addr_1 addr_2
+ addr_3 addr_4 addr_5 addr_6 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73
+ wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87
+ wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101
+ wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113
+ wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125
+ wl_126 wl_127 rbl_wl wl_64 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10
+ wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24
+ wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38
+ wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52
+ wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 vdd_uq2 vdd_uq4
+ vdd_uq76 vdd_uq8 vdd vdd_uq406 vdd_uq407 gnd_uq9 gnd_uq3 gnd_uq20 gnd_uq26 vdd_uq78
+ vdd_uq35 vdd_uq27 vdd_uq51 gnd_uq37 vdd_uq34 vdd_uq3 gnd vdd_uq405
Xsky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0 addr_0 addr_1 addr_2 addr_3
+ addr_4 addr_5 addr_6 sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_1 sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_2
+ sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_3 sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_4
+ sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_5 sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_6
+ sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_7 sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_8
+ sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_9 sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_10
+ sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_11 sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_12
+ sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_13 sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_14
+ sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_15 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_64
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_65 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_66
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_67 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_68
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_69 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_70
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_71 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_72
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_73 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_74
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_75 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_76
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_77 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_78
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_79 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_80
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_81 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_82
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_83 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_84
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_85 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_86
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_87 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_88
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_89 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_90
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_91 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_92
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_93 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_94
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_95 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_96
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_97 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_98
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_99 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_100
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_101 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_102
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_103 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_104
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_105 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_106
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_107 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_108
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_109 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_110
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_111 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_112
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_113 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_114
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_115 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_116
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_117 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_118
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_119 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_120
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_121 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_122
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_123 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_124
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_125 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_126
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_0 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_2 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_3
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_4 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_5
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_6 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_7
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_8 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_9
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_10 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_11
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_12 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_13
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_14 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_15
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_16 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_17
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_18 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_19
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_20 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_21
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_22 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_23
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_24 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_25
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_26 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_27
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_28 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_29
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_30 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_31
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_32 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_33
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_34 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_35
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_36 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_37
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_38 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_39
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_40 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_41
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_42 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_43
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_44 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_45
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_46 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_47
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_48 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_49
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_50 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_51
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_52 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_53
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_54 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_55
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_56 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_57
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_58 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_59
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_60 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_61
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_62 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_63
+ vdd_uq2 vdd_uq3 vdd_uq34 vdd_uq35 vdd_uq27 vdd_uq76 vdd_uq8 sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/gnd_uq2
+ gnd_uq3 gnd_uq9 gnd_uq26 gnd_uq26 gnd_uq20 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_127
+ vdd_uq78 vdd_uq51 vdd_uq4 gnd_uq37 vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder
Xsky130_sram_1kbyte_1rw1r_32x256_8_and2_dec_0_0 wl_en vdd_uq407 vdd_uq405 vdd_uq406
+ gnd rbl_wl sky130_sram_1kbyte_1rw1r_32x256_8_and2_dec_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0 wl_en wl_64 wl_65 wl_66
+ wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80
+ wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94
+ wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107
+ wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119
+ wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_96
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_80 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_97
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_98 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_81
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_99 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_100
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_82 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_101
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_102 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_83
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_103 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_104
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_84 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_105
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_74 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_85
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_86 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_75
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_110 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_87
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_65 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_88
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_76 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_90
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_77 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_91
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_92 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_121
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_78 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_93
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_79 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_95
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_64 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_6
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_7 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_8
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_9 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_10
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_11 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_12
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_13 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_14
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_15 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_16
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_20 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_34
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_35 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_36
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_37 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_38
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_39 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_40
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_41 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_42
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_43 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_44
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_45 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_46
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_47 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_50
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_51 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_62
+ wl_0 wl_32 wl_16 wl_33 wl_8 wl_34 wl_17 wl_35 wl_4 wl_36 wl_18 wl_37 wl_9 wl_38
+ wl_19 wl_39 wl_2 wl_40 wl_20 wl_41 wl_10 wl_42 wl_21 wl_43 wl_5 wl_44 wl_22 wl_45
+ wl_11 wl_46 wl_23 wl_47 wl_1 wl_48 wl_24 wl_49 wl_12 wl_50 wl_25 wl_51 wl_6 wl_52
+ wl_26 wl_53 wl_13 wl_54 wl_27 wl_55 wl_3 wl_56 wl_28 wl_57 wl_14 wl_58 wl_29 wl_59
+ wl_7 wl_60 wl_30 wl_61 wl_15 wl_62 wl_31 wl_63 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_106
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_17 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_107
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_18 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_108
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_48 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_19
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_109 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_49
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_27 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_89
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_111 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_28
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_21 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_122
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_112 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_29
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_22 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_123
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_113 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_52
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_30 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_23
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_124 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_114
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_53 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_2
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_24 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_125
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_54 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_115
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_3 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_25
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_126 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_94
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_55 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_116
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_4 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_26
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_127 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_56
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_117 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_68 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_66
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_57 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_118
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_1 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_69
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_67 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_58
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_119 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_5
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_70 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_31
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_59 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_71
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_120 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_63
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_32 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_60
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_72 vdd_uq406 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_33
+ vdd_uq405 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_61 gnd sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_73
+ gnd sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array
.ends

.subckt sky130_fd_bd_sram__openram_sense_amp bl br dout en vdd vdd_uq0 gnd
X0 a_154_1298# a_96_1689# vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X1 gnd en a_184_1689# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_154_1298# a_96_1689# a_184_1689# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 gnd a_154_1298# dout gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 bl en a_96_1689# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 a_154_1298# en br vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 vdd a_154_1298# a_96_1689# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X7 a_184_1689# a_154_1298# a_96_1689# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 vdd_uq0 a_154_1298# dout vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array vdd data_0 bl_1 bl_2 data_2
+ bl_3 br_3 data_3 br_4 data_4 bl_5 br_5 data_5 br_6 data_6 br_7 data_7 br_8 data_8
+ bl_9 br_9 data_9 data_10 data_11 data_12 data_13 br_14 data_14 bl_15 br_15 data_15
+ bl_16 br_16 data_16 bl_17 br_17 data_17 br_18 data_18 bl_19 br_19 data_20 data_21
+ data_22 data_23 data_24 br_25 data_25 bl_26 br_26 data_26 bl_27 br_27 data_27 bl_28
+ br_28 data_28 bl_29 br_29 data_29 data_30 data_31 vdd_uq0 vdd_uq1 vdd_uq2 vdd_uq3
+ vdd_uq4 vdd_uq5 vdd_uq6 vdd_uq7 vdd_uq8 vdd_uq9 vdd_uq10 vdd_uq11 vdd_uq12 vdd_uq13
+ vdd_uq14 vdd_uq15 vdd_uq16 vdd_uq17 vdd_uq18 vdd_uq19 vdd_uq20 vdd_uq21 vdd_uq22
+ vdd_uq23 vdd_uq24 vdd_uq25 vdd_uq26 vdd_uq27 vdd_uq28 vdd_uq29 vdd_uq30 br_23 br_22
+ br_12 br_2 br_20 br_1 bl_23 bl_22 bl_12 bl_20 br_24 br_13 br_30 br_10 bl_24 bl_30
+ bl_13 bl_7 bl_10 bl_6 data_19 br_21 br_31 br_11 br_0 bl_25 bl_21 bl_18 bl_14 bl_31
+ bl_8 bl_4 bl_11 data_1 bl_0 gnd en vdd_uq62
Xsky130_fd_bd_sram__openram_sense_amp_21 bl_31 br_31 data_31 en vdd_uq62 vdd_uq0 gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_10 bl_11 br_11 data_11 en vdd_uq62 vdd_uq19
+ gnd sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_5 bl_3 br_3 data_3 en vdd_uq62 vdd_uq27 gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_22 bl_30 br_30 data_30 en vdd_uq62 vdd gnd sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_11 bl_10 br_10 data_10 en vdd_uq62 vdd_uq20
+ gnd sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_6 bl_2 br_2 data_2 en vdd_uq62 vdd_uq28 gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_23 bl_29 br_29 data_29 en vdd_uq62 vdd_uq1 gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_7 bl_14 br_14 data_14 en vdd_uq62 vdd_uq16 gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_12 bl_9 br_9 data_9 en vdd_uq62 vdd_uq21 gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_24 bl_28 br_28 data_28 en vdd_uq62 vdd_uq2 gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_8 bl_13 br_13 data_13 en vdd_uq62 vdd_uq17 gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_9 bl_12 br_12 data_12 en vdd_uq62 vdd_uq18 gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_13 bl_8 br_8 data_8 en vdd_uq62 vdd_uq22 gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_25 bl_27 br_27 data_27 en vdd_uq62 vdd_uq3 gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_26 bl_26 br_26 data_26 en vdd_uq62 vdd_uq4 gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_15 bl_19 br_19 data_19 en vdd_uq62 vdd_uq11
+ gnd sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_14 bl_7 br_7 data_7 en vdd_uq62 vdd_uq23 gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_27 bl_25 br_25 data_25 en vdd_uq62 vdd_uq5 gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_16 bl_18 br_18 data_18 en vdd_uq62 vdd_uq12
+ gnd sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_28 bl_24 br_24 data_24 en vdd_uq62 vdd_uq6 gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_17 bl_17 br_17 data_17 en vdd_uq62 vdd_uq13
+ gnd sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_29 bl_23 br_23 data_23 en vdd_uq62 vdd_uq7 gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_18 bl_22 br_22 data_22 en vdd_uq62 vdd_uq8 gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_19 bl_21 br_21 data_21 en vdd_uq62 vdd_uq9 gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_0 bl_1 br_1 data_1 en vdd_uq62 vdd_uq29 gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_1 bl_0 br_0 data_0 en vdd_uq62 vdd_uq30 gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_2 bl_6 br_6 data_6 en vdd_uq62 vdd_uq24 gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_30 bl_16 br_16 data_16 en vdd_uq62 vdd_uq14
+ gnd sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_3 bl_5 br_5 data_5 en vdd_uq62 vdd_uq25 gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_20 bl_20 br_20 data_20 en vdd_uq62 vdd_uq10
+ gnd sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_31 bl_15 br_15 data_15 en vdd_uq62 vdd_uq15
+ gnd sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_4 bl_4 br_4 data_4 en vdd_uq62 vdd_uq26 gnd
+ sky130_fd_bd_sram__openram_sense_amp
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sli_dactive S G a_90_0# w_n26_n26#
+ VSUBS
X0 a_90_0# G S VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sactive_dli D G w_n26_n26#
+ a_0_0# VSUBS
X0 D G a_0_0# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli S D G w_n59_28#
X0 D G S w_n59_28# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pnand2 Z gnd vdd A B w_n36_538# VSUBS
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sli_dactive_0 gnd A sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sactive_dli_0/a_0_0#
+ sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sli_dactive_0/w_n26_n26# VSUBS
+ sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sli_dactive
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sactive_dli_0 Z B sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sli_dactive_0/w_n26_n26#
+ sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sactive_dli_0/a_0_0# VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sactive_dli
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli_0 Z vdd B w_n36_538# sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli_1 vdd Z A w_n36_538# sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pinv A Z gnd vdd
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m2_w0_740_sli_dli_da_p_0 gnd Z A gnd gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m2_w0_740_sli_dli_da_p
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m2_w1_260_sli_dli_da_p_0 vdd Z A vdd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m2_w1_260_sli_dli_da_p
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pdriver Z A vdd gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_0 A Z gnd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pinv
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pand2 Z A B vdd gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_pnand2_0 sky130_sram_1kbyte_1rw1r_32x256_8_pnand2_0/Z
+ gnd vdd A B vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pnand2
Xsky130_sram_1kbyte_1rw1r_32x256_8_pdriver_0 Z sky130_sram_1kbyte_1rw1r_32x256_8_pnand2_0/Z
+ vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pdriver
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_write_mask_and_array wmask_in_0 wmask_in_1
+ wmask_in_2 wmask_in_3 wmask_out_0 wmask_out_1 wmask_out_2 wmask_out_3 vdd en gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_pand2_0 wmask_out_3 wmask_in_3 en vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pand2
Xsky130_sram_1kbyte_1rw1r_32x256_8_pand2_1 wmask_out_2 wmask_in_2 en vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pand2
Xsky130_sram_1kbyte_1rw1r_32x256_8_pand2_2 wmask_out_1 wmask_in_1 en vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pand2
Xsky130_sram_1kbyte_1rw1r_32x256_8_pand2_3 wmask_out_0 wmask_in_0 en vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pand2
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w0_550_sli_dli S D G w_n59_n29#
X0 D G S w_n59_n29# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0 vdd en_bar br bl
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w0_550_sli_dli_0 vdd br en_bar vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w0_550_sli_dli
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w0_550_sli_dli_2 bl br en_bar vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w0_550_sli_dli
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w0_550_sli_dli_1 bl vdd en_bar vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w0_550_sli_dli
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_precharge_array bl_0 br_0 bl_1 br_1 bl_2
+ br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10
+ br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17
+ br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24
+ br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31
+ br_31 br_32 bl_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 br_36 bl_37 br_37 bl_38 br_38
+ bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45
+ bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52
+ bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59
+ bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 vdd bl_36 en_bar
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_39 vdd en_bar br_58 bl_58 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_17 vdd en_bar br_15 bl_15 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_28 vdd en_bar br_4 bl_4 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_18 vdd en_bar br_14 bl_14 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_19 vdd en_bar br_13 bl_13 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_29 vdd en_bar br_3 bl_3 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_0 vdd en_bar br_0 bl_0 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_60 vdd en_bar br_37 bl_37 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_1 vdd en_bar br_31 bl_31 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_50 vdd en_bar br_47 bl_47 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_61 vdd en_bar br_36 bl_36 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_2 vdd en_bar br_30 bl_30 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_3 vdd en_bar br_29 bl_29 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_40 vdd en_bar br_57 bl_57 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_51 vdd en_bar br_46 bl_46 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_62 vdd en_bar br_35 bl_35 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_4 vdd en_bar br_28 bl_28 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_41 vdd en_bar br_56 bl_56 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_52 vdd en_bar br_45 bl_45 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_63 vdd en_bar br_34 bl_34 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_5 vdd en_bar br_27 bl_27 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_30 vdd en_bar br_2 bl_2 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_42 vdd en_bar br_55 bl_55 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_53 vdd en_bar br_44 bl_44 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_64 vdd en_bar br_32 bl_32 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_6 vdd en_bar br_26 bl_26 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_20 vdd en_bar br_12 bl_12 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_31 vdd en_bar br_1 bl_1 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_33 vdd en_bar br_64 bl_64 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_43 vdd en_bar br_54 bl_54 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_44 vdd en_bar br_53 bl_53 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_54 vdd en_bar br_43 bl_43 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_55 vdd en_bar br_42 bl_42 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_32 vdd en_bar br_33 bl_33 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_7 vdd en_bar br_25 bl_25 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_10 vdd en_bar br_22 bl_22 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_11 vdd en_bar br_21 bl_21 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_21 vdd en_bar br_11 bl_11 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_22 vdd en_bar br_10 bl_10 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_34 vdd en_bar br_63 bl_63 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_45 vdd en_bar br_52 bl_52 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_56 vdd en_bar br_41 bl_41 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_8 vdd en_bar br_24 bl_24 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_12 vdd en_bar br_20 bl_20 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_23 vdd en_bar br_9 bl_9 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_35 vdd en_bar br_62 bl_62 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_46 vdd en_bar br_51 bl_51 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_57 vdd en_bar br_40 bl_40 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_9 vdd en_bar br_23 bl_23 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_13 vdd en_bar br_19 bl_19 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_24 vdd en_bar br_8 bl_8 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_36 vdd en_bar br_61 bl_61 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_47 vdd en_bar br_50 bl_50 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_58 vdd en_bar br_39 bl_39 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_14 vdd en_bar br_18 bl_18 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_25 vdd en_bar br_7 bl_7 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_37 vdd en_bar br_60 bl_60 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_48 vdd en_bar br_49 bl_49 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_59 vdd en_bar br_38 bl_38 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_15 vdd en_bar br_17 bl_17 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_26 vdd en_bar br_6 bl_6 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_38 vdd en_bar br_59 bl_59 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_49 vdd en_bar br_48 bl_48 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_16 vdd en_bar br_16 bl_16 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_0_27 vdd en_bar br_5 bl_5 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_0
.ends

.subckt sky130_fd_bd_sram__openram_write_driver din bl br en vdd gnd_uq0 gnd vdd_uq0
X0 a_213_736# en a_129_736# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1 a_271_690# din gnd_uq0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2 vdd a_41_1120# a_121_1585# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3 a_271_690# din vdd_uq0 vdd_uq0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X4 a_129_736# a_271_690# vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X5 a_41_1120# en vdd_uq0 vdd_uq0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X6 br a_121_1585# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_183_1687# a_129_736# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8 gnd_uq0 din a_145_492# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X9 vdd en a_129_736# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X10 gnd a_271_690# a_213_736# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X11 a_183_1687# a_129_736# vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X12 gnd a_183_1687# bl gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 gnd a_41_1120# a_121_1585# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14 vdd_uq0 din a_41_1120# vdd_uq0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X15 a_145_492# en a_41_1120# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_write_driver_array gnd data_0 bl_0 br_0
+ data_1 bl_1 br_1 bl_2 br_2 data_3 bl_3 br_3 data_4 bl_4 br_4 data_5 bl_5 br_5 data_6
+ bl_6 br_6 data_7 bl_7 br_7 data_8 bl_8 br_8 data_9 bl_9 br_9 data_10 bl_10 br_10
+ data_11 bl_11 br_11 data_12 bl_12 br_12 data_13 bl_13 br_13 data_14 bl_14 br_14
+ data_15 bl_15 br_15 data_16 bl_16 br_16 data_17 bl_17 br_17 bl_18 br_18 data_19
+ bl_19 br_19 data_20 bl_20 br_20 data_21 bl_21 br_21 data_22 bl_22 br_22 data_23
+ bl_23 br_23 data_24 bl_24 br_24 data_25 bl_25 br_25 data_26 bl_26 br_26 data_27
+ bl_27 br_27 data_28 bl_28 br_28 data_29 bl_29 br_29 data_30 bl_30 br_30 data_31
+ bl_31 br_31 vdd gnd_uq0 gnd_uq1 gnd_uq2 gnd_uq3 gnd_uq4 gnd_uq5 gnd_uq6 gnd_uq7
+ gnd_uq8 gnd_uq9 gnd_uq10 gnd_uq11 gnd_uq12 gnd_uq13 gnd_uq14 gnd_uq15 gnd_uq16 gnd_uq17
+ gnd_uq18 gnd_uq19 gnd_uq20 gnd_uq21 gnd_uq22 gnd_uq23 gnd_uq24 gnd_uq25 gnd_uq26
+ gnd_uq27 gnd_uq28 gnd_uq29 gnd_uq30 data_18 data_2 vdd_uq62 en_3 en_2 en_1 en_0
+ VSUBS
Xsky130_fd_bd_sram__openram_write_driver_7 data_14 bl_14 br_14 en_1 vdd_uq62 gnd_uq16
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_8 data_13 bl_13 br_13 en_1 vdd_uq62 gnd_uq17
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_9 data_12 bl_12 br_12 en_1 vdd_uq62 gnd_uq18
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_30 data_16 bl_16 br_16 en_2 vdd_uq62 gnd_uq14
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_20 data_20 bl_20 br_20 en_2 vdd_uq62 gnd_uq10
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_31 data_15 bl_15 br_15 en_1 vdd_uq62 gnd_uq15
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_21 data_31 bl_31 br_31 en_3 vdd_uq62 gnd_uq0
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_10 data_11 bl_11 br_11 en_1 vdd_uq62 gnd_uq19
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_22 data_30 bl_30 br_30 en_3 vdd_uq62 gnd
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_11 data_10 bl_10 br_10 en_1 vdd_uq62 gnd_uq20
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_23 data_29 bl_29 br_29 en_3 vdd_uq62 gnd_uq1
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_12 data_9 bl_9 br_9 en_1 vdd_uq62 gnd_uq21
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_24 data_28 bl_28 br_28 en_3 vdd_uq62 gnd_uq2
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_13 data_8 bl_8 br_8 en_1 vdd_uq62 gnd_uq22
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_25 data_27 bl_27 br_27 en_3 vdd_uq62 gnd_uq3
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_26 data_26 bl_26 br_26 en_3 vdd_uq62 gnd_uq4
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_15 data_19 bl_19 br_19 en_2 vdd_uq62 gnd_uq11
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_14 data_7 bl_7 br_7 en_0 vdd_uq62 gnd_uq23
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_27 data_25 bl_25 br_25 en_3 vdd_uq62 gnd_uq5
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_16 data_18 bl_18 br_18 en_2 vdd_uq62 gnd_uq12
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_28 data_24 bl_24 br_24 en_3 vdd_uq62 gnd_uq6
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_17 data_17 bl_17 br_17 en_2 vdd_uq62 gnd_uq13
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_29 data_23 bl_23 br_23 en_2 vdd_uq62 gnd_uq7
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_18 data_22 bl_22 br_22 en_2 vdd_uq62 gnd_uq8
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_19 data_21 bl_21 br_21 en_2 vdd_uq62 gnd_uq9
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_0 data_1 bl_1 br_1 en_0 vdd_uq62 gnd_uq29
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_1 data_0 bl_0 br_0 en_0 vdd_uq62 gnd_uq30
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_2 data_4 bl_4 br_4 en_0 vdd_uq62 gnd_uq26
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_3 data_3 bl_3 br_3 en_0 vdd_uq62 gnd_uq27
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_5 data_6 bl_6 br_6 en_0 vdd_uq62 gnd_uq24
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_4 data_2 bl_2 br_2 en_0 vdd_uq62 gnd_uq28
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_6 data_5 bl_5 br_5 en_0 vdd_uq62 gnd_uq25
+ VSUBS vdd sky130_fd_bd_sram__openram_write_driver
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w2_880_sli_dli S D G VSUBS
X0 D G S VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.88e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_column_mux gnd bl br bl_out br_out sel
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w2_880_sli_dli_0 bl_out bl sel gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w2_880_sli_dli
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w2_880_sli_dli_1 br_out br sel gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w2_880_sli_dli
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_array bl_out_16 bl_out_17 bl_out_18
+ bl_out_19 bl_out_20 bl_out_21 bl_out_22 bl_out_23 bl_out_24 bl_out_25 bl_out_26
+ bl_out_27 bl_out_28 bl_out_29 bl_out_30 bl_out_31 bl_32 br_32 bl_33 br_33 bl_34
+ br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41
+ br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48
+ br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55
+ br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62
+ br_62 bl_63 br_63 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29
+ br_29 bl_30 br_30 bl_31 br_31 bl_out_0 bl_out_1 bl_out_2 bl_out_3 bl_out_4 bl_out_5
+ bl_out_6 bl_out_7 bl_out_8 bl_out_9 bl_out_10 bl_out_11 bl_out_12 bl_out_13 bl_out_14
+ bl_out_15 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6
+ bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14
+ br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21
+ br_21 bl_22 br_22 bl_23 br_23 br_out_0 br_out_8 br_out_4 br_out_9 br_out_2 br_out_10
+ br_out_5 br_out_11 br_out_1 br_out_12 br_out_6 br_out_13 br_out_3 br_out_14 br_out_7
+ br_out_15 br_out_16 br_out_24 br_out_20 br_out_25 br_out_18 br_out_26 br_out_21
+ br_out_27 br_out_17 br_out_28 br_out_22 br_out_29 br_out_19 br_out_30 br_out_23
+ br_out_31 sel_1 sel_0 gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_60 gnd bl_59 br_59 bl_out_29 br_out_29
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_61 gnd bl_58 br_58 bl_out_29 br_out_29
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_50 gnd bl_53 br_53 bl_out_26 br_out_26
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_62 gnd bl_57 br_57 bl_out_28 br_out_28
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_51 gnd bl_52 br_52 bl_out_26 br_out_26
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_40 gnd bl_47 br_47 bl_out_23 br_out_23
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_63 gnd bl_56 br_56 bl_out_28 br_out_28
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_52 gnd bl_51 br_51 bl_out_25 br_out_25
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_41 gnd bl_46 br_46 bl_out_23 br_out_23
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_30 gnd bl_25 br_25 bl_out_12 br_out_12
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_53 gnd bl_50 br_50 bl_out_25 br_out_25
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_42 gnd bl_45 br_45 bl_out_22 br_out_22
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_31 gnd bl_24 br_24 bl_out_12 br_out_12
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_20 gnd bl_19 br_19 bl_out_9 br_out_9
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_54 gnd bl_49 br_49 bl_out_24 br_out_24
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_55 gnd bl_48 br_48 bl_out_24 br_out_24
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_43 gnd bl_44 br_44 bl_out_22 br_out_22
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_44 gnd bl_43 br_43 bl_out_21 br_out_21
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_32 gnd bl_39 br_39 bl_out_19 br_out_19
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_33 gnd bl_38 br_38 bl_out_19 br_out_19
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_21 gnd bl_18 br_18 bl_out_9 br_out_9
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_22 gnd bl_17 br_17 bl_out_8 br_out_8
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_10 gnd bl_13 br_13 bl_out_6 br_out_6
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_11 gnd bl_12 br_12 bl_out_6 br_out_6
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_56 gnd bl_63 br_63 bl_out_31 br_out_31
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_45 gnd bl_42 br_42 bl_out_21 br_out_21
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_34 gnd bl_37 br_37 bl_out_18 br_out_18
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_23 gnd bl_16 br_16 bl_out_8 br_out_8
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_12 gnd bl_11 br_11 bl_out_5 br_out_5
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_57 gnd bl_62 br_62 bl_out_31 br_out_31
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_46 gnd bl_41 br_41 bl_out_20 br_out_20
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_35 gnd bl_36 br_36 bl_out_18 br_out_18
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_24 gnd bl_31 br_31 bl_out_15 br_out_15
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_13 gnd bl_10 br_10 bl_out_5 br_out_5
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_58 gnd bl_61 br_61 bl_out_30 br_out_30
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_47 gnd bl_40 br_40 bl_out_20 br_out_20
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_36 gnd bl_35 br_35 bl_out_17 br_out_17
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_25 gnd bl_30 br_30 bl_out_15 br_out_15
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_14 gnd bl_9 br_9 bl_out_4 br_out_4 sel_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_59 gnd bl_60 br_60 bl_out_30 br_out_30
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_48 gnd bl_55 br_55 bl_out_27 br_out_27
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_37 gnd bl_34 br_34 bl_out_17 br_out_17
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_26 gnd bl_29 br_29 bl_out_14 br_out_14
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_15 gnd bl_8 br_8 bl_out_4 br_out_4 sel_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_49 gnd bl_54 br_54 bl_out_27 br_out_27
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_38 gnd bl_33 br_33 bl_out_16 br_out_16
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_27 gnd bl_28 br_28 bl_out_14 br_out_14
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_16 gnd bl_23 br_23 bl_out_11 br_out_11
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_39 gnd bl_32 br_32 bl_out_16 br_out_16
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_28 gnd bl_27 br_27 bl_out_13 br_out_13
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_17 gnd bl_22 br_22 bl_out_11 br_out_11
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_29 gnd bl_26 br_26 bl_out_13 br_out_13
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_18 gnd bl_21 br_21 bl_out_10 br_out_10
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_19 gnd bl_20 br_20 bl_out_10 br_out_10
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0 gnd bl_7 br_7 bl_out_3 br_out_3 sel_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_1 gnd bl_6 br_6 bl_out_3 br_out_3 sel_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_2 gnd bl_5 br_5 bl_out_2 br_out_2 sel_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_3 gnd bl_4 br_4 bl_out_2 br_out_2 sel_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_4 gnd bl_3 br_3 bl_out_1 br_out_1 sel_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_5 gnd bl_2 br_2 bl_out_1 br_out_1 sel_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_6 gnd bl_1 br_1 bl_out_0 br_out_0 sel_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_7 gnd bl_0 br_0 bl_out_0 br_out_0 sel_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_8 gnd bl_15 br_15 bl_out_7 br_out_7
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_9 gnd bl_14 br_14 bl_out_7 br_out_7
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_port_data sel_0 sel_1 bank_wmask_0 bank_wmask_1
+ bank_wmask_2 bank_wmask_3 wdriver_sel_2 wdriver_sel_3 din_16 din_17 din_19 din_20
+ din_21 din_22 din_23 din_24 din_25 din_26 din_27 din_28 din_29 din_30 din_31 dout_16
+ dout_17 dout_18 dout_19 dout_20 dout_21 dout_22 dout_23 dout_24 dout_25 dout_26
+ dout_27 dout_28 dout_29 dout_30 dout_31 din_12 din_13 dout_0 dout_1 dout_2 dout_3
+ dout_4 dout_5 dout_6 dout_7 dout_8 dout_9 dout_10 dout_11 dout_12 dout_13 dout_14
+ dout_15 din_14 din_15 wdriver_sel_0 wdriver_sel_1 din_0 din_1 din_2 din_3 din_4
+ din_5 din_6 din_7 din_8 din_9 din_10 din_11 rbl_bl rbl_br bl_0 br_0 bl_1 br_1 bl_2
+ br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10
+ br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17
+ br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24
+ br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 br_31
+ bl_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38
+ br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45
+ br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52
+ br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59
+ br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 vdd vdd_uq96 vdd_uq97 vdd_uq98
+ vdd_uq100 vdd_uq101 vdd_uq102 vdd_uq103 vdd_uq104 vdd_uq105 vdd_uq106 vdd_uq107
+ vdd_uq108 vdd_uq109 vdd_uq110 vdd_uq111 vdd_uq112 vdd_uq113 vdd_uq114 vdd_uq115
+ vdd_uq116 vdd_uq117 vdd_uq118 vdd_uq119 vdd_uq120 vdd_uq121 vdd_uq122 vdd_uq123
+ vdd_uq124 vdd_uq125 vdd_uq126 vdd_uq127 vdd_uq159 gnd_uq159 gnd_uq160 gnd_uq161
+ gnd_uq162 gnd_uq163 gnd_uq164 gnd_uq165 gnd_uq166 gnd_uq167 gnd_uq168 gnd_uq169
+ gnd_uq170 gnd_uq171 gnd_uq172 gnd_uq173 gnd_uq174 gnd_uq175 gnd_uq176 gnd_uq177
+ gnd_uq178 gnd_uq179 gnd_uq180 gnd_uq181 gnd_uq182 gnd_uq183 gnd_uq184 gnd_uq185
+ gnd_uq186 gnd_uq187 gnd_uq188 gnd_uq189 gnd_uq190 din_18 vdd_uq193 vdd_uq191 vdd_uq95
+ w_en s_en vdd_uq99 gnd p_en_bar
Xsky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0 vdd_uq97 dout_0 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_2 dout_2 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_3
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_3 dout_3 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_4
+ dout_4 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_5 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_5
+ dout_5 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_6 dout_6 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_7
+ dout_7 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_8 dout_8 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_9
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_9 dout_9 dout_10 dout_11
+ dout_12 dout_13 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_14 dout_14
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_15 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_15
+ dout_15 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_16 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_16
+ dout_16 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_17 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_17
+ dout_17 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_18 dout_18 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_19
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_19 dout_20 dout_21 dout_22
+ dout_23 dout_24 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_25 dout_25
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_26 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_26
+ dout_26 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_27 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_27
+ dout_27 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_28 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_28
+ dout_28 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_29 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_29
+ dout_29 dout_30 dout_31 vdd_uq96 vdd_uq98 vdd_uq99 vdd_uq100 vdd_uq101 vdd_uq102
+ vdd_uq103 vdd_uq104 vdd_uq105 vdd_uq106 vdd_uq107 vdd_uq108 vdd_uq109 vdd_uq110
+ vdd_uq111 vdd_uq112 vdd_uq113 vdd_uq114 vdd_uq115 vdd_uq116 vdd_uq117 vdd_uq118
+ vdd_uq119 vdd_uq120 vdd_uq121 vdd_uq122 vdd_uq123 vdd_uq124 vdd_uq125 vdd_uq126
+ vdd_uq127 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_23 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_22
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_12 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_2
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_20 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_23 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_22
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_12 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_20
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_24 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_13
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_30 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_10
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_24 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_30
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_13 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_7
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_10 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_6
+ dout_19 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_21 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_31
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_11 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_25 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_21
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_18 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_14
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_31 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_8
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_4 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_11
+ dout_1 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_0 gnd s_en vdd_uq95
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array
Xsky130_sram_1kbyte_1rw1r_32x256_8_write_mask_and_array_0 bank_wmask_0 bank_wmask_1
+ bank_wmask_2 bank_wmask_3 wdriver_sel_0 wdriver_sel_1 wdriver_sel_2 wdriver_sel_3
+ vdd_uq193 w_en gnd sky130_sram_1kbyte_1rw1r_32x256_8_write_mask_and_array
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_array_0 rbl_bl rbl_br bl_0 br_0 bl_1
+ br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9
+ br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16
+ br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23
+ br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30
+ br_30 br_31 bl_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 br_35 bl_36 br_36 bl_37 br_37
+ bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44
+ bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51
+ bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58
+ bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 vdd bl_35 p_en_bar sky130_sram_1kbyte_1rw1r_32x256_8_precharge_array
Xsky130_sram_1kbyte_1rw1r_32x256_8_write_driver_array_0 gnd_uq160 din_0 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_0 din_1 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_1 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_2
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_2 din_3 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_3
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_3 din_4 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_4
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_4 din_5 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_5
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_5 din_6 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_6
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_6 din_7 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_7
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_7 din_8 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_8
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_8 din_9 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_9
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_9 din_10 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_10
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_10 din_11 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_11
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_11 din_12 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_12
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_12 din_13 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_13
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_13 din_14 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_14
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_14 din_15 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_15
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_15 din_16 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_16
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_16 din_17 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_17
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_17 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_18
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_18 din_19 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_19
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_19 din_20 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_20
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_20 din_21 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_21
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_21 din_22 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_22
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_22 din_23 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_23
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_23 din_24 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_24
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_24 din_25 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_25
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_25 din_26 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_26
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_26 din_27 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_27
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_27 din_28 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_28
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_28 din_29 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_29
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_29 din_30 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_30
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_30 din_31 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_31
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_31 vdd_uq191 gnd_uq159 gnd_uq161
+ gnd_uq162 gnd_uq163 gnd_uq164 gnd_uq165 gnd_uq166 gnd_uq167 gnd_uq168 gnd_uq169
+ gnd_uq170 gnd_uq171 gnd_uq172 gnd_uq173 gnd_uq174 gnd_uq175 gnd_uq176 gnd_uq177
+ gnd_uq178 gnd_uq179 gnd_uq180 gnd_uq181 gnd_uq182 gnd_uq183 gnd_uq184 gnd_uq185
+ gnd_uq186 gnd_uq187 gnd_uq188 gnd_uq189 gnd_uq190 din_18 din_2 vdd_uq159 wdriver_sel_3
+ wdriver_sel_2 wdriver_sel_1 wdriver_sel_0 gnd sky130_sram_1kbyte_1rw1r_32x256_8_write_driver_array
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_array_0 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_16
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_17 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_18
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_19 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_20
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_21 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_22
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_23 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_24
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_25 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_26
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_27 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_28
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_29 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_30
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_31 bl_32 br_32 bl_33 br_33
+ bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40
+ bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47
+ bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54
+ bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61
+ bl_62 br_62 bl_63 br_63 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28
+ bl_29 br_29 bl_30 br_30 bl_31 br_31 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_1 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_2
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_3 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_4
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_5 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_6
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_7 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_8
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_9 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_10
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_11 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_12
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_13 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_14
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_15 bl_0 br_0 bl_1 br_1 bl_2
+ br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10
+ br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17
+ br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_8 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_4
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_9 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_2
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_10 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_5
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_11 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_12 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_6
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_13 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_3
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_14 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_7
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_15 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_16
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_24 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_20
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_25 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_18
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_26 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_21
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_27 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_17
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_28 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_22
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_29 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_19
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_30 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_23
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_31 sel_1 sel_0 gnd sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_array
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0 gnd bl br bl_out br_out sel
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w2_880_sli_dli_0 bl_out bl sel gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w2_880_sli_dli
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w2_880_sli_dli_1 br_out br sel gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w2_880_sli_dli
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_array_0 bl_out_16 bl_out_17 bl_out_18
+ bl_out_19 bl_out_20 bl_out_21 bl_out_22 bl_out_23 bl_out_24 bl_out_25 bl_out_26
+ bl_out_27 bl_out_28 bl_out_29 bl_out_30 bl_out_31 bl_32 br_32 bl_33 br_33 bl_34
+ br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41
+ br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48
+ br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55
+ br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62
+ br_62 bl_63 br_63 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29
+ br_29 bl_30 br_30 bl_31 br_31 bl_out_0 bl_out_1 bl_out_2 bl_out_3 bl_out_4 bl_out_5
+ bl_out_6 bl_out_7 bl_out_8 bl_out_9 bl_out_10 bl_out_11 bl_out_12 bl_out_13 bl_out_14
+ bl_out_15 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6
+ bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14
+ br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21
+ br_21 bl_22 br_22 bl_23 br_23 br_out_0 br_out_8 br_out_4 br_out_9 br_out_2 br_out_10
+ br_out_5 br_out_11 br_out_1 br_out_12 br_out_6 br_out_13 br_out_3 br_out_14 br_out_7
+ br_out_15 br_out_16 br_out_24 br_out_20 br_out_25 br_out_18 br_out_26 br_out_21
+ br_out_27 br_out_17 br_out_28 br_out_22 br_out_29 br_out_19 br_out_30 br_out_23
+ br_out_31 sel_1 sel_0 gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_0 gnd bl_7 br_7 bl_out_3 br_out_3
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_1 gnd bl_6 br_6 bl_out_3 br_out_3
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_60 gnd bl_59 br_59 bl_out_29 br_out_29
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_2 gnd bl_5 br_5 bl_out_2 br_out_2
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_61 gnd bl_58 br_58 bl_out_29 br_out_29
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_50 gnd bl_53 br_53 bl_out_26 br_out_26
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_3 gnd bl_4 br_4 bl_out_2 br_out_2
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_62 gnd bl_57 br_57 bl_out_28 br_out_28
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_51 gnd bl_52 br_52 bl_out_26 br_out_26
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_40 gnd bl_47 br_47 bl_out_23 br_out_23
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_4 gnd bl_3 br_3 bl_out_1 br_out_1
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_5 gnd bl_2 br_2 bl_out_1 br_out_1
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_63 gnd bl_56 br_56 bl_out_28 br_out_28
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_52 gnd bl_51 br_51 bl_out_25 br_out_25
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_41 gnd bl_46 br_46 bl_out_23 br_out_23
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_30 gnd bl_25 br_25 bl_out_12 br_out_12
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_6 gnd bl_1 br_1 bl_out_0 br_out_0
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_53 gnd bl_50 br_50 bl_out_25 br_out_25
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_42 gnd bl_45 br_45 bl_out_22 br_out_22
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_31 gnd bl_24 br_24 bl_out_12 br_out_12
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_20 gnd bl_19 br_19 bl_out_9 br_out_9
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_7 gnd bl_0 br_0 bl_out_0 br_out_0
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_54 gnd bl_49 br_49 bl_out_24 br_out_24
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_55 gnd bl_48 br_48 bl_out_24 br_out_24
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_43 gnd bl_44 br_44 bl_out_22 br_out_22
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_44 gnd bl_43 br_43 bl_out_21 br_out_21
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_32 gnd bl_39 br_39 bl_out_19 br_out_19
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_33 gnd bl_38 br_38 bl_out_19 br_out_19
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_21 gnd bl_18 br_18 bl_out_9 br_out_9
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_22 gnd bl_17 br_17 bl_out_8 br_out_8
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_8 gnd bl_15 br_15 bl_out_7 br_out_7
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_10 gnd bl_13 br_13 bl_out_6 br_out_6
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_11 gnd bl_12 br_12 bl_out_6 br_out_6
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_56 gnd bl_63 br_63 bl_out_31 br_out_31
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_45 gnd bl_42 br_42 bl_out_21 br_out_21
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_34 gnd bl_37 br_37 bl_out_18 br_out_18
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_23 gnd bl_16 br_16 bl_out_8 br_out_8
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_9 gnd bl_14 br_14 bl_out_7 br_out_7
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_12 gnd bl_11 br_11 bl_out_5 br_out_5
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_57 gnd bl_62 br_62 bl_out_31 br_out_31
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_46 gnd bl_41 br_41 bl_out_20 br_out_20
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_35 gnd bl_36 br_36 bl_out_18 br_out_18
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_24 gnd bl_31 br_31 bl_out_15 br_out_15
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_13 gnd bl_10 br_10 bl_out_5 br_out_5
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_58 gnd bl_61 br_61 bl_out_30 br_out_30
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_47 gnd bl_40 br_40 bl_out_20 br_out_20
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_36 gnd bl_35 br_35 bl_out_17 br_out_17
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_25 gnd bl_30 br_30 bl_out_15 br_out_15
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_14 gnd bl_9 br_9 bl_out_4 br_out_4
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_59 gnd bl_60 br_60 bl_out_30 br_out_30
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_48 gnd bl_55 br_55 bl_out_27 br_out_27
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_37 gnd bl_34 br_34 bl_out_17 br_out_17
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_26 gnd bl_29 br_29 bl_out_14 br_out_14
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_15 gnd bl_8 br_8 bl_out_4 br_out_4
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_49 gnd bl_54 br_54 bl_out_27 br_out_27
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_38 gnd bl_33 br_33 bl_out_16 br_out_16
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_27 gnd bl_28 br_28 bl_out_14 br_out_14
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_16 gnd bl_23 br_23 bl_out_11 br_out_11
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_39 gnd bl_32 br_32 bl_out_16 br_out_16
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_28 gnd bl_27 br_27 bl_out_13 br_out_13
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_17 gnd bl_22 br_22 bl_out_11 br_out_11
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_29 gnd bl_26 br_26 bl_out_13 br_out_13
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_18 gnd bl_21 br_21 bl_out_10 br_out_10
+ sel_1 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0_19 gnd bl_20 br_20 bl_out_10 br_out_10
+ sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_0
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1 vdd en_bar br bl
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w0_550_sli_dli_0 vdd br en_bar vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w0_550_sli_dli
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w0_550_sli_dli_2 bl br en_bar vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w0_550_sli_dli
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w0_550_sli_dli_1 bl vdd en_bar vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w0_550_sli_dli
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_precharge_array_0 bl_0 br_0 bl_1 br_1 bl_2
+ br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10
+ br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17
+ br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24
+ br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31
+ br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38
+ br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45
+ br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52
+ br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59
+ bl_60 br_60 bl_61 br_61 bl_62 bl_63 br_63 bl_64 br_64 bl_56 br_62 vdd en_bar
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_60 vdd en_bar br_37 bl_37 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_50 vdd en_bar br_47 bl_47 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_61 vdd en_bar br_36 bl_36 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_40 vdd en_bar br_57 bl_57 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_51 vdd en_bar br_46 bl_46 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_62 vdd en_bar br_35 bl_35 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_0 vdd en_bar br_0 bl_0 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_41 vdd en_bar br_56 bl_56 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_42 vdd en_bar br_55 bl_55 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_52 vdd en_bar br_45 bl_45 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_53 vdd en_bar br_44 bl_44 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_63 vdd en_bar br_34 bl_34 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_64 vdd en_bar br_32 bl_32 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_1 vdd en_bar br_31 bl_31 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_20 vdd en_bar br_12 bl_12 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_30 vdd en_bar br_2 bl_2 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_31 vdd en_bar br_1 bl_1 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_43 vdd en_bar br_54 bl_54 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_54 vdd en_bar br_43 bl_43 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_32 vdd en_bar br_33 bl_33 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_2 vdd en_bar br_30 bl_30 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_10 vdd en_bar br_22 bl_22 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_21 vdd en_bar br_11 bl_11 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_33 vdd en_bar br_64 bl_64 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_44 vdd en_bar br_53 bl_53 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_55 vdd en_bar br_42 bl_42 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_3 vdd en_bar br_29 bl_29 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_11 vdd en_bar br_21 bl_21 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_22 vdd en_bar br_10 bl_10 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_34 vdd en_bar br_63 bl_63 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_45 vdd en_bar br_52 bl_52 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_56 vdd en_bar br_41 bl_41 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_4 vdd en_bar br_28 bl_28 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_12 vdd en_bar br_20 bl_20 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_23 vdd en_bar br_9 bl_9 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_35 vdd en_bar br_62 bl_62 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_46 vdd en_bar br_51 bl_51 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_57 vdd en_bar br_40 bl_40 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_5 vdd en_bar br_27 bl_27 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_13 vdd en_bar br_19 bl_19 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_24 vdd en_bar br_8 bl_8 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_36 vdd en_bar br_61 bl_61 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_47 vdd en_bar br_50 bl_50 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_58 vdd en_bar br_39 bl_39 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_6 vdd en_bar br_26 bl_26 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_14 vdd en_bar br_18 bl_18 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_25 vdd en_bar br_7 bl_7 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_37 vdd en_bar br_60 bl_60 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_48 vdd en_bar br_49 bl_49 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_59 vdd en_bar br_38 bl_38 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_7 vdd en_bar br_25 bl_25 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_8 vdd en_bar br_24 bl_24 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_15 vdd en_bar br_17 bl_17 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_26 vdd en_bar br_6 bl_6 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_38 vdd en_bar br_59 bl_59 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_49 vdd en_bar br_48 bl_48 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_9 vdd en_bar br_23 bl_23 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_16 vdd en_bar br_16 bl_16 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_27 vdd en_bar br_5 bl_5 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_39 vdd en_bar br_58 bl_58 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_17 vdd en_bar br_15 bl_15 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_18 vdd en_bar br_14 bl_14 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_28 vdd en_bar br_4 bl_4 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_29 vdd en_bar br_3 bl_3 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_1_19 vdd en_bar br_13 bl_13 sky130_sram_1kbyte_1rw1r_32x256_8_precharge_1
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0 sel_0 sel_1 dout_17 dout_18
+ dout_19 dout_20 dout_21 dout_22 dout_23 dout_24 dout_25 dout_26 dout_27 dout_28
+ dout_29 dout_30 dout_31 dout_15 dout_16 dout_0 dout_1 dout_2 dout_3 dout_4 dout_5
+ dout_6 dout_7 dout_8 dout_9 dout_10 dout_11 dout_12 dout_13 dout_14 bl_0 br_0 bl_1
+ br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9
+ br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16
+ br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23
+ br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30
+ br_30 bl_31 br_31 bl_32 rbl_br rbl_bl br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35
+ bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42
+ bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49
+ bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56
+ bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63
+ vdd vdd_uq96 vdd_uq97 vdd_uq98 vdd_uq100 vdd_uq101 vdd_uq102 vdd_uq103 vdd_uq104
+ vdd_uq105 vdd_uq106 vdd_uq107 vdd_uq108 vdd_uq109 vdd_uq110 vdd_uq111 vdd_uq112
+ vdd_uq113 vdd_uq114 vdd_uq115 vdd_uq116 vdd_uq117 vdd_uq118 vdd_uq119 vdd_uq120
+ vdd_uq121 vdd_uq122 vdd_uq123 vdd_uq124 vdd_uq125 vdd_uq126 vdd_uq127 vdd_uq95 s_en
+ p_en_bar vdd_uq99 gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0 vdd_uq97 dout_0 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_2 dout_2 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_3
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_3 dout_3 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_4
+ dout_4 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_5 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_5
+ dout_5 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_6 dout_6 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_7
+ dout_7 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_8 dout_8 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_9
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_9 dout_9 dout_10 dout_11
+ dout_12 dout_13 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_14 dout_14
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_15 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_15
+ dout_15 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_16 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_16
+ dout_16 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_17 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_17
+ dout_17 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_18 dout_18 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_19
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_19 dout_20 dout_21 dout_22
+ dout_23 dout_24 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_25 dout_25
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_26 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_26
+ dout_26 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_27 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_27
+ dout_27 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_28 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_28
+ dout_28 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_29 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_29
+ dout_29 dout_30 dout_31 vdd_uq96 vdd_uq98 vdd_uq99 vdd_uq100 vdd_uq101 vdd_uq102
+ vdd_uq103 vdd_uq104 vdd_uq105 vdd_uq106 vdd_uq107 vdd_uq108 vdd_uq109 vdd_uq110
+ vdd_uq111 vdd_uq112 vdd_uq113 vdd_uq114 vdd_uq115 vdd_uq116 vdd_uq117 vdd_uq118
+ vdd_uq119 vdd_uq120 vdd_uq121 vdd_uq122 vdd_uq123 vdd_uq124 vdd_uq125 vdd_uq126
+ vdd_uq127 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_23 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_22
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_12 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_2
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_20 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_23 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_22
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_12 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_20
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_24 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_13
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_30 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_10
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_24 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_30
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_13 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_7
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_10 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_6
+ dout_19 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_21 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_31
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_11 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_25 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_21
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_18 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_14
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_31 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_8
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_4 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_11
+ dout_1 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_0 gnd s_en vdd_uq95
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array
Xsky130_sram_1kbyte_1rw1r_32x256_8_column_mux_array_0_0 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_16
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_17 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_18
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_19 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_20
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_21 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_22
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_23 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_24
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_25 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_26
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_27 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_28
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_29 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_30
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_31 bl_32 br_32 bl_33 br_33
+ bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40
+ bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47
+ bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54
+ bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61
+ bl_62 br_62 bl_63 br_63 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28
+ bl_29 br_29 bl_30 br_30 bl_31 br_31 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_1 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_2
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_3 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_4
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_5 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_6
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_7 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_8
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_9 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_10
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_11 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_12
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_13 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_14
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/bl_15 bl_0 br_0 bl_1 br_1 bl_2
+ br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10
+ br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17
+ br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_8 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_4
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_9 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_2
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_10 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_5
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_11 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_12 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_6
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_13 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_3
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_14 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_7
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_15 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_16
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_24 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_20
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_25 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_18
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_26 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_21
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_27 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_17
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_28 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_22
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_29 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_19
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_30 sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_23
+ sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0/br_31 sel_1 sel_0 gnd sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_array_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_precharge_array_0_0 bl_0 br_0 bl_1 br_1 bl_2 br_2
+ bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10
+ bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17
+ bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24
+ bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31
+ bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38
+ bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45
+ bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52
+ bl_53 br_53 bl_54 br_54 bl_55 br_55 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60
+ br_60 bl_61 br_61 bl_62 bl_63 br_63 rbl_bl rbl_br bl_56 br_62 vdd p_en_bar sky130_sram_1kbyte_1rw1r_32x256_8_precharge_array_0
.ends

.subckt sky130_fd_bd_sram__openram_dp_cell_replica wl0 wl1 bl0 bl1 br0 br1 a_38_n79#
+ vdd gnd a_400_n79# VSUBS
X0 gnd gnd bl1 gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=80000u
X1 a_38_133# wl0 a_38_133# vdd sky130_fd_pr__special_pfet_pass ad=0p pd=0u as=0p ps=0u w=70000u l=150000u
X2 vdd wl1 br1 gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
X3 gnd gnd a_400_n79# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=80000u
X4 vdd a_38_133# gnd gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
X5 vdd wl1 vdd vdd sky130_fd_pr__special_pfet_pass ad=0p pd=0u as=0p ps=0u w=70000u l=150000u
X6 a_38_133# wl1 bl1 gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
X7 gnd gnd a_38_n79# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=80000u
X8 gnd gnd br1 gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=80000u
X9 a_38_133# vdd gnd gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
X10 br0 wl0 vdd gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
X11 gnd a_38_133# vdd gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
X12 a_38_133# vdd vdd vdd sky130_fd_pr__special_pfet_pass ad=0p pd=0u as=0p ps=0u w=140000u l=150000u
X13 vdd a_38_133# vdd vdd sky130_fd_pr__special_pfet_pass ad=0p pd=0u as=0p ps=0u w=140000u l=150000u
X14 bl0 wl0 a_38_133# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
X15 gnd vdd a_38_133# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
.ends

.subckt sky130_fd_bd_sram__openram_dp_cell_dummy wl0 wl1 vdd bl0 bl1 br0 br1 a_38_n79#
+ w_144_n79# gnd a_400_n79# VSUBS
X0 gnd gnd bl1 gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=80000u
X1 a_400_133# wl1 br1 gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
X2 gnd gnd a_400_n79# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=80000u
X3 a_400_291# gnd gnd gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
X4 a_38_133# wl1 bl1 gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
X5 gnd gnd a_38_n79# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=80000u
X6 gnd gnd br1 gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=80000u
X7 a_38_291# gnd gnd gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
X8 br0 wl0 a_400_291# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
X9 gnd gnd a_400_133# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
X10 bl0 wl0 a_38_291# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
X11 gnd gnd a_38_133# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_replica_column_0 wl_0_97 wl_0_98 wl_0_99
+ wl_0_100 wl_0_101 wl_0_102 wl_0_103 wl_0_104 wl_0_105 wl_0_106 wl_0_107 wl_0_108
+ wl_0_109 wl_0_110 wl_0_111 wl_0_112 wl_0_113 wl_0_114 wl_0_115 wl_0_116 wl_0_117
+ wl_0_118 wl_0_119 wl_0_120 wl_0_121 wl_0_122 wl_0_123 wl_0_124 wl_0_125 wl_0_126
+ wl_0_127 wl_0_128 wl_0_129 wl_1_98 wl_1_99 wl_1_100 wl_1_101 wl_1_102 wl_1_103 wl_1_104
+ wl_1_106 wl_1_107 wl_1_108 wl_1_109 wl_1_110 wl_1_111 wl_1_112 wl_1_113 wl_1_114
+ wl_1_115 wl_1_116 wl_1_117 wl_1_118 wl_1_119 wl_1_120 wl_1_121 wl_1_122 wl_1_123
+ wl_1_124 wl_1_125 wl_1_126 wl_1_127 wl_1_128 wl_1_129 wl_1_65 wl_1_66 wl_1_67 wl_1_68
+ wl_1_69 wl_1_70 wl_1_71 wl_1_72 wl_1_73 wl_1_74 wl_1_75 wl_1_76 wl_1_77 wl_1_78
+ wl_1_79 wl_1_80 wl_1_81 wl_1_82 wl_1_83 wl_1_84 wl_1_85 wl_1_86 wl_1_87 wl_1_88
+ wl_1_89 wl_1_90 wl_1_91 wl_1_92 wl_1_93 wl_1_95 wl_1_96 wl_1_97 wl_0_66 wl_0_67
+ wl_0_68 wl_0_70 wl_0_71 wl_0_72 wl_0_73 wl_0_74 wl_0_75 wl_0_76 wl_0_77 wl_0_78
+ wl_0_79 wl_0_80 wl_0_81 wl_0_82 wl_0_83 wl_0_85 wl_0_86 wl_0_87 wl_0_88 wl_0_89
+ wl_0_90 wl_0_91 wl_0_92 wl_0_93 wl_0_94 wl_0_95 wl_0_96 wl_0_65 wl_0_33 wl_0_34
+ wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43 wl_0_44
+ wl_0_45 wl_0_46 wl_0_47 wl_0_48 wl_0_49 wl_0_50 wl_0_51 wl_0_53 wl_0_54 wl_0_55
+ wl_0_56 wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 wl_1_32
+ wl_1_33 wl_1_34 wl_1_35 wl_1_36 wl_1_37 wl_1_38 wl_1_39 wl_1_40 wl_1_41 wl_1_42
+ wl_1_43 wl_1_44 wl_1_45 wl_1_46 wl_1_47 wl_1_49 wl_1_50 wl_1_51 wl_1_52 wl_1_53
+ wl_1_54 wl_1_55 wl_1_56 wl_1_57 wl_1_58 wl_1_59 wl_1_60 wl_1_61 wl_1_62 wl_1_63
+ wl_1_64 wl_1_0 wl_1_1 wl_1_2 wl_1_3 wl_1_4 wl_1_5 wl_1_6 wl_1_7 wl_1_8 wl_1_9 wl_1_10
+ wl_1_11 wl_1_12 wl_1_13 wl_1_14 wl_1_15 wl_1_16 wl_1_17 wl_1_18 wl_1_19 wl_1_20
+ wl_1_21 wl_1_22 wl_1_23 wl_1_24 wl_1_25 wl_1_26 wl_1_28 wl_1_29 wl_1_30 wl_1_31
+ wl_0_32 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10
+ wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20
+ wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30
+ wl_0_31 vdd wl_1_105 wl_0_84 wl_0_69 wl_0_52 wl_1_27 wl_1_48 wl_1_94 bl_1_0 br_1_0
+ gnd bl_0_0 br_0_0
Xsky130_fd_bd_sram__openram_dp_cell_replica_126 wl_0_66 wl_1_66 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_126/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_115 wl_0_77 wl_1_77 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_115/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_104 wl_0_88 wl_1_88 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_104/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_127 wl_0_65 wl_1_65 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_127/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_116 wl_0_76 wl_1_76 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_116/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_105 wl_0_87 wl_1_87 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_105/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_128 wl_0_64 wl_1_64 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_128/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_117 wl_0_75 wl_1_75 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_117/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_106 wl_0_86 wl_1_86 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_106/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_118 wl_0_74 wl_1_74 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_118/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_107 wl_0_85 wl_1_85 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_107/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_119 wl_0_73 wl_1_73 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_119/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_108 wl_0_84 wl_1_84 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_108/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_109 wl_0_83 wl_1_83 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_109/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_90 wl_0_102 wl_1_102 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_90/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_80 wl_0_112 wl_1_112 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_80/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_91 wl_0_101 wl_1_101 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_91/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_70 wl_0_122 wl_1_122 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_70/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_81 wl_0_111 wl_1_111 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_81/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_92 wl_0_100 wl_1_100 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_92/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_71 wl_0_121 wl_1_121 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_71/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_82 wl_0_110 wl_1_110 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_82/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_93 wl_0_99 wl_1_99 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_93/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_60 wl_0_4 wl_1_4 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_60/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_72 wl_0_120 wl_1_120 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_72/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_83 wl_0_109 wl_1_109 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_83/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_94 wl_0_98 wl_1_98 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_94/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_61 wl_0_3 wl_1_3 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_61/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_50 wl_0_14 wl_1_14 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_50/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_73 wl_0_119 wl_1_119 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_73/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_84 wl_0_108 wl_1_108 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_84/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_95 wl_0_97 wl_1_97 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_95/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_62 wl_0_2 wl_1_2 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_62/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_51 wl_0_13 wl_1_13 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_51/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_40 wl_0_24 wl_1_24 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_40/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_63 wl_0_129 wl_1_129 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_63/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_74 wl_0_118 wl_1_118 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_74/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_85 wl_0_107 wl_1_107 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_85/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_96 wl_0_96 wl_1_96 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_96/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_52 wl_0_12 wl_1_12 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_52/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_41 wl_0_23 wl_1_23 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_41/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_30 wl_0_34 wl_1_34 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_30/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_64 wl_0_128 wl_1_128 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_64/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_75 wl_0_117 wl_1_117 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_75/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_86 wl_0_106 wl_1_106 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_86/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_97 wl_0_95 wl_1_95 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_97/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_dummy_0 wl_0_0 wl_1_0 vdd bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 gnd sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_replica_53 wl_0_11 wl_1_11 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_53/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_42 wl_0_22 wl_1_22 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_42/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_31 wl_0_33 wl_1_33 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_31/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_20 wl_0_44 wl_1_44 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_20/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_65 wl_0_127 wl_1_127 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_65/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_76 wl_0_116 wl_1_116 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_76/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_87 wl_0_105 wl_1_105 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_87/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_54 wl_0_10 wl_1_10 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_54/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_43 wl_0_21 wl_1_21 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_43/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_32 wl_0_32 wl_1_32 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_32/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_21 wl_0_43 wl_1_43 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_21/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_10 wl_0_54 wl_1_54 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_10/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_98 wl_0_94 wl_1_94 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_98/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_66 wl_0_126 wl_1_126 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_66/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_77 wl_0_115 wl_1_115 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_77/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_88 wl_0_104 wl_1_104 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_88/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_55 wl_0_9 wl_1_9 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_55/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_44 wl_0_20 wl_1_20 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_44/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_33 wl_0_31 wl_1_31 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_33/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_22 wl_0_42 wl_1_42 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_22/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_11 wl_0_53 wl_1_53 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_11/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_99 wl_0_93 wl_1_93 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_99/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_67 wl_0_125 wl_1_125 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_67/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_78 wl_0_114 wl_1_114 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_78/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_89 wl_0_103 wl_1_103 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_89/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_56 wl_0_8 wl_1_8 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_56/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_45 wl_0_19 wl_1_19 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_45/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_34 wl_0_30 wl_1_30 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_34/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_23 wl_0_41 wl_1_41 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_23/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_12 wl_0_52 wl_1_52 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_12/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_68 wl_0_124 wl_1_124 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_68/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_79 wl_0_113 wl_1_113 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_79/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_57 wl_0_7 wl_1_7 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_57/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_46 wl_0_18 wl_1_18 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_46/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_35 wl_0_29 wl_1_29 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_35/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_24 wl_0_40 wl_1_40 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_24/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_13 wl_0_51 wl_1_51 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_13/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_69 wl_0_123 wl_1_123 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_69/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_58 wl_0_6 wl_1_6 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_58/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_47 wl_0_17 wl_1_17 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_47/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_36 wl_0_28 wl_1_28 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_36/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_25 wl_0_39 wl_1_39 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_25/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_14 wl_0_50 wl_1_50 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_14/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_0 wl_0_1 wl_1_1 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_0/VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_59 wl_0_5 wl_1_5 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_59/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_48 wl_0_16 wl_1_16 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_48/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_37 wl_0_27 wl_1_27 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_37/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_26 wl_0_38 wl_1_38 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_26/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_15 wl_0_49 wl_1_49 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_15/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_1 wl_0_63 wl_1_63 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_1/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_49 wl_0_15 wl_1_15 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_49/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_38 wl_0_26 wl_1_26 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_38/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_27 wl_0_37 wl_1_37 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_27/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_16 wl_0_48 wl_1_48 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_16/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_39 wl_0_25 wl_1_25 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_39/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_28 wl_0_36 wl_1_36 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_28/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_17 wl_0_47 wl_1_47 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_17/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_2 wl_0_62 wl_1_62 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_2/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_3 wl_0_61 wl_1_61 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_3/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_29 wl_0_35 wl_1_35 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_29/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_18 wl_0_46 wl_1_46 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_18/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_19 wl_0_45 wl_1_45 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_19/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_4 wl_0_60 wl_1_60 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_4/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_5 wl_0_59 wl_1_59 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_5/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_6 wl_0_58 wl_1_58 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_6/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_7 wl_0_57 wl_1_57 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_7/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_120 wl_0_72 wl_1_72 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_120/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_8 wl_0_56 wl_1_56 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_8/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_121 wl_0_71 wl_1_71 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_121/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_110 wl_0_82 wl_1_82 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_110/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_9 wl_0_55 wl_1_55 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_9/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_122 wl_0_70 wl_1_70 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_122/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_111 wl_0_81 wl_1_81 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_111/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_100 wl_0_92 wl_1_92 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_100/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_123 wl_0_69 wl_1_69 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_123/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_112 wl_0_80 wl_1_80 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_112/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_101 wl_0_91 wl_1_91 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_101/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_124 wl_0_68 wl_1_68 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_124/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_113 wl_0_79 wl_1_79 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_113/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_102 wl_0_90 wl_1_90 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_102/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_125 wl_0_67 wl_1_67 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_125/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_114 wl_0_78 wl_1_78 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_114/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_103 wl_0_89 wl_1_89 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica_103/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_replica
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_dummy_array vdd bl_0_0 br_0_0 bl_1_0 br_1_0
+ bl_0_1 br_0_1 bl_1_1 br_1_1 bl_0_2 br_0_2 br_1_2 bl_0_3 br_0_3 bl_1_3 br_1_3 bl_0_4
+ br_0_4 bl_1_4 br_1_4 bl_0_5 br_0_5 bl_1_5 br_1_5 bl_0_6 br_0_6 bl_1_6 br_1_6 bl_0_7
+ br_0_7 bl_1_7 br_1_7 bl_0_8 br_0_8 bl_1_8 br_1_8 bl_0_9 br_0_9 bl_1_9 br_1_9 bl_0_10
+ br_0_10 bl_1_10 br_1_10 bl_0_11 br_0_11 bl_1_11 br_1_11 bl_0_12 br_0_12 bl_1_12
+ br_1_12 bl_0_13 br_0_13 bl_1_13 br_1_13 bl_0_14 br_0_14 bl_1_14 br_1_14 bl_0_15
+ br_0_15 bl_1_15 br_1_15 bl_0_16 br_0_16 bl_1_16 br_1_16 bl_0_17 br_0_17 bl_1_17
+ br_1_17 bl_0_18 br_0_18 bl_1_18 br_1_18 bl_0_19 br_0_19 bl_1_19 br_1_19 bl_0_20
+ br_0_20 br_1_20 bl_0_21 br_0_21 bl_1_21 br_1_21 bl_0_22 br_0_22 br_1_22 bl_0_23
+ br_0_23 bl_1_23 br_1_23 bl_0_24 br_0_24 bl_1_24 br_1_24 bl_0_25 br_0_25 bl_1_25
+ br_1_25 bl_0_26 br_0_26 bl_1_26 br_1_26 bl_0_27 br_0_27 bl_1_27 br_1_27 bl_0_28
+ br_0_28 bl_1_28 br_1_28 bl_0_29 br_0_29 bl_1_29 br_1_29 bl_0_30 br_0_30 bl_1_30
+ br_1_30 bl_0_31 br_0_31 bl_1_31 br_1_31 bl_0_32 br_0_32 bl_1_32 br_1_32 bl_0_33
+ br_0_33 br_1_33 bl_0_34 br_0_34 bl_1_34 br_1_34 br_0_35 bl_1_35 br_1_35 bl_0_36
+ br_0_36 bl_1_36 br_1_36 bl_0_37 br_0_37 bl_1_37 br_1_37 bl_0_38 br_0_38 bl_1_38
+ br_1_38 bl_0_39 br_0_39 bl_1_39 br_1_39 bl_0_40 br_0_40 br_1_40 bl_0_41 br_0_41
+ bl_1_41 br_1_41 bl_0_42 br_0_42 bl_1_42 br_1_42 bl_0_43 br_0_43 bl_1_43 br_1_43
+ bl_0_44 br_0_44 bl_1_44 br_1_44 bl_0_45 br_0_45 bl_1_45 br_1_45 bl_0_46 br_0_46
+ bl_1_46 br_1_46 bl_0_47 br_0_47 bl_1_47 br_1_47 bl_0_48 br_0_48 bl_1_48 br_1_48
+ bl_0_49 br_0_49 bl_1_49 br_1_49 bl_0_50 br_0_50 bl_1_50 br_1_50 bl_0_51 br_0_51
+ br_1_51 bl_0_52 br_0_52 bl_1_52 br_1_52 bl_0_53 br_0_53 br_1_53 bl_0_54 br_0_54
+ bl_1_54 br_1_54 bl_0_55 br_0_55 bl_1_55 br_1_55 bl_0_56 br_0_56 bl_1_56 br_1_56
+ bl_0_57 br_0_57 bl_1_57 br_1_57 bl_0_58 bl_1_58 br_1_58 bl_0_59 br_0_59 bl_1_59
+ br_1_59 bl_0_60 br_0_60 bl_1_60 br_1_60 bl_0_61 br_0_61 bl_1_61 br_1_61 bl_0_62
+ br_0_62 bl_1_62 br_1_62 bl_0_63 br_0_63 bl_1_63 br_1_63 vdd_uq0 vdd_uq1 vdd_uq2
+ vdd_uq3 vdd_uq4 vdd_uq5 vdd_uq6 vdd_uq7 vdd_uq8 vdd_uq9 vdd_uq10 vdd_uq11 vdd_uq12
+ vdd_uq13 vdd_uq14 vdd_uq15 vdd_uq16 vdd_uq17 vdd_uq18 vdd_uq19 vdd_uq20 vdd_uq21
+ vdd_uq22 vdd_uq23 vdd_uq24 vdd_uq25 vdd_uq26 vdd_uq27 vdd_uq28 vdd_uq29 vdd_uq30
+ vdd_uq31 vdd_uq32 vdd_uq33 vdd_uq34 vdd_uq35 vdd_uq36 vdd_uq37 vdd_uq38 vdd_uq39
+ vdd_uq40 vdd_uq41 vdd_uq42 vdd_uq43 vdd_uq44 vdd_uq45 vdd_uq46 vdd_uq47 vdd_uq48
+ vdd_uq49 vdd_uq50 vdd_uq51 vdd_uq52 vdd_uq53 vdd_uq54 vdd_uq55 vdd_uq56 vdd_uq57
+ vdd_uq58 vdd_uq59 vdd_uq60 vdd_uq61 vdd_uq62 sky130_fd_bd_sram__openram_dp_cell_dummy_0/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_44/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_36/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_54/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_15/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_5/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_32/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_25/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_61/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_10/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_17/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_0/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_35/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_20/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_45/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_13/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_46/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_30/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_55/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_16/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_6/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_42/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_40/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_26/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_50/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_11/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_27/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_1/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_36/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_9/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_21/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_60/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_23/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_46/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_56/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_31/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_5/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_56/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_17/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_7/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_52/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_41/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_27/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_1/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_12/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_51/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_37/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_2/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_37/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_61/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_22/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_47/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_33/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_32/w_144_n79# bl_1_51 sky130_fd_bd_sram__openram_dp_cell_dummy_57/a_400_n79#
+ bl_1_33 sky130_fd_bd_sram__openram_dp_cell_dummy_18/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_8/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_62/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_18/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_42/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_28/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_52/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_14/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_13/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_47/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_3/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_38/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_23/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_62/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_10/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_43/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_48/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_33/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_19/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_58/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_9/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_28/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_43/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_29/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_24/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_14/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_53/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_57/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_4/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_39/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_6/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_63/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_24/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_20/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_53/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_49/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_34/w_144_n79# bl_0_35 sky130_fd_bd_sram__openram_dp_cell_dummy_2/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_59/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_38/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_44/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_54/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_34/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_15/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_5/w_144_n79# bl_1_20 bl_1_2 sky130_fd_bd_sram__openram_dp_cell_dummy_25/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_30/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_63/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_19/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_35/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_10/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_0/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_15/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_48/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_45/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_20/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_11/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_55/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_44/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_16/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_6/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_30/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_26/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_40/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_40/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_29/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_36/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_50/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_11/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_1/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_25/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_58/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_46/w_144_n79# bl_1_53 sky130_fd_bd_sram__openram_dp_cell_dummy_60/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_21/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_7/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_21/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_54/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_56/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_17/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_7/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_31/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_3/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_27/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_50/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_41/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_39/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_37/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_51/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_12/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_2/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_35/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_47/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_61/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_22/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_31/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_57/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_18/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_8/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_32/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_28/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_60/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_42/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_16/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_49/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_38/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_52/a_400_n79# br_0_58 sky130_fd_bd_sram__openram_dp_cell_dummy_13/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_3/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_12/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_45/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_48/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_62/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_23/a_400_n79#
+ wl_1_0 sky130_fd_bd_sram__openram_dp_cell_dummy_41/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_19/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_58/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_9/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_33/a_400_n79# wl_0_0 sky130_fd_bd_sram__openram_dp_cell_dummy_29/w_144_n79#
+ bl_1_40 sky130_fd_bd_sram__openram_dp_cell_dummy_43/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_26/a_38_n79#
+ bl_1_22 sky130_fd_bd_sram__openram_dp_cell_dummy_59/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_39/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_53/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_14/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_8/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_4/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_22/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_55/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_49/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_63/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_24/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_4/a_38_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_51/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_59/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_34/a_400_n79#
Xsky130_fd_bd_sram__openram_dp_cell_dummy_60 wl_0_0 wl_1_0 vdd_uq59 bl_0_3 bl_1_3
+ br_0_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell_dummy_60/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_60/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_60/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_60/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_50 wl_0_0 wl_1_0 vdd_uq49 bl_0_13 bl_1_13
+ br_0_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell_dummy_50/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_50/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_50/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_50/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_61 wl_0_0 wl_1_0 vdd_uq60 bl_0_2 bl_1_2
+ br_0_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell_dummy_61/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_61/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_61/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_61/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_40 wl_0_0 wl_1_0 vdd_uq39 bl_0_23 bl_1_23
+ br_0_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell_dummy_40/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_40/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_40/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_40/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_51 wl_0_0 wl_1_0 vdd_uq50 bl_0_12 bl_1_12
+ br_0_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell_dummy_51/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_51/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_51/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_51/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_62 wl_0_0 wl_1_0 vdd_uq61 bl_0_1 bl_1_1
+ br_0_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell_dummy_62/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_62/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_62/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_62/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_30 wl_0_0 wl_1_0 vdd_uq29 bl_0_33 bl_1_33
+ br_0_33 br_1_33 sky130_fd_bd_sram__openram_dp_cell_dummy_30/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_30/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_30/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_30/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_41 wl_0_0 wl_1_0 vdd_uq40 bl_0_22 bl_1_22
+ br_0_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell_dummy_41/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_41/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_41/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_41/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_52 wl_0_0 wl_1_0 vdd_uq51 bl_0_11 bl_1_11
+ br_0_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell_dummy_52/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_52/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_52/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_52/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_63 wl_0_0 wl_1_0 vdd_uq62 bl_0_0 bl_1_0
+ br_0_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_dummy_63/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_63/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_63/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_63/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_10 wl_0_0 wl_1_0 vdd_uq9 bl_0_53 bl_1_53
+ br_0_53 br_1_53 sky130_fd_bd_sram__openram_dp_cell_dummy_10/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_10/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_10/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_10/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_20 wl_0_0 wl_1_0 vdd_uq19 bl_0_43 bl_1_43
+ br_0_43 br_1_43 sky130_fd_bd_sram__openram_dp_cell_dummy_20/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_20/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_20/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_20/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_21 wl_0_0 wl_1_0 vdd_uq20 bl_0_42 bl_1_42
+ br_0_42 br_1_42 sky130_fd_bd_sram__openram_dp_cell_dummy_21/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_21/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_21/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_21/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_31 wl_0_0 wl_1_0 vdd_uq30 bl_0_32 bl_1_32
+ br_0_32 br_1_32 sky130_fd_bd_sram__openram_dp_cell_dummy_31/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_31/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_31/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_31/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_32 wl_0_0 wl_1_0 vdd_uq31 bl_0_31 bl_1_31
+ br_0_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell_dummy_32/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_32/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_32/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_32/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_42 wl_0_0 wl_1_0 vdd_uq41 bl_0_21 bl_1_21
+ br_0_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell_dummy_42/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_42/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_42/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_42/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_43 wl_0_0 wl_1_0 vdd_uq42 bl_0_20 bl_1_20
+ br_0_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell_dummy_43/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_43/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_43/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_43/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_53 wl_0_0 wl_1_0 vdd_uq52 bl_0_10 bl_1_10
+ br_0_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell_dummy_53/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_53/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_53/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_53/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_54 wl_0_0 wl_1_0 vdd_uq53 bl_0_9 bl_1_9
+ br_0_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell_dummy_54/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_54/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_54/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_54/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_11 wl_0_0 wl_1_0 vdd_uq10 bl_0_52 bl_1_52
+ br_0_52 br_1_52 sky130_fd_bd_sram__openram_dp_cell_dummy_11/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_11/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_11/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_11/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_22 wl_0_0 wl_1_0 vdd_uq21 bl_0_41 bl_1_41
+ br_0_41 br_1_41 sky130_fd_bd_sram__openram_dp_cell_dummy_22/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_22/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_22/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_22/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_33 wl_0_0 wl_1_0 vdd_uq32 bl_0_30 bl_1_30
+ br_0_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell_dummy_33/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_33/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_33/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_33/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_44 wl_0_0 wl_1_0 vdd_uq43 bl_0_19 bl_1_19
+ br_0_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell_dummy_44/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_44/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_44/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_44/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_55 wl_0_0 wl_1_0 vdd_uq54 bl_0_8 bl_1_8
+ br_0_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell_dummy_55/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_55/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_55/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_55/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_0 wl_0_0 wl_1_0 vdd_uq0 bl_0_63 bl_1_63
+ br_0_63 br_1_63 sky130_fd_bd_sram__openram_dp_cell_dummy_0/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_0/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_0/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_0/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_12 wl_0_0 wl_1_0 vdd_uq11 bl_0_51 bl_1_51
+ br_0_51 br_1_51 sky130_fd_bd_sram__openram_dp_cell_dummy_12/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_12/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_12/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_12/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_23 wl_0_0 wl_1_0 vdd_uq22 bl_0_40 bl_1_40
+ br_0_40 br_1_40 sky130_fd_bd_sram__openram_dp_cell_dummy_23/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_23/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_23/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_23/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_34 wl_0_0 wl_1_0 vdd_uq33 bl_0_29 bl_1_29
+ br_0_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell_dummy_34/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_34/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_34/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_34/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_45 wl_0_0 wl_1_0 vdd_uq44 bl_0_18 bl_1_18
+ br_0_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell_dummy_45/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_45/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_45/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_45/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_56 wl_0_0 wl_1_0 vdd_uq55 bl_0_7 bl_1_7
+ br_0_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell_dummy_56/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_56/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_56/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_56/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_1 wl_0_0 wl_1_0 vdd bl_0_62 bl_1_62 br_0_62
+ br_1_62 sky130_fd_bd_sram__openram_dp_cell_dummy_1/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_1/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_1/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_1/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_13 wl_0_0 wl_1_0 vdd_uq12 bl_0_50 bl_1_50
+ br_0_50 br_1_50 sky130_fd_bd_sram__openram_dp_cell_dummy_13/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_13/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_13/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_13/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_24 wl_0_0 wl_1_0 vdd_uq23 bl_0_39 bl_1_39
+ br_0_39 br_1_39 sky130_fd_bd_sram__openram_dp_cell_dummy_24/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_24/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_24/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_24/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_35 wl_0_0 wl_1_0 vdd_uq34 bl_0_28 bl_1_28
+ br_0_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell_dummy_35/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_35/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_35/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_35/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_46 wl_0_0 wl_1_0 vdd_uq45 bl_0_17 bl_1_17
+ br_0_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell_dummy_46/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_46/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_46/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_46/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_57 wl_0_0 wl_1_0 vdd_uq56 bl_0_6 bl_1_6
+ br_0_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell_dummy_57/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_57/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_57/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_57/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_2 wl_0_0 wl_1_0 vdd_uq1 bl_0_61 bl_1_61
+ br_0_61 br_1_61 sky130_fd_bd_sram__openram_dp_cell_dummy_2/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_2/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_2/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_2/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_14 wl_0_0 wl_1_0 vdd_uq13 bl_0_49 bl_1_49
+ br_0_49 br_1_49 sky130_fd_bd_sram__openram_dp_cell_dummy_14/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_14/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_14/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_14/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_25 wl_0_0 wl_1_0 vdd_uq24 bl_0_38 bl_1_38
+ br_0_38 br_1_38 sky130_fd_bd_sram__openram_dp_cell_dummy_25/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_25/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_25/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_25/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_36 wl_0_0 wl_1_0 vdd_uq35 bl_0_27 bl_1_27
+ br_0_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell_dummy_36/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_36/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_36/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_36/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_47 wl_0_0 wl_1_0 vdd_uq46 bl_0_16 bl_1_16
+ br_0_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell_dummy_47/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_47/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_47/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_47/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_58 wl_0_0 wl_1_0 vdd_uq57 bl_0_5 bl_1_5
+ br_0_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell_dummy_58/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_58/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_58/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_58/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_3 wl_0_0 wl_1_0 vdd_uq2 bl_0_60 bl_1_60
+ br_0_60 br_1_60 sky130_fd_bd_sram__openram_dp_cell_dummy_3/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_3/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_3/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_3/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_15 wl_0_0 wl_1_0 vdd_uq14 bl_0_48 bl_1_48
+ br_0_48 br_1_48 sky130_fd_bd_sram__openram_dp_cell_dummy_15/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_15/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_15/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_15/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_26 wl_0_0 wl_1_0 vdd_uq25 bl_0_37 bl_1_37
+ br_0_37 br_1_37 sky130_fd_bd_sram__openram_dp_cell_dummy_26/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_26/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_26/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_26/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_37 wl_0_0 wl_1_0 vdd_uq36 bl_0_26 bl_1_26
+ br_0_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell_dummy_37/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_37/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_37/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_37/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_48 wl_0_0 wl_1_0 vdd_uq47 bl_0_15 bl_1_15
+ br_0_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell_dummy_48/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_48/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_48/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_48/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_59 wl_0_0 wl_1_0 vdd_uq58 bl_0_4 bl_1_4
+ br_0_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell_dummy_59/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_59/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_59/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_59/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_4 wl_0_0 wl_1_0 vdd_uq3 bl_0_59 bl_1_59
+ br_0_59 br_1_59 sky130_fd_bd_sram__openram_dp_cell_dummy_4/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_4/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_4/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_4/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_16 wl_0_0 wl_1_0 vdd_uq15 bl_0_47 bl_1_47
+ br_0_47 br_1_47 sky130_fd_bd_sram__openram_dp_cell_dummy_16/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_16/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_16/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_16/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_27 wl_0_0 wl_1_0 vdd_uq26 bl_0_36 bl_1_36
+ br_0_36 br_1_36 sky130_fd_bd_sram__openram_dp_cell_dummy_27/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_27/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_27/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_27/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_38 wl_0_0 wl_1_0 vdd_uq37 bl_0_25 bl_1_25
+ br_0_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell_dummy_38/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_38/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_38/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_38/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_49 wl_0_0 wl_1_0 vdd_uq48 bl_0_14 bl_1_14
+ br_0_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell_dummy_49/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_49/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_49/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_49/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_5 wl_0_0 wl_1_0 vdd_uq4 bl_0_58 bl_1_58
+ br_0_58 br_1_58 sky130_fd_bd_sram__openram_dp_cell_dummy_5/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_5/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_5/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_5/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_6 wl_0_0 wl_1_0 vdd_uq5 bl_0_57 bl_1_57
+ br_0_57 br_1_57 sky130_fd_bd_sram__openram_dp_cell_dummy_6/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_6/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_6/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_6/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_17 wl_0_0 wl_1_0 vdd_uq16 bl_0_46 bl_1_46
+ br_0_46 br_1_46 sky130_fd_bd_sram__openram_dp_cell_dummy_17/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_17/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_17/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_17/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_28 wl_0_0 wl_1_0 vdd_uq27 bl_0_35 bl_1_35
+ br_0_35 br_1_35 sky130_fd_bd_sram__openram_dp_cell_dummy_28/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_28/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_28/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_28/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_39 wl_0_0 wl_1_0 vdd_uq38 bl_0_24 bl_1_24
+ br_0_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell_dummy_39/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_39/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_39/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_39/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_7 wl_0_0 wl_1_0 vdd_uq6 bl_0_56 bl_1_56
+ br_0_56 br_1_56 sky130_fd_bd_sram__openram_dp_cell_dummy_7/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_7/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_7/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_7/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_18 wl_0_0 wl_1_0 vdd_uq17 bl_0_45 bl_1_45
+ br_0_45 br_1_45 sky130_fd_bd_sram__openram_dp_cell_dummy_18/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_18/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_18/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_18/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_19 wl_0_0 wl_1_0 vdd_uq18 bl_0_44 bl_1_44
+ br_0_44 br_1_44 sky130_fd_bd_sram__openram_dp_cell_dummy_19/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_19/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_19/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_19/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_29 wl_0_0 wl_1_0 vdd_uq28 bl_0_34 bl_1_34
+ br_0_34 br_1_34 sky130_fd_bd_sram__openram_dp_cell_dummy_29/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_29/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_29/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_29/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_8 wl_0_0 wl_1_0 vdd_uq7 bl_0_55 bl_1_55
+ br_0_55 br_1_55 sky130_fd_bd_sram__openram_dp_cell_dummy_8/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_8/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_8/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_8/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_9 wl_0_0 wl_1_0 vdd_uq8 bl_0_54 bl_1_54
+ br_0_54 br_1_54 sky130_fd_bd_sram__openram_dp_cell_dummy_9/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_9/w_144_n79#
+ gnd sky130_fd_bd_sram__openram_dp_cell_dummy_9/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_9/VSUBS
+ sky130_fd_bd_sram__openram_dp_cell_dummy
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_replica_column wl_1_98 wl_1_99 wl_1_100
+ wl_1_106 wl_1_109 wl_1_112 wl_1_115 wl_1_118 wl_1_121 wl_1_123 wl_1_124 wl_1_127
+ wl_0_97 wl_0_103 wl_0_104 wl_0_105 wl_0_106 wl_0_107 wl_0_108 wl_0_109 wl_0_114
+ wl_0_115 wl_0_116 wl_0_117 wl_0_118 wl_0_119 wl_0_125 wl_0_126 wl_0_127 wl_0_128
+ wl_0_129 wl_1_97 wl_0_67 wl_0_70 wl_0_76 wl_0_82 wl_0_85 wl_0_91 wl_1_65 wl_1_66
+ wl_1_67 wl_1_68 wl_1_69 wl_1_70 wl_1_71 wl_1_72 wl_1_74 wl_1_75 wl_1_76 wl_1_77
+ wl_1_78 wl_1_79 wl_1_80 wl_1_81 wl_1_82 wl_1_83 wl_1_84 wl_1_85 wl_1_86 wl_1_87
+ wl_1_88 wl_1_91 wl_1_92 wl_1_93 wl_1_95 wl_1_96 wl_0_37 wl_0_38 wl_0_39 wl_0_48
+ wl_0_49 wl_0_55 wl_0_59 wl_0_60 wl_0_63 wl_1_32 wl_1_33 wl_1_35 wl_1_36 wl_1_38
+ wl_1_39 wl_1_40 wl_1_41 wl_1_42 wl_1_44 wl_1_45 wl_1_47 wl_1_48 wl_1_50 wl_1_51
+ wl_1_53 wl_1_54 wl_1_55 wl_1_56 wl_1_58 wl_1_59 wl_1_60 wl_1_61 wl_1_62 wl_1_63
+ wl_1_1 wl_1_2 wl_1_3 wl_1_6 wl_1_9 wl_1_10 wl_1_11 wl_1_12 wl_1_14 wl_1_15 wl_1_17
+ wl_1_18 wl_1_20 wl_1_21 wl_1_23 wl_1_24 wl_1_26 wl_1_27 wl_1_29 wl_1_30 wl_0_1 wl_0_2
+ wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_15 wl_0_16 wl_0_17 wl_0_18
+ wl_0_19 wl_0_26 wl_0_27 wl_0_28 wl_0_29 vdd wl_0_124 wl_0_88 wl_0_79 wl_0_36 wl_0_100
+ wl_0_30 wl_0_21 wl_0_12 wl_0_121 wl_0_112 wl_0_56 wl_0_51 wl_0_42 wl_0_93 wl_0_33
+ wl_0_24 wl_1_114 wl_1_105 wl_0_84 wl_0_75 wl_0_66 wl_0_123 wl_0_54 wl_0_45 wl_0_96
+ wl_1_8 wl_1_126 wl_1_117 wl_1_108 wl_0_87 wl_0_69 wl_0_78 wl_0_62 wl_0_99 wl_1_90
+ wl_1_120 wl_1_111 wl_1_102 wl_0_90 wl_0_81 wl_0_72 wl_0_47 wl_0_20 wl_0_11 wl_0_120
+ wl_0_111 wl_0_102 wl_1_129 wl_1_5 wl_0_50 wl_0_41 wl_0_32 wl_0_14 wl_0_23 wl_1_113
+ wl_1_104 wl_0_83 wl_0_74 wl_0_65 wl_0_58 wl_0_113 wl_0_53 wl_0_44 wl_0_35 wl_0_95
+ wl_1_16 wl_1_7 wl_1_125 wl_1_116 wl_1_107 wl_0_86 wl_0_77 wl_0_68 wl_0_61 wl_0_98
+ wl_1_89 wl_1_46 wl_1_0 wl_1_37 wl_1_28 wl_1_19 wl_1_128 wl_1_119 wl_1_110 wl_1_101
+ wl_0_89 wl_0_80 wl_0_71 wl_0_0 wl_0_46 wl_0_10 wl_0_110 wl_0_101 wl_1_49 wl_1_31
+ wl_1_22 wl_1_13 wl_1_4 wl_1_122 wl_0_92 wl_0_40 wl_0_31 wl_0_22 wl_0_13 wl_0_122
+ wl_1_73 wl_1_64 wl_1_57 wl_1_52 wl_1_103 wl_1_43 wl_1_94 wl_1_34 wl_1_25 wl_0_73
+ wl_0_64 wl_0_57 wl_0_52 wl_0_43 wl_0_34 wl_0_94 wl_0_25 bl_1_0 br_1_0 br_0_0 bl_0_0
+ gnd
Xsky130_fd_bd_sram__openram_dp_cell_replica_126 wl_0_66 wl_1_66 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_115 wl_0_77 wl_1_77 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_104 wl_0_88 wl_1_88 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_127 wl_0_65 wl_1_65 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_116 wl_0_76 wl_1_76 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_105 wl_0_87 wl_1_87 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_128 wl_0_64 wl_1_64 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_117 wl_0_75 wl_1_75 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_106 wl_0_86 wl_1_86 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_118 wl_0_74 wl_1_74 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_107 wl_0_85 wl_1_85 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_119 wl_0_73 wl_1_73 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_108 wl_0_84 wl_1_84 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_109 wl_0_83 wl_1_83 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_90 wl_0_102 wl_1_102 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_80 wl_0_112 wl_1_112 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_91 wl_0_101 wl_1_101 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_70 wl_0_122 wl_1_122 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_81 wl_0_111 wl_1_111 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_92 wl_0_100 wl_1_100 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_71 wl_0_121 wl_1_121 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_82 wl_0_110 wl_1_110 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_93 wl_0_99 wl_1_99 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_60 wl_0_5 wl_1_5 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_72 wl_0_120 wl_1_120 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_83 wl_0_109 wl_1_109 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_94 wl_0_98 wl_1_98 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_61 wl_0_4 wl_1_4 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_50 wl_0_15 wl_1_15 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_73 wl_0_119 wl_1_119 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_84 wl_0_108 wl_1_108 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_95 wl_0_97 wl_1_97 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_62 wl_0_3 wl_1_3 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_51 wl_0_14 wl_1_14 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_40 wl_0_25 wl_1_25 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_74 wl_0_118 wl_1_118 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_85 wl_0_107 wl_1_107 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_96 wl_0_96 wl_1_96 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_63 wl_0_2 wl_1_2 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_52 wl_0_13 wl_1_13 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_41 wl_0_24 wl_1_24 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_30 wl_0_35 wl_1_35 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_dummy_0 wl_0_129 wl_1_129 vdd bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_replica_64 wl_0_128 wl_1_128 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_75 wl_0_117 wl_1_117 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_86 wl_0_106 wl_1_106 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_97 wl_0_95 wl_1_95 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_53 wl_0_12 wl_1_12 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_42 wl_0_23 wl_1_23 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_31 wl_0_34 wl_1_34 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_20 wl_0_45 wl_1_45 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_65 wl_0_127 wl_1_127 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_76 wl_0_116 wl_1_116 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_87 wl_0_105 wl_1_105 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_54 wl_0_11 wl_1_11 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_43 wl_0_22 wl_1_22 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_32 wl_0_33 wl_1_33 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_21 wl_0_44 wl_1_44 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_10 wl_0_55 wl_1_55 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_98 wl_0_94 wl_1_94 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_66 wl_0_126 wl_1_126 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_77 wl_0_115 wl_1_115 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_88 wl_0_104 wl_1_104 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_55 wl_0_10 wl_1_10 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_44 wl_0_21 wl_1_21 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_33 wl_0_32 wl_1_32 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_22 wl_0_43 wl_1_43 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_11 wl_0_54 wl_1_54 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_99 wl_0_93 wl_1_93 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_67 wl_0_125 wl_1_125 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_78 wl_0_114 wl_1_114 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_89 wl_0_103 wl_1_103 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_56 wl_0_9 wl_1_9 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_45 wl_0_20 wl_1_20 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_34 wl_0_31 wl_1_31 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_23 wl_0_42 wl_1_42 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_12 wl_0_53 wl_1_53 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_68 wl_0_124 wl_1_124 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_79 wl_0_113 wl_1_113 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_57 wl_0_8 wl_1_8 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_46 wl_0_19 wl_1_19 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_35 wl_0_30 wl_1_30 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_24 wl_0_41 wl_1_41 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_13 wl_0_52 wl_1_52 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_69 wl_0_123 wl_1_123 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_58 wl_0_7 wl_1_7 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_47 wl_0_18 wl_1_18 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_36 wl_0_29 wl_1_29 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_25 wl_0_40 wl_1_40 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_14 wl_0_51 wl_1_51 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_0 wl_0_1 wl_1_1 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_59 wl_0_6 wl_1_6 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_48 wl_0_17 wl_1_17 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_37 wl_0_28 wl_1_28 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_26 wl_0_39 wl_1_39 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_15 wl_0_50 wl_1_50 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_1 wl_0_0 wl_1_0 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_49 wl_0_16 wl_1_16 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_38 wl_0_27 wl_1_27 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_27 wl_0_38 wl_1_38 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_16 wl_0_49 wl_1_49 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_39 wl_0_26 wl_1_26 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_28 wl_0_37 wl_1_37 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_17 wl_0_48 wl_1_48 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_2 wl_0_63 wl_1_63 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_3 wl_0_62 wl_1_62 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_29 wl_0_36 wl_1_36 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_18 wl_0_47 wl_1_47 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_19 wl_0_46 wl_1_46 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_4 wl_0_61 wl_1_61 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_5 wl_0_60 wl_1_60 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_6 wl_0_59 wl_1_59 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_7 wl_0_58 wl_1_58 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_120 wl_0_72 wl_1_72 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_8 wl_0_57 wl_1_57 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_121 wl_0_71 wl_1_71 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_110 wl_0_82 wl_1_82 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_9 wl_0_56 wl_1_56 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_122 wl_0_70 wl_1_70 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_111 wl_0_81 wl_1_81 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_100 wl_0_92 wl_1_92 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_123 wl_0_69 wl_1_69 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_112 wl_0_80 wl_1_80 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_101 wl_0_91 wl_1_91 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_124 wl_0_68 wl_1_68 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_113 wl_0_79 wl_1_79 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_102 wl_0_90 wl_1_90 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_125 wl_0_67 wl_1_67 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_114 wl_0_78 wl_1_78 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_103 wl_0_89 wl_1_89 bl_0_0 bl_1_0 br_0_0
+ br_1_0 bl_1_0 vdd gnd br_1_0 VSUBS sky130_fd_bd_sram__openram_dp_cell_replica
.ends

.subckt sky130_fd_bd_sram__openram_dp_cell wl0 wl1 bl0 bl1 br0 br1 a_38_n79# vdd gnd
+ a_400_n79#
X0 gnd gnd bl1 gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=80000u
X1 a_38_133# wl0 a_38_133# vdd sky130_fd_pr__special_pfet_pass ad=0p pd=0u as=0p ps=0u w=70000u l=150000u
X2 a_16_183# wl1 br1 gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
X3 gnd gnd a_400_n79# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=80000u
X4 a_16_183# a_38_133# gnd gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
X5 a_16_183# wl1 a_16_183# vdd sky130_fd_pr__special_pfet_pass ad=0p pd=0u as=0p ps=0u w=70000u l=150000u
X6 a_38_133# wl1 bl1 gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
X7 gnd gnd a_38_n79# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=80000u
X8 gnd gnd br1 gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=80000u
X9 a_38_133# a_16_183# gnd gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
X10 br0 wl0 a_16_183# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
X11 gnd a_38_133# a_16_183# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
X12 a_38_133# a_16_183# vdd vdd sky130_fd_pr__special_pfet_pass ad=0p pd=0u as=0p ps=0u w=140000u l=150000u
X13 vdd a_38_133# a_16_183# vdd sky130_fd_pr__special_pfet_pass ad=0p pd=0u as=0p ps=0u w=140000u l=150000u
X14 bl0 wl0 a_38_133# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
X15 gnd a_16_183# a_38_133# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_bitcell_array wl_0_125 wl_1_80 wl_1_81 wl_0_59
+ wl_0_48 wl_0_49 wl_1_51 wl_0_37 wl_0_28 wl_0_26 wl_0_19 wl_0_15 wl_0_4 br_1_30 br_0_19
+ bl_1_12 bl_1_4 bl_1_5 bl_1_56 bl_1_57 br_1_51 bl_1_45 br_1_40 br_1_41 bl_1_37 bl_1_34
+ gnd vdd vdd_uq99 vdd_uq190 vdd_uq254 vdd_uq318 vdd_uq382 vdd_uq446 vdd_uq510 vdd_uq574
+ vdd_uq638 vdd_uq702 vdd_uq766 vdd_uq830 vdd_uq894 vdd_uq958 vdd_uq999 vdd_uq1086
+ vdd_uq1150 vdd_uq1214 vdd_uq1278 vdd_uq1342 vdd_uq1470 vdd_uq1534 vdd_uq1598 vdd_uq1662
+ vdd_uq1726 vdd_uq1790 vdd_uq1918 vdd_uq2046 vdd_uq2110 vdd_uq2174 vdd_uq2238 vdd_uq2302
+ vdd_uq2366 vdd_uq2430 vdd_uq2494 vdd_uq2558 vdd_uq2622 vdd_uq2750 vdd_uq2814 vdd_uq2878
+ vdd_uq2942 vdd_uq3006 vdd_uq3070 vdd_uq3134 vdd_uq3198 vdd_uq3262 vdd_uq3326 vdd_uq3390
+ vdd_uq3454 vdd_uq3518 vdd_uq3582 vdd_uq3646 vdd_uq3710 vdd_uq3774 vdd_uq3902 vdd_uq3966
+ vdd_uq4030 vdd_uq4094 sky130_fd_bd_sram__openram_dp_cell_154/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_2487/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_6982/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_7479/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_7523/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_2099/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_7556/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_15/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_476/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_2099/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1974/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_8001/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_6953/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_5070/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5449/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_2452/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_7508/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_6963/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_184/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_7723/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5516/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_5126/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_2404/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_891/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_7076/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_2040/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_636/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_4990/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_5487/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5409/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_7003/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5003/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_607/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5778/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_21/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1972/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_3857/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_3790/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_7057/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_7523/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_5468/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_99/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_10/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5603/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_2414/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1904/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_7359/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_117/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_7476/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_8129/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_638/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_7431/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_166/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_413/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_5449/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5550/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_5584/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_2819/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_5013/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_2082/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_7412/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_2071/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_5075/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_2034/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_5603/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5070/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_5143/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_21/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_1993/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_8002/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_2101/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_2557/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_121/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_154/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_638/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_2130/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_6956/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_8001/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_5023/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_6956/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_5499/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5634/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_1974/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_7077/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_640/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_90/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_629/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_2470/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_4993/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_454/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_877/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_483/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_629/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_2082/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_5430/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_2379/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_2480/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_7360/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_7108/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_2040/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_2496/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5713/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_454/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5003/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_483/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_891/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_4993/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1904/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_2563/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_2563/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_6933/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_8002/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_2492/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5013/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_2415/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_7021/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1966/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5023/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_5421/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_2034/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_5533/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5018/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_497/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_484/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_7473/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_518/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_7039/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_2442/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_7473/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_2819/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_33/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1966/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_2452/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_7556/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_3857/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5092/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_5499/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5126/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_7056/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5533/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_5143/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_2108/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_1835/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_2487/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_90/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_7587/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_5210/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1972/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_2404/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_7076/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_184/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_7508/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_5778/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_2492/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_2414/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_6953/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_180/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_640/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_1/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_7057/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_7431/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_7497/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_7360/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_476/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_7393/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5109/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_6982/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_15/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_5038/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_4990/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_484/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5584/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_7077/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_7587/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_121/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_117/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_7412/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5516/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_2342/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_2415/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_7374/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_607/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_6963/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_7660/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_5409/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_2835/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_180/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5177/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_7359/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_636/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_5092/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_7393/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_33/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_99/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_5075/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_7003/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_5109/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5210/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_6911/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_2557/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_7039/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_2470/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_7476/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_7874/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_7723/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_497/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_413/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_2494/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_7488/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5567/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_7374/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5177/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_6911/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5430/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_7660/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5634/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_7874/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_3790/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_542/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_10/a_38_n79# wl_0_83 br_1_50 wl_1_28 sky130_fd_bd_sram__openram_dp_cell_2480/a_38_n79#
+ wl_1_19 wl_1_113 wl_1_4 wl_1_0 br_0_50 wl_1_98 sky130_fd_bd_sram__openram_dp_cell_5018/a_400_n79#
+ wl_1_46 sky130_fd_bd_sram__openram_dp_cell_604/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_166/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_5567/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_2130/a_400_n79#
+ wl_0_67 wl_0_113 sky130_fd_bd_sram__openram_dp_cell_7497/a_400_n79# wl_1_86 wl_0_78
+ bl_0_34 sky130_fd_bd_sram__openram_dp_cell_8129/a_400_n79# wl_0_0 sky130_fd_bd_sram__openram_dp_cell_1835/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_877/a_400_n79# wl_0_98 wl_1_40 wl_0_60 bl_0_10
+ wl_0_46 sky130_fd_bd_sram__openram_dp_cell_2101/a_400_n79# wl_1_58 wl_1_107 sky130_fd_bd_sram__openram_dp_cell_2071/a_38_n79#
+ bl_1_50 sky130_fd_bd_sram__openram_dp_cell_2494/a_38_n79# wl_1_49 wl_1_10 wl_0_9
+ sky130_fd_bd_sram__openram_dp_cell_2835/a_400_n79# wl_1_76 wl_1_64 wl_0_65 sky130_fd_bd_sram__openram_dp_cell_2379/a_38_n79#
+ wl_0_86 bl_0_23 sky130_fd_bd_sram__openram_dp_cell_5038/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_7056/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_7479/a_38_n79# wl_1_43 bl_0_37 wl_1_123 wl_0_40
+ bl_0_56 sky130_fd_bd_sram__openram_dp_cell_5421/a_38_n79# bl_1_16 wl_0_58 wl_1_125
+ wl_0_107 sky130_fd_bd_sram__openram_dp_cell_5487/a_38_n79# bl_0_50 wl_0_10 wl_1_116
+ wl_1_97 br_1_21 wl_0_29 br_1_38 wl_1_13 bl_0_1 wl_0_8 wl_0_34 bl_0_7 wl_0_76 wl_0_63
+ wl_0_95 br_0_52 br_1_18 wl_0_64 sky130_fd_bd_sram__openram_dp_cell_2342/a_38_n79#
+ bl_1_6 bl_1_31 bl_0_45 wl_0_93 br_1_25 bl_0_2 wl_1_75 wl_1_20 wl_1_29 bl_1_42 wl_0_43
+ br_1_4 bl_0_53 wl_1_110 br_0_8 sky130_fd_bd_sram__openram_dp_cell_2496/a_400_n79#
+ bl_0_40 wl_1_36 br_0_32 wl_0_22 wl_0_74 bl_1_63 wl_1_120 vdd_uq2686 wl_0_123 bl_0_58
+ wl_1_54 bl_1_51 bl_1_49 wl_0_69 bl_0_8 bl_1_61 wl_1_56 sky130_fd_bd_sram__openram_dp_cell_7488/a_400_n79#
+ br_1_45 wl_0_106 br_0_56 sky130_fd_bd_sram__openram_dp_cell_604/a_38_n79# wl_1_79
+ bl_0_35 br_1_60 wl_1_101 bl_0_16 wl_1_35 bl_0_43 wl_0_104 wl_0_105 bl_1_0 br_1_2
+ wl_1_100 wl_0_116 wl_0_108 wl_1_42 bl_1_3 wl_0_97 br_1_9 wl_1_31 br_1_59 wl_0_7
+ wl_1_90 wl_0_52 br_1_31 wl_1_119 wl_1_114 br_1_0 wl_1_99 br_1_12 br_0_26 br_0_24
+ bl_0_44 br_0_21 br_1_39 sky130_fd_bd_sram__openram_dp_cell_2442/a_38_n79# wl_1_111
+ br_0_38 wl_1_84 wl_0_13 br_0_36 wl_1_89 br_0_37 bl_1_39 br_1_58 bl_1_27 bl_1_20
+ wl_1_9 bl_0_14 bl_0_47 bl_0_25 wl_0_32 wl_1_68 bl_0_5 bl_0_17 wl_1_17 wl_0_25 br_0_18
+ br_1_16 wl_1_77 br_1_53 bl_0_9 bl_0_6 bl_1_46 bl_0_59 bl_0_31 bl_1_38 br_1_63 br_0_33
+ wl_1_27 wl_1_2 br_0_42 wl_1_12 bl_1_41 br_0_28 bl_1_19 wl_0_47 bl_1_18 wl_0_87 br_0_23
+ br_0_25 wl_0_66 bl_0_13 wl_0_6 wl_1_3 wl_0_45 wl_1_117 wl_1_1 wl_1_112 wl_0_75 wl_0_20
+ sky130_fd_bd_sram__openram_dp_cell_7108/a_38_n79# bl_1_33 wl_0_38 br_1_3 wl_1_50
+ bl_0_42 wl_1_11 wl_0_36 wl_1_103 br_1_20 br_0_30 wl_0_61 wl_0_16 bl_0_4 wl_0_55
+ br_0_4 wl_1_32 wl_1_122 wl_1_14 wl_1_18 wl_0_110 wl_1_108 bl_1_30 sky130_fd_bd_sram__openram_dp_cell_1993/a_38_n79#
+ bl_0_60 wl_0_57 bl_1_17 bl_0_11 br_0_43 wl_1_126 br_1_43 wl_1_30 bl_0_54 wl_0_24
+ br_1_23 bl_0_32 br_0_6 bl_0_63 br_1_26 wl_1_87 wl_0_80 br_1_29 br_0_34 br_0_47 wl_0_120
+ br_1_49 br_1_46 bl_0_12 bl_1_7 wl_1_88 br_1_35 sky130_fd_bd_sram__openram_dp_cell_5550/a_38_n79#
+ wl_0_54 wl_1_109 bl_0_51 bl_0_49 br_1_44 bl_1_35 wl_0_71 wl_1_105 br_0_11 wl_1_121
+ br_0_41 wl_1_45 wl_0_94 bl_0_62 bl_1_48 wl_1_24 wl_1_63 wl_1_61 wl_1_62 wl_0_127
+ bl_1_32 bl_0_61 br_0_31 wl_1_106 br_0_29 wl_0_56 br_1_34 bl_0_48 br_0_45 br_1_27
+ wl_0_51 wl_0_85 br_1_22 wl_1_52 wl_0_102 br_0_14 wl_1_78 wl_0_118 br_1_19 wl_1_5
+ wl_0_5 br_0_51 wl_0_88 wl_0_44 br_0_46 bl_1_15 wl_0_79 br_0_48 br_0_60 wl_0_101
+ wl_1_92 wl_0_70 wl_0_109 sky130_fd_bd_sram__openram_dp_cell_542/a_400_n79# wl_1_94
+ wl_1_47 wl_0_35 wl_1_60 wl_0_33 wl_0_62 wl_1_127 br_1_42 br_0_10 bl_1_14 wl_1_83
+ wl_1_33 bl_0_0 wl_0_100 br_0_2 wl_1_104 wl_1_85 br_1_17 wl_0_92 wl_0_42 vdd_uq1406
+ wl_0_39 br_0_61 bl_0_3 wl_1_7 wl_1_95 br_0_54 wl_0_53 bl_0_52 br_0_9 wl_0_31 br_0_13
+ br_0_59 br_1_7 bl_1_10 wl_0_90 bl_1_47 bl_1_52 bl_1_11 br_1_24 bl_1_36 wl_0_119
+ bl_0_24 bl_1_55 bl_0_28 br_0_49 wl_1_102 wl_0_114 wl_1_53 sky130_fd_bd_sram__openram_dp_cell_2108/a_38_n79#
+ br_1_28 br_0_0 wl_0_99 br_0_12 wl_0_72 wl_1_23 br_1_8 wl_0_81 bl_0_15 br_0_39 wl_0_111
+ br_1_33 bl_1_53 wl_1_8 br_1_57 bl_0_26 br_1_10 br_0_57 wl_0_84 br_1_55 wl_0_89 wl_0_122
+ bl_1_13 bl_0_29 bl_0_39 br_1_62 wl_0_73 br_0_7 wl_1_74 br_0_58 bl_0_27 br_0_55 sky130_fd_bd_sram__openram_dp_cell_5468/a_38_n79#
+ bl_1_1 wl_0_14 bl_0_20 wl_1_59 br_1_5 wl_1_70 bl_1_24 wl_1_26 wl_0_68 bl_0_30 wl_1_65
+ sky130_fd_bd_sram__openram_dp_cell_5713/a_400_n79# bl_1_9 br_1_32 wl_0_91 bl_1_8
+ br_1_61 br_1_37 br_0_5 bl_0_57 wl_0_17 wl_1_38 wl_1_91 br_1_47 bl_1_54 wl_1_66 bl_0_36
+ wl_1_71 br_0_16 bl_0_21 br_1_48 wl_1_41 wl_1_22 wl_0_77 wl_0_82 br_0_53 wl_0_23
+ bl_1_2 bl_1_26 br_1_56 wl_0_21 wl_1_82 wl_1_44 bl_0_46 br_1_11 br_1_13 bl_0_38 wl_1_118
+ br_0_63 wl_1_6 br_0_1 bl_1_62 bl_1_22 sky130_fd_bd_sram__openram_dp_cell_518/a_38_n79#
+ wl_1_21 wl_1_39 wl_0_27 wl_1_93 wl_1_124 wl_0_2 br_0_27 bl_1_25 wl_0_12 wl_1_73
+ wl_0_126 sky130_fd_bd_sram__openram_dp_cell_7021/a_400_n79# bl_1_43 bl_0_41 wl_1_69
+ br_1_52 bl_0_19 wl_0_96 br_0_22 wl_0_41 br_0_62 bl_0_22 bl_0_18 bl_1_21 vdd_uq1982
+ br_1_14 br_1_6 wl_0_18 wl_1_34 wl_1_48 wl_1_115 bl_1_59 wl_0_3 br_0_15 wl_0_117
+ wl_0_121 wl_1_96 br_1_15 wl_0_1 wl_0_112 br_1_36 wl_0_124 bl_0_33 bl_1_40 br_0_3
+ bl_1_29 wl_1_25 wl_1_72 br_0_40 wl_1_15 wl_1_37 br_0_17 wl_0_30 br_0_35 br_1_54
+ wl_0_50 wl_1_57 vdd_uq3838 wl_0_11 bl_1_58 sky130_fd_bd_sram__openram_dp_cell_6933/a_400_n79#
+ bl_1_28 br_0_44 bl_1_23 bl_1_44 wl_0_103 br_0_20 bl_1_60 bl_0_55 wl_1_55 wl_0_115
+ wl_1_16 vdd_uq1854 wl_1_67 br_1_1
Xsky130_fd_bd_sram__openram_dp_cell_7215 wl_0_108 wl_1_108 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7204 wl_0_101 wl_1_101 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7248 wl_0_108 wl_1_108 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7237 wl_0_106 wl_1_106 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7226 wl_0_97 wl_1_97 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6503 wl_0_87 wl_1_87 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5802 wl_0_103 wl_1_103 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7259 wl_0_97 wl_1_97 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6547 wl_0_81 wl_1_81 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6514 wl_0_84 wl_1_84 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6525 wl_0_85 wl_1_85 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6536 wl_0_92 wl_1_92 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5835 wl_0_70 wl_1_70 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5824 wl_0_81 wl_1_81 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6558 wl_0_86 wl_1_86 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5813 wl_0_92 wl_1_92 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6569 wl_0_91 wl_1_91 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5868 wl_0_72 wl_1_72 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5857 wl_0_96 wl_1_96 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5846 wl_0_95 wl_1_95 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5879 wl_0_77 wl_1_77 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7771 wl_0_79 wl_1_79 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7760 wl_0_90 wl_1_90 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7793 wl_0_95 wl_1_95 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7782 wl_0_68 wl_1_68 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_240 wl_0_22 wl_1_22 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_251 wl_0_18 wl_1_18 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_273 wl_0_26 wl_1_26 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_262 wl_0_27 wl_1_27 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_295 wl_0_25 wl_1_25 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_284 wl_0_28 wl_1_28 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5109 wl_0_127 wl_1_127 bl_0_12 bl_1_12 br_0_12
+ br_1_12 sky130_fd_bd_sram__openram_dp_cell_5109/a_38_n79# vdd_uq3326 gnd sky130_fd_bd_sram__openram_dp_cell_5109/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4419 wl_0_67 wl_1_67 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4408 wl_0_77 wl_1_77 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3718 wl_0_46 wl_1_46 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3707 wl_0_57 wl_1_57 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3729 wl_0_61 wl_1_61 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7023 wl_0_125 wl_1_125 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7001 wl_0_122 wl_1_122 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7012 wl_0_118 wl_1_118 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7056 wl_0_127 wl_1_127 bl_0_41 bl_1_41 br_0_41
+ br_1_41 sky130_fd_bd_sram__openram_dp_cell_7056/a_38_n79# vdd_uq1470 gnd sky130_fd_bd_sram__openram_dp_cell_7056/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7045 wl_0_121 wl_1_121 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7034 wl_0_114 wl_1_114 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6311 wl_0_70 wl_1_70 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6300 wl_0_79 wl_1_79 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7078 wl_0_126 wl_1_126 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5610 wl_0_120 wl_1_120 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7067 wl_0_117 wl_1_117 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7089 wl_0_115 wl_1_115 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6355 wl_0_67 wl_1_67 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6322 wl_0_70 wl_1_70 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6344 wl_0_73 wl_1_73 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6333 wl_0_75 wl_1_75 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5643 wl_0_118 wl_1_118 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5621 wl_0_109 wl_1_109 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5632 wl_0_98 wl_1_98 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6366 wl_0_69 wl_1_69 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6377 wl_0_69 wl_1_69 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6388 wl_0_73 wl_1_73 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5665 wl_0_112 wl_1_112 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4931 wl_0_110 wl_1_110 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5654 wl_0_107 wl_1_107 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4920 wl_0_101 wl_1_101 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4942 wl_0_101 wl_1_101 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6399 wl_0_75 wl_1_75 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5676 wl_0_95 wl_1_95 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4975 wl_0_117 wl_1_117 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4964 wl_0_116 wl_1_116 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4953 wl_0_104 wl_1_104 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5698 wl_0_95 wl_1_95 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5687 wl_0_96 wl_1_96 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4997 wl_0_123 wl_1_123 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4986 wl_0_115 wl_1_115 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7590 wl_0_124 wl_1_124 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4227 wl_0_85 wl_1_85 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4216 wl_0_86 wl_1_86 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4205 wl_0_90 wl_1_90 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3515 wl_0_49 wl_1_49 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3526 wl_0_56 wl_1_56 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3504 wl_0_60 wl_1_60 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4249 wl_0_89 wl_1_89 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4238 wl_0_94 wl_1_94 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2803 wl_0_17 wl_1_17 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2814 wl_0_5 wl_1_5 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3548 wl_0_50 wl_1_50 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3559 wl_0_59 wl_1_59 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3537 wl_0_61 wl_1_61 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2836 wl_0_16 wl_1_16 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2847 wl_0_15 wl_1_15 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2825 wl_0_10 wl_1_10 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2869 wl_0_36 wl_1_36 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2858 wl_0_44 wl_1_44 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6130 wl_0_91 wl_1_91 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6152 wl_0_81 wl_1_81 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6163 wl_0_85 wl_1_85 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6141 wl_0_88 wl_1_88 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5440 wl_0_119 wl_1_119 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5451 wl_0_119 wl_1_119 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6185 wl_0_82 wl_1_82 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6196 wl_0_89 wl_1_89 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6174 wl_0_93 wl_1_93 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5473 wl_0_124 wl_1_124 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5495 wl_0_121 wl_1_121 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5462 wl_0_116 wl_1_116 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5484 wl_0_113 wl_1_113 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4750 wl_0_82 wl_1_82 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4783 wl_0_102 wl_1_102 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4761 wl_0_71 wl_1_71 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4772 wl_0_80 wl_1_80 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4794 wl_0_101 wl_1_101 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1409 wl_0_44 wl_1_44 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_806 wl_0_28 wl_1_28 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4002 wl_0_66 wl_1_66 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_839 wl_0_16 wl_1_16 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_817 wl_0_16 wl_1_16 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_828 wl_0_27 wl_1_27 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3301 wl_0_47 wl_1_47 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4024 wl_0_65 wl_1_65 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4013 wl_0_71 wl_1_71 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4035 wl_0_76 wl_1_76 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3323 wl_0_35 wl_1_35 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3334 wl_0_40 wl_1_40 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3312 wl_0_46 wl_1_46 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4046 wl_0_67 wl_1_67 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4057 wl_0_70 wl_1_70 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4068 wl_0_74 wl_1_74 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4079 wl_0_94 wl_1_94 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2600 wl_0_23 wl_1_23 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2622 wl_0_21 wl_1_21 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2611 wl_0_27 wl_1_27 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3356 wl_0_36 wl_1_36 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3367 wl_0_37 wl_1_37 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3345 wl_0_45 wl_1_45 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2633 wl_0_23 wl_1_23 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2655 wl_0_22 wl_1_22 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2666 wl_0_18 wl_1_18 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2644 wl_0_26 wl_1_26 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1910 wl_0_31 wl_1_31 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1921 wl_0_32 wl_1_32 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3389 wl_0_36 wl_1_36 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3378 wl_0_36 wl_1_36 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2677 wl_0_20 wl_1_20 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1954 wl_0_12 wl_1_12 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2699 wl_0_27 wl_1_27 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2688 wl_0_29 wl_1_29 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1932 wl_0_31 wl_1_31 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1943 wl_0_32 wl_1_32 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1976 wl_0_14 wl_1_14 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1987 wl_0_6 wl_1_6 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1965 wl_0_1 wl_1_1 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1998 wl_0_11 wl_1_11 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5270 wl_0_108 wl_1_108 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5292 wl_0_106 wl_1_106 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5281 wl_0_97 wl_1_97 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4580 wl_0_92 wl_1_92 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4591 wl_0_93 wl_1_93 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3890 wl_0_32 wl_1_32 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1217 wl_0_51 wl_1_51 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1206 wl_0_59 wl_1_59 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1239 wl_0_53 wl_1_53 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1228 wl_0_58 wl_1_58 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_614 wl_0_11 wl_1_11 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_603 wl_0_1 wl_1_1 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_636 wl_0_0 wl_1_0 bl_0_35 bl_1_35 br_0_35 br_1_35
+ sky130_fd_bd_sram__openram_dp_cell_636/a_38_n79# vdd_uq1854 gnd sky130_fd_bd_sram__openram_dp_cell_636/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_625 wl_0_4 wl_1_4 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_647 wl_0_28 wl_1_28 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_669 wl_0_21 wl_1_21 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_658 wl_0_28 wl_1_28 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3131 wl_0_53 wl_1_53 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3142 wl_0_53 wl_1_53 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3120 wl_0_57 wl_1_57 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2430 wl_0_12 wl_1_12 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2441 wl_0_1 wl_1_1 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3164 wl_0_51 wl_1_51 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3153 wl_0_57 wl_1_57 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3175 wl_0_57 wl_1_57 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2463 wl_0_7 wl_1_7 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2452 wl_0_0 wl_1_0 bl_0_11 bl_1_11 br_0_11 br_1_11
+ sky130_fd_bd_sram__openram_dp_cell_2452/a_38_n79# vdd_uq3390 gnd sky130_fd_bd_sram__openram_dp_cell_2452/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2474 wl_0_1 wl_1_1 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3186 wl_0_54 wl_1_54 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3197 wl_0_61 wl_1_61 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2485 wl_0_1 wl_1_1 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2496 wl_0_0 wl_1_0 bl_0_0 bl_1_0 br_0_0 br_1_0
+ sky130_fd_bd_sram__openram_dp_cell_2496/a_38_n79# vdd_uq4094 gnd sky130_fd_bd_sram__openram_dp_cell_2496/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1762 wl_0_37 wl_1_37 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1751 wl_0_48 wl_1_48 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1740 wl_0_59 wl_1_59 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1795 wl_0_38 wl_1_38 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1784 wl_0_49 wl_1_49 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1773 wl_0_60 wl_1_60 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8109 wl_0_20 wl_1_20 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7419 wl_0_118 wl_1_118 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7408 wl_0_114 wl_1_114 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6729 wl_0_99 wl_1_99 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6718 wl_0_76 wl_1_76 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6707 wl_0_87 wl_1_87 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1014 wl_0_34 wl_1_34 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1003 wl_0_41 wl_1_41 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1025 wl_0_43 wl_1_43 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1036 wl_0_35 wl_1_35 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1058 wl_0_42 wl_1_42 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1047 wl_0_43 wl_1_43 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1069 wl_0_59 wl_1_59 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7920 wl_0_81 wl_1_81 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7953 wl_0_48 wl_1_48 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7942 wl_0_59 wl_1_59 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7931 wl_0_70 wl_1_70 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7986 wl_0_15 wl_1_15 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7975 wl_0_26 wl_1_26 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7964 wl_0_37 wl_1_37 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7997 wl_0_4 wl_1_4 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_411 wl_0_16 wl_1_16 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_422 wl_0_16 wl_1_16 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_400 wl_0_9 wl_1_9 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_433 wl_0_21 wl_1_21 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_455 wl_0_16 wl_1_16 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_444 wl_0_10 wl_1_10 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_499 wl_0_9 wl_1_9 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_488 wl_0_6 wl_1_6 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_477 wl_0_6 wl_1_6 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_466 wl_0_5 wl_1_5 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2260 wl_0_23 wl_1_23 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2282 wl_0_20 wl_1_20 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2271 wl_0_27 wl_1_27 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2293 wl_0_26 wl_1_26 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1581 wl_0_53 wl_1_53 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1570 wl_0_62 wl_1_62 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1592 wl_0_57 wl_1_57 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7205 wl_0_100 wl_1_100 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7216 wl_0_107 wl_1_107 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7249 wl_0_107 wl_1_107 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7227 wl_0_107 wl_1_107 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7238 wl_0_105 wl_1_105 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6504 wl_0_86 wl_1_86 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6515 wl_0_83 wl_1_83 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6526 wl_0_84 wl_1_84 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6537 wl_0_91 wl_1_91 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5803 wl_0_102 wl_1_102 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5825 wl_0_80 wl_1_80 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6548 wl_0_82 wl_1_82 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6559 wl_0_85 wl_1_85 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5814 wl_0_91 wl_1_91 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5836 wl_0_69 wl_1_69 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5869 wl_0_71 wl_1_71 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5858 wl_0_95 wl_1_95 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5847 wl_0_96 wl_1_96 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7750 wl_0_100 wl_1_100 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7761 wl_0_89 wl_1_89 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7794 wl_0_96 wl_1_96 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7783 wl_0_67 wl_1_67 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7772 wl_0_78 wl_1_78 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_230 wl_0_24 wl_1_24 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_241 wl_0_21 wl_1_21 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_263 wl_0_19 wl_1_19 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_252 wl_0_17 wl_1_17 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_274 wl_0_25 wl_1_25 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_296 wl_0_24 wl_1_24 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_285 wl_0_27 wl_1_27 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2090 wl_0_8 wl_1_8 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4409 wl_0_70 wl_1_70 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3708 wl_0_56 wl_1_56 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3719 wl_0_45 wl_1_45 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7002 wl_0_121 wl_1_121 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7013 wl_0_117 wl_1_117 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7057 wl_0_127 wl_1_127 bl_0_46 bl_1_46 br_0_46
+ br_1_46 sky130_fd_bd_sram__openram_dp_cell_7057/a_38_n79# vdd_uq1150 gnd sky130_fd_bd_sram__openram_dp_cell_7057/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7024 wl_0_124 wl_1_124 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7046 wl_0_120 wl_1_120 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7035 wl_0_113 wl_1_113 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6312 wl_0_69 wl_1_69 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6301 wl_0_80 wl_1_80 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7079 wl_0_125 wl_1_125 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7068 wl_0_116 wl_1_116 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5600 wl_0_111 wl_1_111 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6323 wl_0_69 wl_1_69 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6345 wl_0_72 wl_1_72 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6334 wl_0_74 wl_1_74 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5611 wl_0_119 wl_1_119 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5644 wl_0_117 wl_1_117 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5622 wl_0_108 wl_1_108 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5633 wl_0_97 wl_1_97 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6356 wl_0_66 wl_1_66 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6367 wl_0_68 wl_1_68 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6378 wl_0_68 wl_1_68 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6389 wl_0_78 wl_1_78 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5666 wl_0_111 wl_1_111 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4932 wl_0_109 wl_1_109 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5655 wl_0_106 wl_1_106 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4910 wl_0_100 wl_1_100 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4921 wl_0_99 wl_1_99 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5677 wl_0_96 wl_1_96 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4965 wl_0_115 wl_1_115 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4954 wl_0_103 wl_1_103 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4943 wl_0_100 wl_1_100 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5699 wl_0_96 wl_1_96 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5688 wl_0_95 wl_1_95 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4998 wl_0_122 wl_1_122 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4976 wl_0_116 wl_1_116 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4987 wl_0_114 wl_1_114 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7591 wl_0_123 wl_1_123 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7580 wl_0_103 wl_1_103 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6890 wl_0_107 wl_1_107 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4228 wl_0_84 wl_1_84 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4217 wl_0_85 wl_1_85 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4206 wl_0_89 wl_1_89 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3516 wl_0_58 wl_1_58 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3505 wl_0_59 wl_1_59 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4239 wl_0_93 wl_1_93 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2804 wl_0_16 wl_1_16 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2815 wl_0_4 wl_1_4 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3549 wl_0_49 wl_1_49 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3527 wl_0_55 wl_1_55 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3538 wl_0_60 wl_1_60 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2848 wl_0_16 wl_1_16 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2837 wl_0_15 wl_1_15 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2826 wl_0_9 wl_1_9 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2859 wl_0_46 wl_1_46 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6120 wl_0_83 wl_1_83 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6142 wl_0_87 wl_1_87 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6131 wl_0_90 wl_1_90 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6153 wl_0_94 wl_1_94 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5430 wl_0_127 wl_1_127 bl_0_22 bl_1_22 br_0_22
+ br_1_22 sky130_fd_bd_sram__openram_dp_cell_5430/a_38_n79# vdd_uq2686 gnd sky130_fd_bd_sram__openram_dp_cell_5430/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5452 wl_0_126 wl_1_126 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5441 wl_0_118 wl_1_118 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6186 wl_0_81 wl_1_81 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6164 wl_0_84 wl_1_84 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6197 wl_0_88 wl_1_88 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6175 wl_0_92 wl_1_92 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5474 wl_0_123 wl_1_123 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5463 wl_0_115 wl_1_115 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5485 wl_0_116 wl_1_116 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4740 wl_0_92 wl_1_92 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5496 wl_0_120 wl_1_120 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4784 wl_0_101 wl_1_101 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4762 wl_0_70 wl_1_70 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4773 wl_0_79 wl_1_79 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4751 wl_0_81 wl_1_81 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4795 wl_0_100 wl_1_100 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4003 wl_0_65 wl_1_65 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_818 wl_0_15 wl_1_15 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_829 wl_0_26 wl_1_26 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_807 wl_0_27 wl_1_27 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4025 wl_0_69 wl_1_69 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4014 wl_0_70 wl_1_70 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4036 wl_0_75 wl_1_75 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3324 wl_0_34 wl_1_34 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3302 wl_0_40 wl_1_40 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3313 wl_0_45 wl_1_45 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4047 wl_0_66 wl_1_66 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4058 wl_0_69 wl_1_69 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4069 wl_0_73 wl_1_73 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2601 wl_0_22 wl_1_22 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2623 wl_0_20 wl_1_20 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2612 wl_0_26 wl_1_26 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3357 wl_0_35 wl_1_35 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3335 wl_0_39 wl_1_39 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3346 wl_0_46 wl_1_46 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3368 wl_0_46 wl_1_46 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2634 wl_0_22 wl_1_22 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2656 wl_0_21 wl_1_21 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1900 wl_0_4 wl_1_4 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2645 wl_0_25 wl_1_25 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1911 wl_0_32 wl_1_32 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3379 wl_0_35 wl_1_35 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2678 wl_0_19 wl_1_19 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2667 wl_0_19 wl_1_19 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1955 wl_0_11 wl_1_11 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2689 wl_0_28 wl_1_28 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1933 wl_0_32 wl_1_32 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1944 wl_0_31 wl_1_31 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1922 wl_0_31 wl_1_31 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1977 wl_0_13 wl_1_13 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1966 wl_0_0 wl_1_0 bl_0_29 bl_1_29 br_0_29 br_1_29
+ sky130_fd_bd_sram__openram_dp_cell_1966/a_38_n79# vdd_uq2238 gnd sky130_fd_bd_sram__openram_dp_cell_1966/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1988 wl_0_5 wl_1_5 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1999 wl_0_10 wl_1_10 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5260 wl_0_100 wl_1_100 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5271 wl_0_107 wl_1_107 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5282 wl_0_107 wl_1_107 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5293 wl_0_105 wl_1_105 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4570 wl_0_90 wl_1_90 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4592 wl_0_92 wl_1_92 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4581 wl_0_91 wl_1_91 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3880 wl_0_32 wl_1_32 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3891 wl_0_32 wl_1_32 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1207 wl_0_58 wl_1_58 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1218 wl_0_50 wl_1_50 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1229 wl_0_57 wl_1_57 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_604 wl_0_0 wl_1_0 bl_0_36 bl_1_36 br_0_36 br_1_36
+ sky130_fd_bd_sram__openram_dp_cell_604/a_38_n79# vdd_uq1790 gnd sky130_fd_bd_sram__openram_dp_cell_604/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_615 wl_0_10 wl_1_10 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_637 wl_0_1 wl_1_1 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_626 wl_0_3 wl_1_3 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_648 wl_0_27 wl_1_27 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_659 wl_0_27 wl_1_27 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3143 wl_0_52 wl_1_52 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3121 wl_0_56 wl_1_56 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3110 wl_0_57 wl_1_57 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3132 wl_0_58 wl_1_58 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2431 wl_0_11 wl_1_11 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2420 wl_0_10 wl_1_10 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3165 wl_0_50 wl_1_50 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3176 wl_0_56 wl_1_56 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3154 wl_0_61 wl_1_61 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2453 wl_0_14 wl_1_14 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2464 wl_0_6 wl_1_6 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2442 wl_0_0 wl_1_0 bl_0_12 bl_1_12 br_0_12 br_1_12
+ sky130_fd_bd_sram__openram_dp_cell_2442/a_38_n79# vdd_uq3326 gnd sky130_fd_bd_sram__openram_dp_cell_2442/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1730 wl_0_39 wl_1_39 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3187 wl_0_53 wl_1_53 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3198 wl_0_60 wl_1_60 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2475 wl_0_14 wl_1_14 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2497 wl_0_3 wl_1_3 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2486 wl_0_4 wl_1_4 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1763 wl_0_36 wl_1_36 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1752 wl_0_47 wl_1_47 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1741 wl_0_58 wl_1_58 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1796 wl_0_37 wl_1_37 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1785 wl_0_48 wl_1_48 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1774 wl_0_59 wl_1_59 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5090 wl_0_122 wl_1_122 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7409 wl_0_113 wl_1_113 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6719 wl_0_75 wl_1_75 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6708 wl_0_86 wl_1_86 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1015 wl_0_33 wl_1_33 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1004 wl_0_40 wl_1_40 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1037 wl_0_34 wl_1_34 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1059 wl_0_41 wl_1_41 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1026 wl_0_42 wl_1_42 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1048 wl_0_46 wl_1_46 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7910 wl_0_91 wl_1_91 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7943 wl_0_58 wl_1_58 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7932 wl_0_69 wl_1_69 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7921 wl_0_80 wl_1_80 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7987 wl_0_14 wl_1_14 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7976 wl_0_25 wl_1_25 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7965 wl_0_36 wl_1_36 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7954 wl_0_47 wl_1_47 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7998 wl_0_3 wl_1_3 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_412 wl_0_15 wl_1_15 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_423 wl_0_15 wl_1_15 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_401 wl_0_8 wl_1_8 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_434 wl_0_20 wl_1_20 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_456 wl_0_15 wl_1_15 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_445 wl_0_9 wl_1_9 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_467 wl_0_4 wl_1_4 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_478 wl_0_5 wl_1_5 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_489 wl_0_5 wl_1_5 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2250 wl_0_24 wl_1_24 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2261 wl_0_22 wl_1_22 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2283 wl_0_19 wl_1_19 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2272 wl_0_26 wl_1_26 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2294 wl_0_25 wl_1_25 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1560 wl_0_55 wl_1_55 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1571 wl_0_62 wl_1_62 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1582 wl_0_52 wl_1_52 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1593 wl_0_56 wl_1_56 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_990 wl_0_44 wl_1_44 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7206 wl_0_99 wl_1_99 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7217 wl_0_106 wl_1_106 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7228 wl_0_106 wl_1_106 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7239 wl_0_104 wl_1_104 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6527 wl_0_83 wl_1_83 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6505 wl_0_85 wl_1_85 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6538 wl_0_90 wl_1_90 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6516 wl_0_94 wl_1_94 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5804 wl_0_101 wl_1_101 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5826 wl_0_79 wl_1_79 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6549 wl_0_81 wl_1_81 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5815 wl_0_90 wl_1_90 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5837 wl_0_68 wl_1_68 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5859 wl_0_67 wl_1_67 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5848 wl_0_95 wl_1_95 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7740 wl_0_110 wl_1_110 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7751 wl_0_99 wl_1_99 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7762 wl_0_88 wl_1_88 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7795 wl_0_95 wl_1_95 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7784 wl_0_66 wl_1_66 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7773 wl_0_77 wl_1_77 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_231 wl_0_23 wl_1_23 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_220 wl_0_27 wl_1_27 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_242 wl_0_20 wl_1_20 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_264 wl_0_18 wl_1_18 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_253 wl_0_26 wl_1_26 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_275 wl_0_24 wl_1_24 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_297 wl_0_23 wl_1_23 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_286 wl_0_26 wl_1_26 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2091 wl_0_7 wl_1_7 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2080 wl_0_2 wl_1_2 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1390 wl_0_43 wl_1_43 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3709 wl_0_55 wl_1_55 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7003 wl_0_127 wl_1_127 bl_0_44 bl_1_44 br_0_44
+ br_1_44 sky130_fd_bd_sram__openram_dp_cell_7003/a_38_n79# vdd_uq1278 gnd sky130_fd_bd_sram__openram_dp_cell_7003/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7014 wl_0_116 wl_1_116 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7025 wl_0_123 wl_1_123 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7047 wl_0_119 wl_1_119 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7036 wl_0_117 wl_1_117 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6302 wl_0_79 wl_1_79 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7058 wl_0_126 wl_1_126 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7069 wl_0_115 wl_1_115 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5601 wl_0_112 wl_1_112 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6324 wl_0_68 wl_1_68 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6313 wl_0_68 wl_1_68 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6346 wl_0_71 wl_1_71 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6335 wl_0_73 wl_1_73 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5634 wl_0_127 wl_1_127 bl_0_23 bl_1_23 br_0_23
+ br_1_23 sky130_fd_bd_sram__openram_dp_cell_5634/a_38_n79# vdd_uq2622 gnd sky130_fd_bd_sram__openram_dp_cell_5634/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5612 wl_0_118 wl_1_118 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5623 wl_0_107 wl_1_107 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6379 wl_0_67 wl_1_67 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6357 wl_0_78 wl_1_78 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6368 wl_0_78 wl_1_78 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5645 wl_0_116 wl_1_116 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5667 wl_0_112 wl_1_112 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4900 wl_0_110 wl_1_110 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4933 wl_0_110 wl_1_110 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4922 wl_0_110 wl_1_110 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5656 wl_0_105 wl_1_105 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4911 wl_0_99 wl_1_99 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4966 wl_0_114 wl_1_114 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4955 wl_0_102 wl_1_102 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4944 wl_0_99 wl_1_99 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5678 wl_0_95 wl_1_95 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5689 wl_0_96 wl_1_96 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4988 wl_0_121 wl_1_121 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4999 wl_0_121 wl_1_121 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4977 wl_0_115 wl_1_115 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7570 wl_0_113 wl_1_113 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7592 wl_0_122 wl_1_122 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7581 wl_0_102 wl_1_102 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6891 wl_0_109 wl_1_109 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6880 wl_0_97 wl_1_97 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4207 wl_0_88 wl_1_88 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4218 wl_0_94 wl_1_94 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3517 wl_0_57 wl_1_57 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3506 wl_0_58 wl_1_58 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4229 wl_0_83 wl_1_83 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2805 wl_0_15 wl_1_15 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3528 wl_0_54 wl_1_54 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3539 wl_0_59 wl_1_59 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2838 wl_0_16 wl_1_16 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2827 wl_0_8 wl_1_8 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2816 wl_0_3 wl_1_3 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2849 wl_0_15 wl_1_15 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6121 wl_0_82 wl_1_82 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6110 wl_0_93 wl_1_93 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6143 wl_0_86 wl_1_86 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6132 wl_0_89 wl_1_89 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6154 wl_0_94 wl_1_94 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5431 wl_0_122 wl_1_122 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5442 wl_0_117 wl_1_117 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5420 wl_0_113 wl_1_113 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6165 wl_0_83 wl_1_83 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6187 wl_0_92 wl_1_92 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6176 wl_0_91 wl_1_91 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5453 wl_0_125 wl_1_125 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5475 wl_0_122 wl_1_122 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5486 wl_0_115 wl_1_115 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5464 wl_0_114 wl_1_114 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4730 wl_0_68 wl_1_68 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6198 wl_0_87 wl_1_87 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4741 wl_0_91 wl_1_91 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5497 wl_0_119 wl_1_119 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4763 wl_0_69 wl_1_69 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4774 wl_0_80 wl_1_80 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4752 wl_0_80 wl_1_80 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4785 wl_0_110 wl_1_110 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4796 wl_0_99 wl_1_99 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8090 wl_0_39 wl_1_39 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_819 wl_0_16 wl_1_16 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_808 wl_0_26 wl_1_26 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4026 wl_0_68 wl_1_68 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4015 wl_0_68 wl_1_68 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4004 wl_0_74 wl_1_74 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3325 wl_0_33 wl_1_33 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3303 wl_0_39 wl_1_39 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3314 wl_0_44 wl_1_44 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4048 wl_0_65 wl_1_65 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4059 wl_0_68 wl_1_68 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4037 wl_0_76 wl_1_76 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2602 wl_0_21 wl_1_21 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2613 wl_0_25 wl_1_25 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3358 wl_0_34 wl_1_34 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3336 wl_0_38 wl_1_38 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3347 wl_0_45 wl_1_45 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2646 wl_0_24 wl_1_24 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2635 wl_0_21 wl_1_21 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2657 wl_0_20 wl_1_20 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1901 wl_0_3 wl_1_3 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2624 wl_0_27 wl_1_27 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1912 wl_0_31 wl_1_31 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3369 wl_0_45 wl_1_45 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2679 wl_0_18 wl_1_18 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2668 wl_0_18 wl_1_18 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1923 wl_0_32 wl_1_32 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1945 wl_0_32 wl_1_32 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1934 wl_0_31 wl_1_31 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1978 wl_0_14 wl_1_14 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1956 wl_0_10 wl_1_10 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1967 wl_0_5 wl_1_5 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1989 wl_0_4 wl_1_4 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5250 wl_0_110 wl_1_110 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5261 wl_0_99 wl_1_99 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5272 wl_0_106 wl_1_106 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5283 wl_0_106 wl_1_106 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5294 wl_0_104 wl_1_104 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4582 wl_0_86 wl_1_86 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4571 wl_0_89 wl_1_89 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4560 wl_0_90 wl_1_90 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3870 wl_0_32 wl_1_32 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3881 wl_0_31 wl_1_31 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4593 wl_0_91 wl_1_91 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3892 wl_0_31 wl_1_31 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1219 wl_0_49 wl_1_49 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1208 wl_0_57 wl_1_57 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_605 wl_0_5 wl_1_5 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_616 wl_0_9 wl_1_9 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_638 wl_0_0 wl_1_0 bl_0_34 bl_1_34 br_0_34 br_1_34
+ sky130_fd_bd_sram__openram_dp_cell_638/a_38_n79# vdd_uq1918 gnd sky130_fd_bd_sram__openram_dp_cell_638/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_627 wl_0_2 wl_1_2 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3100 wl_0_61 wl_1_61 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_649 wl_0_26 wl_1_26 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3111 wl_0_56 wl_1_56 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3133 wl_0_57 wl_1_57 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3122 wl_0_62 wl_1_62 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2432 wl_0_10 wl_1_10 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2421 wl_0_9 wl_1_9 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2410 wl_0_4 wl_1_4 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3166 wl_0_49 wl_1_49 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3144 wl_0_51 wl_1_51 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3155 wl_0_60 wl_1_60 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2454 wl_0_13 wl_1_13 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2443 wl_0_9 wl_1_9 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2465 wl_0_5 wl_1_5 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1720 wl_0_49 wl_1_49 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3188 wl_0_52 wl_1_52 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3177 wl_0_55 wl_1_55 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3199 wl_0_62 wl_1_62 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2476 wl_0_13 wl_1_13 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2487 wl_0_0 wl_1_0 bl_0_5 bl_1_5 br_0_5 br_1_5
+ sky130_fd_bd_sram__openram_dp_cell_2487/a_38_n79# vdd_uq3774 gnd sky130_fd_bd_sram__openram_dp_cell_2487/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2498 wl_0_2 wl_1_2 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1731 wl_0_38 wl_1_38 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1753 wl_0_46 wl_1_46 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1742 wl_0_57 wl_1_57 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1797 wl_0_36 wl_1_36 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1764 wl_0_35 wl_1_35 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1786 wl_0_47 wl_1_47 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1775 wl_0_58 wl_1_58 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5080 wl_0_122 wl_1_122 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5091 wl_0_121 wl_1_121 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4390 wl_0_68 wl_1_68 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6709 wl_0_85 wl_1_85 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1005 wl_0_39 wl_1_39 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1016 wl_0_44 wl_1_44 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1038 wl_0_33 wl_1_33 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1027 wl_0_41 wl_1_41 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1049 wl_0_42 wl_1_42 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7900 wl_0_101 wl_1_101 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7911 wl_0_90 wl_1_90 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7944 wl_0_57 wl_1_57 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7933 wl_0_68 wl_1_68 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7922 wl_0_79 wl_1_79 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7977 wl_0_24 wl_1_24 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7966 wl_0_35 wl_1_35 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7955 wl_0_46 wl_1_46 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7988 wl_0_13 wl_1_13 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7999 wl_0_2 wl_1_2 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_402 wl_0_16 wl_1_16 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_413 wl_0_0 wl_1_0 bl_0_55 bl_1_55 br_0_55 br_1_55
+ sky130_fd_bd_sram__openram_dp_cell_413/a_38_n79# vdd_uq574 gnd sky130_fd_bd_sram__openram_dp_cell_413/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_435 wl_0_19 wl_1_19 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_446 wl_0_8 wl_1_8 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_424 wl_0_30 wl_1_30 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_457 wl_0_16 wl_1_16 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_468 wl_0_3 wl_1_3 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_479 wl_0_4 wl_1_4 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2240 wl_0_21 wl_1_21 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2251 wl_0_23 wl_1_23 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2262 wl_0_21 wl_1_21 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2273 wl_0_25 wl_1_25 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2295 wl_0_24 wl_1_24 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2284 wl_0_18 wl_1_18 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1550 wl_0_52 wl_1_52 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1561 wl_0_54 wl_1_54 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1572 wl_0_62 wl_1_62 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1583 wl_0_51 wl_1_51 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1594 wl_0_55 wl_1_55 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_980 wl_0_39 wl_1_39 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_991 wl_0_43 wl_1_43 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7218 wl_0_105 wl_1_105 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7229 wl_0_105 wl_1_105 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7207 wl_0_98 wl_1_98 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6528 wl_0_82 wl_1_82 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6506 wl_0_84 wl_1_84 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6517 wl_0_93 wl_1_93 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5805 wl_0_100 wl_1_100 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5816 wl_0_89 wl_1_89 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6539 wl_0_89 wl_1_89 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5838 wl_0_67 wl_1_67 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5827 wl_0_78 wl_1_78 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5849 wl_0_96 wl_1_96 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7730 wl_0_120 wl_1_120 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7741 wl_0_109 wl_1_109 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7752 wl_0_98 wl_1_98 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7785 wl_0_65 wl_1_65 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7774 wl_0_76 wl_1_76 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7763 wl_0_87 wl_1_87 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7796 wl_0_96 wl_1_96 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_210 wl_0_25 wl_1_25 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_221 wl_0_30 wl_1_30 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_232 wl_0_22 wl_1_22 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_243 wl_0_19 wl_1_19 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_265 wl_0_17 wl_1_17 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_254 wl_0_25 wl_1_25 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_298 wl_0_22 wl_1_22 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_276 wl_0_23 wl_1_23 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_287 wl_0_25 wl_1_25 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2070 wl_0_1 wl_1_1 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2081 wl_0_1 wl_1_1 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2092 wl_0_6 wl_1_6 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1380 wl_0_36 wl_1_36 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1391 wl_0_42 wl_1_42 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7004 wl_0_126 wl_1_126 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7026 wl_0_122 wl_1_122 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7048 wl_0_118 wl_1_118 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7015 wl_0_115 wl_1_115 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7037 wl_0_116 wl_1_116 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6303 wl_0_80 wl_1_80 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7059 wl_0_125 wl_1_125 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6325 wl_0_67 wl_1_67 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6314 wl_0_67 wl_1_67 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6336 wl_0_72 wl_1_72 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5635 wl_0_126 wl_1_126 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5613 wl_0_117 wl_1_117 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5602 wl_0_111 wl_1_111 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5624 wl_0_106 wl_1_106 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6347 wl_0_70 wl_1_70 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6358 wl_0_77 wl_1_77 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6369 wl_0_77 wl_1_77 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5646 wl_0_115 wl_1_115 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5668 wl_0_111 wl_1_111 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4901 wl_0_109 wl_1_109 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5657 wl_0_104 wl_1_104 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4912 wl_0_98 wl_1_98 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4923 wl_0_98 wl_1_98 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4934 wl_0_109 wl_1_109 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4956 wl_0_101 wl_1_101 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4945 wl_0_98 wl_1_98 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5679 wl_0_96 wl_1_96 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4989 wl_0_122 wl_1_122 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4978 wl_0_114 wl_1_114 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4967 wl_0_113 wl_1_113 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7560 wl_0_123 wl_1_123 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7593 wl_0_121 wl_1_121 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7571 wl_0_112 wl_1_112 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7582 wl_0_101 wl_1_101 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6892 wl_0_110 wl_1_110 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6870 wl_0_105 wl_1_105 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6881 wl_0_99 wl_1_99 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4208 wl_0_87 wl_1_87 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4219 wl_0_93 wl_1_93 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3507 wl_0_57 wl_1_57 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2806 wl_0_13 wl_1_13 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3529 wl_0_53 wl_1_53 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3518 wl_0_62 wl_1_62 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2839 wl_0_15 wl_1_15 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2828 wl_0_7 wl_1_7 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2817 wl_0_2 wl_1_2 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6111 wl_0_92 wl_1_92 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6100 wl_0_92 wl_1_92 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5410 wl_0_126 wl_1_126 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6122 wl_0_81 wl_1_81 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6144 wl_0_85 wl_1_85 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6133 wl_0_88 wl_1_88 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5421 wl_0_127 wl_1_127 bl_0_18 bl_1_18 br_0_18
+ br_1_18 sky130_fd_bd_sram__openram_dp_cell_5421/a_38_n79# vdd_uq2942 gnd sky130_fd_bd_sram__openram_dp_cell_5421/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5432 wl_0_121 wl_1_121 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5443 wl_0_116 wl_1_116 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6166 wl_0_82 wl_1_82 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6177 wl_0_90 wl_1_90 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6188 wl_0_91 wl_1_91 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6155 wl_0_93 wl_1_93 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5454 wl_0_124 wl_1_124 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5476 wl_0_121 wl_1_121 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5465 wl_0_113 wl_1_113 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4731 wl_0_67 wl_1_67 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4720 wl_0_78 wl_1_78 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6199 wl_0_86 wl_1_86 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5487 wl_0_127 wl_1_127 bl_0_19 bl_1_19 br_0_19
+ br_1_19 sky130_fd_bd_sram__openram_dp_cell_5487/a_38_n79# vdd_uq2878 gnd sky130_fd_bd_sram__openram_dp_cell_5487/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5498 wl_0_118 wl_1_118 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4764 wl_0_68 wl_1_68 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4775 wl_0_79 wl_1_79 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4753 wl_0_79 wl_1_79 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4742 wl_0_90 wl_1_90 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4786 wl_0_109 wl_1_109 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4797 wl_0_102 wl_1_102 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8080 wl_0_49 wl_1_49 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8091 wl_0_38 wl_1_38 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7390 wl_0_113 wl_1_113 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_809 wl_0_25 wl_1_25 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4027 wl_0_67 wl_1_67 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4016 wl_0_67 wl_1_67 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4005 wl_0_73 wl_1_73 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3304 wl_0_38 wl_1_38 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3315 wl_0_43 wl_1_43 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4038 wl_0_75 wl_1_75 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4049 wl_0_78 wl_1_78 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2614 wl_0_24 wl_1_24 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2603 wl_0_20 wl_1_20 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3359 wl_0_33 wl_1_33 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3326 wl_0_34 wl_1_34 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3337 wl_0_37 wl_1_37 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3348 wl_0_44 wl_1_44 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2647 wl_0_23 wl_1_23 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2636 wl_0_20 wl_1_20 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1902 wl_0_2 wl_1_2 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2625 wl_0_26 wl_1_26 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2658 wl_0_19 wl_1_19 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2669 wl_0_17 wl_1_17 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1924 wl_0_31 wl_1_31 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1946 wl_0_31 wl_1_31 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1935 wl_0_32 wl_1_32 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1913 wl_0_32 wl_1_32 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1979 wl_0_13 wl_1_13 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1957 wl_0_9 wl_1_9 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1968 wl_0_4 wl_1_4 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5251 wl_0_109 wl_1_109 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5240 wl_0_97 wl_1_97 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5273 wl_0_105 wl_1_105 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5284 wl_0_105 wl_1_105 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5262 wl_0_98 wl_1_98 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4550 wl_0_86 wl_1_86 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5295 wl_0_103 wl_1_103 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4583 wl_0_85 wl_1_85 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4572 wl_0_88 wl_1_88 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4561 wl_0_89 wl_1_89 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3860 wl_0_32 wl_1_32 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3871 wl_0_31 wl_1_31 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4594 wl_0_90 wl_1_90 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3893 wl_0_31 wl_1_31 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3882 wl_0_32 wl_1_32 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1209 wl_0_56 wl_1_56 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_617 wl_0_8 wl_1_8 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_628 wl_0_1 wl_1_1 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_606 wl_0_1 wl_1_1 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_639 wl_0_1 wl_1_1 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3112 wl_0_55 wl_1_55 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3101 wl_0_60 wl_1_60 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3123 wl_0_61 wl_1_61 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3134 wl_0_61 wl_1_61 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2422 wl_0_8 wl_1_8 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2400 wl_0_4 wl_1_4 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2411 wl_0_3 wl_1_3 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3167 wl_0_56 wl_1_56 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3156 wl_0_59 wl_1_59 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3145 wl_0_62 wl_1_62 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2455 wl_0_12 wl_1_12 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2433 wl_0_9 wl_1_9 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2444 wl_0_8 wl_1_8 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1721 wl_0_48 wl_1_48 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3189 wl_0_51 wl_1_51 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3178 wl_0_54 wl_1_54 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1710 wl_0_59 wl_1_59 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2488 wl_0_6 wl_1_6 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2499 wl_0_4 wl_1_4 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2477 wl_0_3 wl_1_3 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2466 wl_0_4 wl_1_4 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1732 wl_0_37 wl_1_37 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1754 wl_0_45 wl_1_45 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1743 wl_0_56 wl_1_56 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1765 wl_0_34 wl_1_34 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1787 wl_0_46 wl_1_46 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1776 wl_0_57 wl_1_57 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1798 wl_0_35 wl_1_35 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5092 wl_0_127 wl_1_127 bl_0_13 bl_1_13 br_0_13
+ br_1_13 sky130_fd_bd_sram__openram_dp_cell_5092/a_38_n79# vdd_uq3262 gnd sky130_fd_bd_sram__openram_dp_cell_5092/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5070 wl_0_127 wl_1_127 bl_0_9 bl_1_9 br_0_9 br_1_9
+ sky130_fd_bd_sram__openram_dp_cell_5070/a_38_n79# vdd_uq3518 gnd sky130_fd_bd_sram__openram_dp_cell_5070/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5081 wl_0_121 wl_1_121 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4380 wl_0_67 wl_1_67 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4391 wl_0_67 wl_1_67 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3690 wl_0_44 wl_1_44 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1006 wl_0_38 wl_1_38 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1028 wl_0_35 wl_1_35 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1017 wl_0_43 wl_1_43 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1039 wl_0_45 wl_1_45 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7901 wl_0_100 wl_1_100 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7934 wl_0_67 wl_1_67 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7923 wl_0_78 wl_1_78 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7912 wl_0_89 wl_1_89 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7978 wl_0_23 wl_1_23 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7967 wl_0_34 wl_1_34 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7956 wl_0_45 wl_1_45 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7945 wl_0_56 wl_1_56 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7989 wl_0_12 wl_1_12 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_403 wl_0_15 wl_1_15 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_414 wl_0_16 wl_1_16 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_436 wl_0_18 wl_1_18 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_447 wl_0_7 wl_1_7 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_425 wl_0_29 wl_1_29 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_458 wl_0_16 wl_1_16 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_469 wl_0_2 wl_1_2 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2230 wl_0_20 wl_1_20 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2274 wl_0_24 wl_1_24 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2252 wl_0_22 wl_1_22 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2241 wl_0_20 wl_1_20 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2263 wl_0_20 wl_1_20 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2296 wl_0_23 wl_1_23 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2285 wl_0_17 wl_1_17 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1551 wl_0_51 wl_1_51 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1562 wl_0_53 wl_1_53 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1540 wl_0_62 wl_1_62 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1584 wl_0_50 wl_1_50 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1595 wl_0_54 wl_1_54 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1573 wl_0_61 wl_1_61 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_970 wl_0_34 wl_1_34 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_981 wl_0_38 wl_1_38 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_992 wl_0_42 wl_1_42 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7219 wl_0_104 wl_1_104 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7208 wl_0_97 wl_1_97 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6507 wl_0_83 wl_1_83 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6518 wl_0_92 wl_1_92 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5806 wl_0_99 wl_1_99 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6529 wl_0_81 wl_1_81 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5817 wl_0_88 wl_1_88 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5839 wl_0_66 wl_1_66 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5828 wl_0_77 wl_1_77 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7731 wl_0_119 wl_1_119 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7742 wl_0_108 wl_1_108 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7753 wl_0_97 wl_1_97 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7720 wl_0_67 wl_1_67 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7786 wl_0_96 wl_1_96 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7775 wl_0_75 wl_1_75 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7764 wl_0_86 wl_1_86 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7797 wl_0_95 wl_1_95 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_200 wl_0_19 wl_1_19 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_211 wl_0_24 wl_1_24 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_222 wl_0_29 wl_1_29 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_233 wl_0_21 wl_1_21 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_244 wl_0_23 wl_1_23 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_255 wl_0_30 wl_1_30 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_277 wl_0_22 wl_1_22 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_288 wl_0_24 wl_1_24 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_266 wl_0_26 wl_1_26 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_299 wl_0_21 wl_1_21 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2060 wl_0_11 wl_1_11 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2071 wl_0_0 wl_1_0 bl_0_18 bl_1_18 br_0_18 br_1_18
+ sky130_fd_bd_sram__openram_dp_cell_2071/a_38_n79# vdd_uq2942 gnd sky130_fd_bd_sram__openram_dp_cell_2071/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2082 wl_0_0 wl_1_0 bl_0_17 bl_1_17 br_0_17 br_1_17
+ sky130_fd_bd_sram__openram_dp_cell_2082/a_38_n79# vdd_uq3006 gnd sky130_fd_bd_sram__openram_dp_cell_2082/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2093 wl_0_5 wl_1_5 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1370 wl_0_46 wl_1_46 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1381 wl_0_35 wl_1_35 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1392 wl_0_41 wl_1_41 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7005 wl_0_125 wl_1_125 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7027 wl_0_121 wl_1_121 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7038 wl_0_115 wl_1_115 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7016 wl_0_114 wl_1_114 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7049 wl_0_117 wl_1_117 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6326 wl_0_66 wl_1_66 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6315 wl_0_66 wl_1_66 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6337 wl_0_71 wl_1_71 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6304 wl_0_79 wl_1_79 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5603 wl_0_127 wl_1_127 bl_0_24 bl_1_24 br_0_24
+ br_1_24 sky130_fd_bd_sram__openram_dp_cell_5603/a_38_n79# vdd_uq2558 gnd sky130_fd_bd_sram__openram_dp_cell_5603/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5614 wl_0_116 wl_1_116 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5625 wl_0_105 wl_1_105 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6348 wl_0_69 wl_1_69 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6359 wl_0_76 wl_1_76 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5636 wl_0_125 wl_1_125 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5647 wl_0_114 wl_1_114 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4902 wl_0_108 wl_1_108 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5658 wl_0_103 wl_1_103 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4913 wl_0_97 wl_1_97 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4924 wl_0_97 wl_1_97 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5669 wl_0_112 wl_1_112 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4935 wl_0_108 wl_1_108 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4957 wl_0_100 wl_1_100 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4946 wl_0_97 wl_1_97 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4968 wl_0_118 wl_1_118 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4979 wl_0_113 wl_1_113 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7561 wl_0_122 wl_1_122 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7550 wl_0_112 wl_1_112 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7594 wl_0_120 wl_1_120 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7572 wl_0_111 wl_1_111 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7583 wl_0_100 wl_1_100 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6893 wl_0_109 wl_1_109 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6871 wl_0_104 wl_1_104 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6860 wl_0_100 wl_1_100 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6882 wl_0_98 wl_1_98 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_90 wl_0_0 wl_1_0 bl_0_60 bl_1_60 br_0_60 br_1_60
+ sky130_fd_bd_sram__openram_dp_cell_90/a_38_n79# vdd_uq254 gnd sky130_fd_bd_sram__openram_dp_cell_90/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4209 wl_0_86 wl_1_86 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3508 wl_0_56 wl_1_56 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3519 wl_0_61 wl_1_61 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2807 wl_0_12 wl_1_12 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2829 wl_0_6 wl_1_6 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2818 wl_0_1 wl_1_1 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6112 wl_0_91 wl_1_91 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6101 wl_0_91 wl_1_91 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5400 wl_0_97 wl_1_97 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6123 wl_0_82 wl_1_82 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6145 wl_0_84 wl_1_84 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6134 wl_0_87 wl_1_87 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5433 wl_0_126 wl_1_126 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5411 wl_0_125 wl_1_125 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5422 wl_0_114 wl_1_114 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6167 wl_0_81 wl_1_81 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6178 wl_0_89 wl_1_89 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6156 wl_0_92 wl_1_92 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5455 wl_0_123 wl_1_123 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5477 wl_0_120 wl_1_120 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5466 wl_0_118 wl_1_118 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5444 wl_0_115 wl_1_115 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4721 wl_0_77 wl_1_77 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4732 wl_0_80 wl_1_80 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4710 wl_0_86 wl_1_86 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6189 wl_0_90 wl_1_90 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5499 wl_0_127 wl_1_127 bl_0_30 bl_1_30 br_0_30
+ br_1_30 sky130_fd_bd_sram__openram_dp_cell_5499/a_38_n79# vdd_uq2174 gnd sky130_fd_bd_sram__openram_dp_cell_5499/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5488 wl_0_116 wl_1_116 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4765 wl_0_67 wl_1_67 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4754 wl_0_78 wl_1_78 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4743 wl_0_89 wl_1_89 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4776 wl_0_109 wl_1_109 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4787 wl_0_108 wl_1_108 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4798 wl_0_101 wl_1_101 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8081 wl_0_48 wl_1_48 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8070 wl_0_59 wl_1_59 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8092 wl_0_37 wl_1_37 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7380 wl_0_121 wl_1_121 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7391 wl_0_117 wl_1_117 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6690 wl_0_80 wl_1_80 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4017 wl_0_66 wl_1_66 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4006 wl_0_72 wl_1_72 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3305 wl_0_37 wl_1_37 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3316 wl_0_42 wl_1_42 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4028 wl_0_66 wl_1_66 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4039 wl_0_74 wl_1_74 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2604 wl_0_19 wl_1_19 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3327 wl_0_33 wl_1_33 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3349 wl_0_43 wl_1_43 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3338 wl_0_46 wl_1_46 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2648 wl_0_22 wl_1_22 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1903 wl_0_1 wl_1_1 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2637 wl_0_25 wl_1_25 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2626 wl_0_30 wl_1_30 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2615 wl_0_30 wl_1_30 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2659 wl_0_18 wl_1_18 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1925 wl_0_32 wl_1_32 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1936 wl_0_31 wl_1_31 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1914 wl_0_31 wl_1_31 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1958 wl_0_8 wl_1_8 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1969 wl_0_3 wl_1_3 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1947 wl_0_32 wl_1_32 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5252 wl_0_108 wl_1_108 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5230 wl_0_107 wl_1_107 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5241 wl_0_101 wl_1_101 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5274 wl_0_104 wl_1_104 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5285 wl_0_104 wl_1_104 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5263 wl_0_97 wl_1_97 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4540 wl_0_90 wl_1_90 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5296 wl_0_102 wl_1_102 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4551 wl_0_85 wl_1_85 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4573 wl_0_87 wl_1_87 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4562 wl_0_88 wl_1_88 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3850 wl_0_7 wl_1_7 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3861 wl_0_31 wl_1_31 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3872 wl_0_32 wl_1_32 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4595 wl_0_89 wl_1_89 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4584 wl_0_90 wl_1_90 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3894 wl_0_32 wl_1_32 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3883 wl_0_31 wl_1_31 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_618 wl_0_7 wl_1_7 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_629 wl_0_0 wl_1_0 bl_0_38 bl_1_38 br_0_38 br_1_38
+ sky130_fd_bd_sram__openram_dp_cell_629/a_38_n79# vdd_uq1662 gnd sky130_fd_bd_sram__openram_dp_cell_629/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_607 wl_0_0 wl_1_0 bl_0_37 bl_1_37 br_0_37 br_1_37
+ sky130_fd_bd_sram__openram_dp_cell_607/a_38_n79# vdd_uq1726 gnd sky130_fd_bd_sram__openram_dp_cell_607/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3113 wl_0_54 wl_1_54 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3124 wl_0_60 wl_1_60 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3102 wl_0_59 wl_1_59 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2423 wl_0_14 wl_1_14 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2412 wl_0_2 wl_1_2 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2401 wl_0_3 wl_1_3 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3146 wl_0_50 wl_1_50 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3157 wl_0_58 wl_1_58 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3135 wl_0_60 wl_1_60 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2456 wl_0_11 wl_1_11 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2434 wl_0_8 wl_1_8 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2445 wl_0_7 wl_1_7 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1700 wl_0_47 wl_1_47 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3179 wl_0_53 wl_1_53 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3168 wl_0_55 wl_1_55 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1711 wl_0_58 wl_1_58 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2478 wl_0_2 wl_1_2 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2467 wl_0_3 wl_1_3 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2489 wl_0_5 wl_1_5 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1733 wl_0_36 wl_1_36 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1722 wl_0_47 wl_1_47 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1744 wl_0_55 wl_1_55 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1766 wl_0_33 wl_1_33 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1755 wl_0_44 wl_1_44 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1788 wl_0_45 wl_1_45 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1777 wl_0_56 wl_1_56 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1799 wl_0_34 wl_1_34 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5060 wl_0_120 wl_1_120 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5093 wl_0_126 wl_1_126 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5071 wl_0_126 wl_1_126 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5082 wl_0_120 wl_1_120 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4392 wl_0_66 wl_1_66 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4370 wl_0_73 wl_1_73 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4381 wl_0_77 wl_1_77 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3680 wl_0_54 wl_1_54 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3691 wl_0_43 wl_1_43 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2990 wl_0_34 wl_1_34 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1007 wl_0_37 wl_1_37 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1029 wl_0_34 wl_1_34 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1018 wl_0_42 wl_1_42 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7902 wl_0_99 wl_1_99 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7935 wl_0_66 wl_1_66 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7924 wl_0_77 wl_1_77 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7913 wl_0_88 wl_1_88 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7968 wl_0_33 wl_1_33 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7957 wl_0_44 wl_1_44 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7946 wl_0_55 wl_1_55 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7979 wl_0_22 wl_1_22 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_404 wl_0_7 wl_1_7 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_437 wl_0_17 wl_1_17 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_415 wl_0_15 wl_1_15 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_426 wl_0_28 wl_1_28 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_459 wl_0_15 wl_1_15 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_448 wl_0_6 wl_1_6 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2231 wl_0_19 wl_1_19 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2220 wl_0_30 wl_1_30 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2242 wl_0_19 wl_1_19 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2264 wl_0_19 wl_1_19 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2253 wl_0_30 wl_1_30 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2275 wl_0_23 wl_1_23 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2297 wl_0_22 wl_1_22 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2286 wl_0_17 wl_1_17 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1552 wl_0_50 wl_1_50 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1563 wl_0_52 wl_1_52 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1530 wl_0_57 wl_1_57 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1541 wl_0_61 wl_1_61 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1596 wl_0_53 wl_1_53 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1585 wl_0_54 wl_1_54 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1574 wl_0_60 wl_1_60 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_960 wl_0_44 wl_1_44 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_971 wl_0_33 wl_1_33 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_982 wl_0_34 wl_1_34 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_993 wl_0_41 wl_1_41 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7209 wl_0_97 wl_1_97 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6508 wl_0_90 wl_1_90 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6519 wl_0_91 wl_1_91 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5807 wl_0_98 wl_1_98 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5829 wl_0_76 wl_1_76 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5818 wl_0_87 wl_1_87 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7710 wl_0_77 wl_1_77 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7732 wl_0_118 wl_1_118 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7743 wl_0_107 wl_1_107 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7721 wl_0_66 wl_1_66 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7754 wl_0_96 wl_1_96 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7776 wl_0_74 wl_1_74 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7765 wl_0_85 wl_1_85 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7787 wl_0_95 wl_1_95 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7798 wl_0_96 wl_1_96 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_201 wl_0_18 wl_1_18 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_212 wl_0_23 wl_1_23 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_245 wl_0_22 wl_1_22 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_234 wl_0_20 wl_1_20 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_223 wl_0_28 wl_1_28 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_256 wl_0_29 wl_1_29 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_278 wl_0_21 wl_1_21 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_289 wl_0_23 wl_1_23 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_267 wl_0_25 wl_1_25 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2050 wl_0_13 wl_1_13 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2061 wl_0_10 wl_1_10 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2072 wl_0_10 wl_1_10 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2083 wl_0_10 wl_1_10 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2094 wl_0_4 wl_1_4 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1360 wl_0_43 wl_1_43 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1371 wl_0_45 wl_1_45 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1382 wl_0_34 wl_1_34 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1393 wl_0_40 wl_1_40 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_790 wl_0_21 wl_1_21 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7039 wl_0_127 wl_1_127 bl_0_42 bl_1_42 br_0_42
+ br_1_42 sky130_fd_bd_sram__openram_dp_cell_7039/a_38_n79# vdd_uq1406 gnd sky130_fd_bd_sram__openram_dp_cell_7039/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7006 wl_0_124 wl_1_124 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7028 wl_0_120 wl_1_120 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7017 wl_0_113 wl_1_113 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6327 wl_0_65 wl_1_65 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6316 wl_0_65 wl_1_65 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6305 wl_0_80 wl_1_80 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5604 wl_0_126 wl_1_126 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5615 wl_0_115 wl_1_115 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5626 wl_0_104 wl_1_104 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6349 wl_0_68 wl_1_68 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6338 wl_0_70 wl_1_70 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5637 wl_0_124 wl_1_124 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5648 wl_0_113 wl_1_113 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4914 wl_0_110 wl_1_110 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4903 wl_0_107 wl_1_107 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5659 wl_0_102 wl_1_102 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4947 wl_0_108 wl_1_108 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4936 wl_0_107 wl_1_107 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4925 wl_0_102 wl_1_102 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4969 wl_0_118 wl_1_118 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4958 wl_0_117 wl_1_117 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7540 wl_0_112 wl_1_112 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7551 wl_0_111 wl_1_111 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7562 wl_0_121 wl_1_121 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7595 wl_0_119 wl_1_119 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7573 wl_0_110 wl_1_110 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6850 wl_0_105 wl_1_105 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7584 wl_0_99 wl_1_99 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6883 wl_0_108 wl_1_108 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6861 wl_0_99 wl_1_99 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6872 wl_0_97 wl_1_97 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6894 wl_0_106 wl_1_106 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_80 wl_0_10 wl_1_10 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_91 wl_0_8 wl_1_8 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1190 wl_0_55 wl_1_55 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3509 wl_0_55 wl_1_55 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2808 wl_0_11 wl_1_11 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2819 wl_0_0 wl_1_0 bl_0_7 bl_1_7 br_0_7 br_1_7
+ sky130_fd_bd_sram__openram_dp_cell_2819/a_38_n79# vdd_uq3646 gnd sky130_fd_bd_sram__openram_dp_cell_2819/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6102 wl_0_89 wl_1_89 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5401 wl_0_110 wl_1_110 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6135 wl_0_86 wl_1_86 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6113 wl_0_90 wl_1_90 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6124 wl_0_94 wl_1_94 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5434 wl_0_125 wl_1_125 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5412 wl_0_124 wl_1_124 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5423 wl_0_113 wl_1_113 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6146 wl_0_83 wl_1_83 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6179 wl_0_88 wl_1_88 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6157 wl_0_91 wl_1_91 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6168 wl_0_93 wl_1_93 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5456 wl_0_122 wl_1_122 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5467 wl_0_117 wl_1_117 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5445 wl_0_114 wl_1_114 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4722 wl_0_76 wl_1_76 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4700 wl_0_80 wl_1_80 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4711 wl_0_85 wl_1_85 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5478 wl_0_119 wl_1_119 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5489 wl_0_115 wl_1_115 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4766 wl_0_66 wl_1_66 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4755 wl_0_77 wl_1_77 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4733 wl_0_79 wl_1_79 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4744 wl_0_88 wl_1_88 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4788 wl_0_107 wl_1_107 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4777 wl_0_108 wl_1_108 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4799 wl_0_100 wl_1_100 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8071 wl_0_58 wl_1_58 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8060 wl_0_69 wl_1_69 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8093 wl_0_36 wl_1_36 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8082 wl_0_47 wl_1_47 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7381 wl_0_122 wl_1_122 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7392 wl_0_116 wl_1_116 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7370 wl_0_113 wl_1_113 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6680 wl_0_78 wl_1_78 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6691 wl_0_79 wl_1_79 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5990 wl_0_68 wl_1_68 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4018 wl_0_65 wl_1_65 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4007 wl_0_71 wl_1_71 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3306 wl_0_36 wl_1_36 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4029 wl_0_78 wl_1_78 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2605 wl_0_30 wl_1_30 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3317 wl_0_41 wl_1_41 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3339 wl_0_45 wl_1_45 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3328 wl_0_46 wl_1_46 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2638 wl_0_24 wl_1_24 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2627 wl_0_29 wl_1_29 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2616 wl_0_29 wl_1_29 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2649 wl_0_21 wl_1_21 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1904 wl_0_0 wl_1_0 bl_0_47 bl_1_47 br_0_47 br_1_47
+ sky130_fd_bd_sram__openram_dp_cell_1904/a_38_n79# vdd_uq1086 gnd sky130_fd_bd_sram__openram_dp_cell_1904/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1915 wl_0_32 wl_1_32 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1926 wl_0_31 wl_1_31 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1937 wl_0_32 wl_1_32 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1959 wl_0_7 wl_1_7 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1948 wl_0_31 wl_1_31 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5220 wl_0_117 wl_1_117 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5231 wl_0_106 wl_1_106 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5242 wl_0_100 wl_1_100 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5253 wl_0_107 wl_1_107 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5275 wl_0_103 wl_1_103 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5264 wl_0_97 wl_1_97 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4530 wl_0_88 wl_1_88 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5297 wl_0_110 wl_1_110 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5286 wl_0_103 wl_1_103 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4552 wl_0_84 wl_1_84 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4574 wl_0_86 wl_1_86 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4563 wl_0_87 wl_1_87 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4541 wl_0_89 wl_1_89 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3840 wl_0_17 wl_1_17 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3851 wl_0_6 wl_1_6 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3862 wl_0_32 wl_1_32 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4596 wl_0_88 wl_1_88 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4585 wl_0_89 wl_1_89 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3884 wl_0_32 wl_1_32 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3895 wl_0_31 wl_1_31 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3873 wl_0_31 wl_1_31 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_619 wl_0_6 wl_1_6 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_608 wl_0_3 wl_1_3 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3114 wl_0_53 wl_1_53 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3103 wl_0_58 wl_1_58 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3125 wl_0_59 wl_1_59 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2413 wl_0_1 wl_1_1 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2402 wl_0_2 wl_1_2 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3147 wl_0_49 wl_1_49 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3158 wl_0_57 wl_1_57 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3136 wl_0_59 wl_1_59 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2424 wl_0_13 wl_1_13 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2435 wl_0_7 wl_1_7 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2446 wl_0_6 wl_1_6 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1701 wl_0_48 wl_1_48 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3169 wl_0_54 wl_1_54 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1712 wl_0_57 wl_1_57 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2457 wl_0_10 wl_1_10 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2479 wl_0_1 wl_1_1 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2468 wl_0_2 wl_1_2 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1734 wl_0_35 wl_1_35 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1723 wl_0_46 wl_1_46 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1745 wl_0_54 wl_1_54 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1756 wl_0_43 wl_1_43 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1767 wl_0_48 wl_1_48 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1778 wl_0_55 wl_1_55 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1789 wl_0_44 wl_1_44 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5050 wl_0_115 wl_1_115 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5094 wl_0_125 wl_1_125 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5072 wl_0_125 wl_1_125 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5083 wl_0_119 wl_1_119 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5061 wl_0_120 wl_1_120 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4371 wl_0_72 wl_1_72 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4360 wl_0_74 wl_1_74 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4382 wl_0_76 wl_1_76 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3670 wl_0_48 wl_1_48 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4393 wl_0_65 wl_1_65 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3692 wl_0_42 wl_1_42 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3681 wl_0_53 wl_1_53 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2991 wl_0_33 wl_1_33 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2980 wl_0_44 wl_1_44 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1008 wl_0_36 wl_1_36 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1019 wl_0_41 wl_1_41 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7903 wl_0_98 wl_1_98 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7925 wl_0_76 wl_1_76 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7914 wl_0_87 wl_1_87 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7969 wl_0_32 wl_1_32 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7958 wl_0_43 wl_1_43 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7947 wl_0_54 wl_1_54 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7936 wl_0_65 wl_1_65 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_405 wl_0_6 wl_1_6 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_438 wl_0_16 wl_1_16 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_416 wl_0_16 wl_1_16 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_427 wl_0_27 wl_1_27 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_449 wl_0_5 wl_1_5 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2210 wl_0_19 wl_1_19 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2221 wl_0_29 wl_1_29 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2243 wl_0_18 wl_1_18 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2265 wl_0_18 wl_1_18 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2232 wl_0_18 wl_1_18 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2254 wl_0_29 wl_1_29 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1520 wl_0_49 wl_1_49 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2276 wl_0_22 wl_1_22 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2298 wl_0_21 wl_1_21 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2287 wl_0_30 wl_1_30 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1553 wl_0_49 wl_1_49 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1531 wl_0_56 wl_1_56 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1542 wl_0_60 wl_1_60 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1564 wl_0_51 wl_1_51 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1586 wl_0_53 wl_1_53 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1575 wl_0_59 wl_1_59 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1597 wl_0_52 wl_1_52 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_950 wl_0_42 wl_1_42 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_994 wl_0_40 wl_1_40 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_972 wl_0_39 wl_1_39 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_983 wl_0_44 wl_1_44 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_961 wl_0_43 wl_1_43 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4190 wl_0_86 wl_1_86 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6509 wl_0_89 wl_1_89 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5808 wl_0_97 wl_1_97 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5819 wl_0_86 wl_1_86 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7700 wl_0_87 wl_1_87 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7733 wl_0_117 wl_1_117 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7744 wl_0_106 wl_1_106 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7722 wl_0_65 wl_1_65 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7711 wl_0_76 wl_1_76 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7755 wl_0_95 wl_1_95 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7777 wl_0_73 wl_1_73 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7766 wl_0_84 wl_1_84 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7788 wl_0_96 wl_1_96 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7799 wl_0_95 wl_1_95 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_213 wl_0_22 wl_1_22 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_202 wl_0_17 wl_1_17 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_246 wl_0_21 wl_1_21 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_235 wl_0_19 wl_1_19 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_224 wl_0_27 wl_1_27 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_257 wl_0_28 wl_1_28 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_279 wl_0_29 wl_1_29 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_268 wl_0_30 wl_1_30 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2051 wl_0_12 wl_1_12 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2062 wl_0_9 wl_1_9 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2073 wl_0_9 wl_1_9 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2040 wl_0_0 wl_1_0 bl_0_25 bl_1_25 br_0_25 br_1_25
+ sky130_fd_bd_sram__openram_dp_cell_2040/a_38_n79# vdd_uq2494 gnd sky130_fd_bd_sram__openram_dp_cell_2040/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2084 wl_0_9 wl_1_9 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2095 wl_0_3 wl_1_3 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1350 wl_0_33 wl_1_33 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1361 wl_0_42 wl_1_42 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1383 wl_0_33 wl_1_33 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1394 wl_0_39 wl_1_39 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1372 wl_0_44 wl_1_44 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_780 wl_0_20 wl_1_20 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_791 wl_0_20 wl_1_20 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7007 wl_0_123 wl_1_123 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7029 wl_0_119 wl_1_119 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7018 wl_0_120 wl_1_120 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6317 wl_0_75 wl_1_75 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6328 wl_0_77 wl_1_77 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6306 wl_0_79 wl_1_79 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5605 wl_0_125 wl_1_125 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5616 wl_0_114 wl_1_114 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6339 wl_0_78 wl_1_78 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5638 wl_0_123 wl_1_123 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5649 wl_0_112 wl_1_112 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4915 wl_0_109 wl_1_109 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4904 wl_0_106 wl_1_106 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5627 wl_0_103 wl_1_103 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4948 wl_0_107 wl_1_107 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4937 wl_0_106 wl_1_106 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4926 wl_0_104 wl_1_104 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4959 wl_0_116 wl_1_116 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7530 wl_0_120 wl_1_120 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7541 wl_0_111 wl_1_111 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7552 wl_0_112 wl_1_112 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7563 wl_0_120 wl_1_120 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7574 wl_0_109 wl_1_109 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7585 wl_0_98 wl_1_98 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6840 wl_0_98 wl_1_98 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7596 wl_0_118 wl_1_118 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6851 wl_0_104 wl_1_104 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6873 wl_0_103 wl_1_103 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6884 wl_0_102 wl_1_102 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6862 wl_0_98 wl_1_98 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6895 wl_0_110 wl_1_110 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_70 wl_0_14 wl_1_14 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_81 wl_0_9 wl_1_9 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_92 wl_0_7 wl_1_7 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1180 wl_0_49 wl_1_49 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1191 wl_0_54 wl_1_54 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2809 wl_0_10 wl_1_10 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6103 wl_0_88 wl_1_88 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6136 wl_0_85 wl_1_85 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6114 wl_0_89 wl_1_89 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6125 wl_0_90 wl_1_90 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5424 wl_0_126 wl_1_126 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5413 wl_0_123 wl_1_123 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5402 wl_0_109 wl_1_109 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6147 wl_0_82 wl_1_82 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6158 wl_0_90 wl_1_90 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6169 wl_0_92 wl_1_92 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5468 wl_0_127 wl_1_127 bl_0_20 bl_1_20 br_0_20
+ br_1_20 sky130_fd_bd_sram__openram_dp_cell_5468/a_38_n79# vdd_uq2814 gnd sky130_fd_bd_sram__openram_dp_cell_5468/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5435 wl_0_124 wl_1_124 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5457 wl_0_121 wl_1_121 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5446 wl_0_113 wl_1_113 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4723 wl_0_75 wl_1_75 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4701 wl_0_79 wl_1_79 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4712 wl_0_84 wl_1_84 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5479 wl_0_118 wl_1_118 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4756 wl_0_76 wl_1_76 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4734 wl_0_80 wl_1_80 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4745 wl_0_87 wl_1_87 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4778 wl_0_107 wl_1_107 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4789 wl_0_106 wl_1_106 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4767 wl_0_65 wl_1_65 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8072 wl_0_57 wl_1_57 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8061 wl_0_68 wl_1_68 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8050 wl_0_79 wl_1_79 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7360 wl_0_127 wl_1_127 bl_0_50 bl_1_50 br_0_50
+ br_1_50 sky130_fd_bd_sram__openram_dp_cell_7360/a_38_n79# vdd_uq894 gnd sky130_fd_bd_sram__openram_dp_cell_7360/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8094 wl_0_35 wl_1_35 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8083 wl_0_46 wl_1_46 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7393 wl_0_127 wl_1_127 bl_0_53 bl_1_53 br_0_53
+ br_1_53 sky130_fd_bd_sram__openram_dp_cell_7393/a_38_n79# vdd_uq702 gnd sky130_fd_bd_sram__openram_dp_cell_7393/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7382 wl_0_121 wl_1_121 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7371 wl_0_120 wl_1_120 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6692 wl_0_68 wl_1_68 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6681 wl_0_77 wl_1_77 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6670 wl_0_88 wl_1_88 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5980 wl_0_71 wl_1_71 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5991 wl_0_74 wl_1_74 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4008 wl_0_70 wl_1_70 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3307 wl_0_35 wl_1_35 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4019 wl_0_69 wl_1_69 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3318 wl_0_40 wl_1_40 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3329 wl_0_45 wl_1_45 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2639 wl_0_23 wl_1_23 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2628 wl_0_28 wl_1_28 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2617 wl_0_28 wl_1_28 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2606 wl_0_29 wl_1_29 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1916 wl_0_31 wl_1_31 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1927 wl_0_32 wl_1_32 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1905 wl_0_32 wl_1_32 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1949 wl_0_32 wl_1_32 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1938 wl_0_31 wl_1_31 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5210 wl_0_127 wl_1_127 bl_0_7 bl_1_7 br_0_7 br_1_7
+ sky130_fd_bd_sram__openram_dp_cell_5210/a_38_n79# vdd_uq3646 gnd sky130_fd_bd_sram__openram_dp_cell_5210/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5221 wl_0_116 wl_1_116 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5232 wl_0_105 wl_1_105 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5243 wl_0_99 wl_1_99 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5265 wl_0_110 wl_1_110 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5254 wl_0_106 wl_1_106 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5276 wl_0_102 wl_1_102 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4531 wl_0_87 wl_1_87 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4520 wl_0_94 wl_1_94 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5298 wl_0_109 wl_1_109 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5287 wl_0_102 wl_1_102 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4553 wl_0_83 wl_1_83 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4564 wl_0_86 wl_1_86 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4542 wl_0_94 wl_1_94 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3841 wl_0_16 wl_1_16 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3852 wl_0_5 wl_1_5 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3830 wl_0_27 wl_1_27 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3863 wl_0_31 wl_1_31 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4575 wl_0_85 wl_1_85 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4597 wl_0_87 wl_1_87 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4586 wl_0_88 wl_1_88 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3885 wl_0_31 wl_1_31 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3896 wl_0_32 wl_1_32 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3874 wl_0_32 wl_1_32 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7190 wl_0_100 wl_1_100 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_609 wl_0_2 wl_1_2 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3104 wl_0_57 wl_1_57 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3115 wl_0_62 wl_1_62 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2414 wl_0_0 wl_1_0 bl_0_14 bl_1_14 br_0_14 br_1_14
+ sky130_fd_bd_sram__openram_dp_cell_2414/a_38_n79# vdd_uq3198 gnd sky130_fd_bd_sram__openram_dp_cell_2414/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2403 wl_0_1 wl_1_1 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3126 wl_0_58 wl_1_58 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3137 wl_0_58 wl_1_58 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3148 wl_0_62 wl_1_62 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2425 wl_0_12 wl_1_12 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2436 wl_0_6 wl_1_6 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2447 wl_0_5 wl_1_5 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1702 wl_0_47 wl_1_47 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3159 wl_0_56 wl_1_56 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2458 wl_0_9 wl_1_9 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2469 wl_0_1 wl_1_1 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1735 wl_0_34 wl_1_34 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1724 wl_0_45 wl_1_45 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1713 wl_0_56 wl_1_56 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1757 wl_0_42 wl_1_42 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1768 wl_0_47 wl_1_47 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1746 wl_0_53 wl_1_53 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1779 wl_0_54 wl_1_54 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5040 wl_0_125 wl_1_125 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5051 wl_0_114 wl_1_114 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5073 wl_0_124 wl_1_124 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5062 wl_0_119 wl_1_119 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5084 wl_0_118 wl_1_118 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5095 wl_0_124 wl_1_124 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4372 wl_0_71 wl_1_71 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4361 wl_0_73 wl_1_73 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4350 wl_0_74 wl_1_74 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3660 wl_0_48 wl_1_48 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3671 wl_0_47 wl_1_47 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4394 wl_0_66 wl_1_66 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4383 wl_0_75 wl_1_75 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3693 wl_0_41 wl_1_41 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3682 wl_0_52 wl_1_52 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2970 wl_0_37 wl_1_37 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2981 wl_0_43 wl_1_43 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2992 wl_0_45 wl_1_45 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1009 wl_0_35 wl_1_35 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7904 wl_0_97 wl_1_97 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7926 wl_0_75 wl_1_75 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7915 wl_0_86 wl_1_86 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7959 wl_0_42 wl_1_42 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7948 wl_0_53 wl_1_53 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7937 wl_0_64 wl_1_64 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_417 wl_0_15 wl_1_15 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_406 wl_0_5 wl_1_5 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_428 wl_0_26 wl_1_26 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_439 wl_0_15 wl_1_15 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2211 wl_0_18 wl_1_18 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2222 wl_0_28 wl_1_28 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2200 wl_0_29 wl_1_29 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2233 wl_0_17 wl_1_17 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2255 wl_0_28 wl_1_28 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2244 wl_0_30 wl_1_30 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1510 wl_0_58 wl_1_58 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2277 wl_0_21 wl_1_21 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2266 wl_0_17 wl_1_17 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2288 wl_0_29 wl_1_29 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1532 wl_0_55 wl_1_55 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1543 wl_0_59 wl_1_59 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1521 wl_0_61 wl_1_61 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1554 wl_0_61 wl_1_61 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2299 wl_0_20 wl_1_20 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1565 wl_0_50 wl_1_50 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1576 wl_0_58 wl_1_58 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1587 wl_0_62 wl_1_62 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1598 wl_0_51 wl_1_51 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_940 wl_0_38 wl_1_38 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_951 wl_0_41 wl_1_41 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_984 wl_0_35 wl_1_35 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_973 wl_0_38 wl_1_38 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_962 wl_0_42 wl_1_42 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4191 wl_0_85 wl_1_85 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4180 wl_0_94 wl_1_94 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_995 wl_0_39 wl_1_39 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3490 wl_0_56 wl_1_56 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5809 wl_0_96 wl_1_96 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7701 wl_0_86 wl_1_86 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7723 wl_0_127 wl_1_127 bl_0_47 bl_1_47 br_0_47
+ br_1_47 sky130_fd_bd_sram__openram_dp_cell_7723/a_38_n79# vdd_uq1086 gnd sky130_fd_bd_sram__openram_dp_cell_7723/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7734 wl_0_116 wl_1_116 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7712 wl_0_75 wl_1_75 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7745 wl_0_105 wl_1_105 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7767 wl_0_83 wl_1_83 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7756 wl_0_94 wl_1_94 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7789 wl_0_95 wl_1_95 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7778 wl_0_72 wl_1_72 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_203 wl_0_20 wl_1_20 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_214 wl_0_21 wl_1_21 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_247 wl_0_20 wl_1_20 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_236 wl_0_18 wl_1_18 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_225 wl_0_26 wl_1_26 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_258 wl_0_27 wl_1_27 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_269 wl_0_30 wl_1_30 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2030 wl_0_4 wl_1_4 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2052 wl_0_11 wl_1_11 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2063 wl_0_8 wl_1_8 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2041 wl_0_6 wl_1_6 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2074 wl_0_8 wl_1_8 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2096 wl_0_2 wl_1_2 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2085 wl_0_5 wl_1_5 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1351 wl_0_38 wl_1_38 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1340 wl_0_40 wl_1_40 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1362 wl_0_41 wl_1_41 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1395 wl_0_38 wl_1_38 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1384 wl_0_39 wl_1_39 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1373 wl_0_43 wl_1_43 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_770 wl_0_20 wl_1_20 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_792 wl_0_19 wl_1_19 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_781 wl_0_30 wl_1_30 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7008 wl_0_122 wl_1_122 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7019 wl_0_119 wl_1_119 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6318 wl_0_74 wl_1_74 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6307 wl_0_80 wl_1_80 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5606 wl_0_124 wl_1_124 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5617 wl_0_113 wl_1_113 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6329 wl_0_76 wl_1_76 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5639 wl_0_122 wl_1_122 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4905 wl_0_105 wl_1_105 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5628 wl_0_102 wl_1_102 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4938 wl_0_105 wl_1_105 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4916 wl_0_105 wl_1_105 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4927 wl_0_103 wl_1_103 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4949 wl_0_108 wl_1_108 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7531 wl_0_119 wl_1_119 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7520 wl_0_115 wl_1_115 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7542 wl_0_112 wl_1_112 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7564 wl_0_119 wl_1_119 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7553 wl_0_111 wl_1_111 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7575 wl_0_108 wl_1_108 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6830 wl_0_99 wl_1_99 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7586 wl_0_97 wl_1_97 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6841 wl_0_97 wl_1_97 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7597 wl_0_117 wl_1_117 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6863 wl_0_110 wl_1_110 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6874 wl_0_103 wl_1_103 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6852 wl_0_100 wl_1_100 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6885 wl_0_110 wl_1_110 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6896 wl_0_109 wl_1_109 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_71 wl_0_13 wl_1_13 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_60 wl_0_9 wl_1_9 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_82 wl_0_8 wl_1_8 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_93 wl_0_6 wl_1_6 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1170 wl_0_58 wl_1_58 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1192 wl_0_53 wl_1_53 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1181 wl_0_57 wl_1_57 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6115 wl_0_88 wl_1_88 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6104 wl_0_87 wl_1_87 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6126 wl_0_89 wl_1_89 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5425 wl_0_125 wl_1_125 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5414 wl_0_117 wl_1_117 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5403 wl_0_100 wl_1_100 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6148 wl_0_81 wl_1_81 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6137 wl_0_84 wl_1_84 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6159 wl_0_89 wl_1_89 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5436 wl_0_123 wl_1_123 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5458 wl_0_120 wl_1_120 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5447 wl_0_120 wl_1_120 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4713 wl_0_83 wl_1_83 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4702 wl_0_94 wl_1_94 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5469 wl_0_118 wl_1_118 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4724 wl_0_74 wl_1_74 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4757 wl_0_75 wl_1_75 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4735 wl_0_79 wl_1_79 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4746 wl_0_86 wl_1_86 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4779 wl_0_106 wl_1_106 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4768 wl_0_80 wl_1_80 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8062 wl_0_67 wl_1_67 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8051 wl_0_78 wl_1_78 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8040 wl_0_89 wl_1_89 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7350 wl_0_120 wl_1_120 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8095 wl_0_34 wl_1_34 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8084 wl_0_45 wl_1_45 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8073 wl_0_56 wl_1_56 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7394 wl_0_126 wl_1_126 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7361 wl_0_126 wl_1_126 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7383 wl_0_120 wl_1_120 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7372 wl_0_119 wl_1_119 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6682 wl_0_76 wl_1_76 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6660 wl_0_80 wl_1_80 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6671 wl_0_87 wl_1_87 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6693 wl_0_67 wl_1_67 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5981 wl_0_70 wl_1_70 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5970 wl_0_71 wl_1_71 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5992 wl_0_73 wl_1_73 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4009 wl_0_69 wl_1_69 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3308 wl_0_34 wl_1_34 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3319 wl_0_39 wl_1_39 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2629 wl_0_27 wl_1_27 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2607 wl_0_28 wl_1_28 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2618 wl_0_27 wl_1_27 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1917 wl_0_32 wl_1_32 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1928 wl_0_31 wl_1_31 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1906 wl_0_31 wl_1_31 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1939 wl_0_32 wl_1_32 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5200 wl_0_106 wl_1_106 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5211 wl_0_126 wl_1_126 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5222 wl_0_115 wl_1_115 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5233 wl_0_104 wl_1_104 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5266 wl_0_109 wl_1_109 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5255 wl_0_105 wl_1_105 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5244 wl_0_98 wl_1_98 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4510 wl_0_82 wl_1_82 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4521 wl_0_93 wl_1_93 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5288 wl_0_110 wl_1_110 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5299 wl_0_108 wl_1_108 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5277 wl_0_101 wl_1_101 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3820 wl_0_35 wl_1_35 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4554 wl_0_82 wl_1_82 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4565 wl_0_85 wl_1_85 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4532 wl_0_86 wl_1_86 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4543 wl_0_93 wl_1_93 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3842 wl_0_15 wl_1_15 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3853 wl_0_4 wl_1_4 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3831 wl_0_26 wl_1_26 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4576 wl_0_84 wl_1_84 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4598 wl_0_86 wl_1_86 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4587 wl_0_87 wl_1_87 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3886 wl_0_32 wl_1_32 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3897 wl_0_31 wl_1_31 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3875 wl_0_31 wl_1_31 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3864 wl_0_32 wl_1_32 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7180 wl_0_110 wl_1_110 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7191 wl_0_99 wl_1_99 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6490 wl_0_86 wl_1_86 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3105 wl_0_56 wl_1_56 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3116 wl_0_61 wl_1_61 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2404 wl_0_0 wl_1_0 bl_0_9 bl_1_9 br_0_9 br_1_9
+ sky130_fd_bd_sram__openram_dp_cell_2404/a_38_n79# vdd_uq3518 gnd sky130_fd_bd_sram__openram_dp_cell_2404/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3127 wl_0_57 wl_1_57 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3138 wl_0_57 wl_1_57 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3149 wl_0_61 wl_1_61 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2426 wl_0_11 wl_1_11 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2415 wl_0_0 wl_1_0 bl_0_10 bl_1_10 br_0_10 br_1_10
+ sky130_fd_bd_sram__openram_dp_cell_2415/a_38_n79# vdd_uq3454 gnd sky130_fd_bd_sram__openram_dp_cell_2415/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2437 wl_0_5 wl_1_5 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1703 wl_0_48 wl_1_48 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2459 wl_0_8 wl_1_8 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2448 wl_0_4 wl_1_4 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1736 wl_0_33 wl_1_33 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1725 wl_0_44 wl_1_44 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1714 wl_0_55 wl_1_55 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1769 wl_0_32 wl_1_32 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1758 wl_0_41 wl_1_41 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1747 wl_0_52 wl_1_52 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5041 wl_0_124 wl_1_124 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5030 wl_0_120 wl_1_120 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5074 wl_0_123 wl_1_123 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5085 wl_0_117 wl_1_117 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5063 wl_0_117 wl_1_117 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5052 wl_0_113 wl_1_113 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4340 wl_0_67 wl_1_67 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5096 wl_0_123 wl_1_123 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4373 wl_0_70 wl_1_70 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4362 wl_0_72 wl_1_72 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4351 wl_0_73 wl_1_73 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3661 wl_0_47 wl_1_47 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3650 wl_0_48 wl_1_48 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4395 wl_0_65 wl_1_65 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4384 wl_0_74 wl_1_74 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2960 wl_0_38 wl_1_38 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3694 wl_0_40 wl_1_40 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3683 wl_0_51 wl_1_51 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3672 wl_0_62 wl_1_62 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2971 wl_0_36 wl_1_36 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2982 wl_0_42 wl_1_42 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2993 wl_0_44 wl_1_44 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7905 wl_0_96 wl_1_96 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7916 wl_0_85 wl_1_85 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7949 wl_0_52 wl_1_52 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7938 wl_0_63 wl_1_63 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7927 wl_0_74 wl_1_74 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_418 wl_0_16 wl_1_16 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_407 wl_0_4 wl_1_4 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_429 wl_0_25 wl_1_25 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2212 wl_0_17 wl_1_17 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2201 wl_0_28 wl_1_28 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2223 wl_0_27 wl_1_27 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2256 wl_0_27 wl_1_27 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2234 wl_0_27 wl_1_27 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2245 wl_0_29 wl_1_29 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1500 wl_0_34 wl_1_34 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1511 wl_0_57 wl_1_57 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2267 wl_0_21 wl_1_21 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2278 wl_0_20 wl_1_20 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2289 wl_0_30 wl_1_30 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1533 wl_0_54 wl_1_54 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1544 wl_0_58 wl_1_58 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1522 wl_0_60 wl_1_60 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1566 wl_0_49 wl_1_49 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1577 wl_0_57 wl_1_57 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1555 wl_0_60 wl_1_60 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1599 wl_0_50 wl_1_50 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1588 wl_0_61 wl_1_61 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_930 wl_0_33 wl_1_33 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_941 wl_0_45 wl_1_45 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_985 wl_0_34 wl_1_34 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_974 wl_0_37 wl_1_37 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_952 wl_0_40 wl_1_40 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_963 wl_0_41 wl_1_41 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4170 wl_0_88 wl_1_88 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4181 wl_0_93 wl_1_93 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_996 wl_0_38 wl_1_38 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3480 wl_0_54 wl_1_54 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4192 wl_0_84 wl_1_84 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3491 wl_0_55 wl_1_55 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2790 wl_0_30 wl_1_30 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7724 wl_0_126 wl_1_126 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7735 wl_0_115 wl_1_115 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7713 wl_0_74 wl_1_74 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7702 wl_0_85 wl_1_85 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7746 wl_0_104 wl_1_104 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7768 wl_0_82 wl_1_82 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7757 wl_0_93 wl_1_93 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7779 wl_0_71 wl_1_71 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_204 wl_0_29 wl_1_29 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_215 wl_0_20 wl_1_20 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_237 wl_0_17 wl_1_17 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_226 wl_0_25 wl_1_25 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_248 wl_0_19 wl_1_19 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_259 wl_0_30 wl_1_30 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2020 wl_0_14 wl_1_14 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2042 wl_0_14 wl_1_14 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2053 wl_0_14 wl_1_14 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2064 wl_0_7 wl_1_7 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2031 wl_0_3 wl_1_3 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2075 wl_0_7 wl_1_7 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2097 wl_0_1 wl_1_1 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2086 wl_0_4 wl_1_4 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1330 wl_0_35 wl_1_35 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1352 wl_0_37 wl_1_37 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1341 wl_0_39 wl_1_39 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1396 wl_0_37 wl_1_37 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1385 wl_0_38 wl_1_38 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1374 wl_0_42 wl_1_42 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1363 wl_0_46 wl_1_46 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_0 wl_0_1 wl_1_1 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_760 wl_0_21 wl_1_21 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_771 wl_0_19 wl_1_19 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_793 wl_0_18 wl_1_18 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_782 wl_0_29 wl_1_29 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7009 wl_0_121 wl_1_121 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6319 wl_0_73 wl_1_73 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6308 wl_0_79 wl_1_79 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5607 wl_0_123 wl_1_123 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5618 wl_0_112 wl_1_112 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4906 wl_0_104 wl_1_104 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5629 wl_0_101 wl_1_101 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4917 wl_0_109 wl_1_109 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4939 wl_0_104 wl_1_104 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4928 wl_0_100 wl_1_100 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7510 wl_0_125 wl_1_125 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7532 wl_0_118 wl_1_118 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7521 wl_0_114 wl_1_114 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7543 wl_0_111 wl_1_111 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7565 wl_0_118 wl_1_118 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7554 wl_0_112 wl_1_112 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6820 wl_0_110 wl_1_110 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7576 wl_0_107 wl_1_107 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6831 wl_0_105 wl_1_105 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7587 wl_0_127 wl_1_127 bl_0_55 bl_1_55 br_0_55
+ br_1_55 sky130_fd_bd_sram__openram_dp_cell_7587/a_38_n79# vdd_uq574 gnd sky130_fd_bd_sram__openram_dp_cell_7587/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7598 wl_0_116 wl_1_116 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6864 wl_0_109 wl_1_109 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6875 wl_0_102 wl_1_102 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6842 wl_0_101 wl_1_101 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6853 wl_0_99 wl_1_99 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6897 wl_0_122 wl_1_122 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6886 wl_0_101 wl_1_101 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_50 wl_0_12 wl_1_12 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_72 wl_0_12 wl_1_12 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_61 wl_0_10 wl_1_10 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_83 wl_0_7 wl_1_7 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_94 wl_0_5 wl_1_5 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1160 wl_0_57 wl_1_57 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1193 wl_0_52 wl_1_52 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1182 wl_0_56 wl_1_56 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1171 wl_0_58 wl_1_58 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_590 wl_0_8 wl_1_8 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6105 wl_0_86 wl_1_86 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6116 wl_0_87 wl_1_87 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6127 wl_0_94 wl_1_94 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5415 wl_0_116 wl_1_116 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5404 wl_0_99 wl_1_99 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6149 wl_0_84 wl_1_84 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6138 wl_0_83 wl_1_83 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5426 wl_0_124 wl_1_124 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5437 wl_0_122 wl_1_122 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5459 wl_0_119 wl_1_119 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5448 wl_0_119 wl_1_119 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4714 wl_0_82 wl_1_82 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4703 wl_0_93 wl_1_93 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4736 wl_0_66 wl_1_66 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4725 wl_0_73 wl_1_73 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4747 wl_0_85 wl_1_85 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4758 wl_0_74 wl_1_74 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4769 wl_0_79 wl_1_79 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8030 wl_0_99 wl_1_99 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8063 wl_0_66 wl_1_66 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8052 wl_0_77 wl_1_77 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8041 wl_0_88 wl_1_88 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7351 wl_0_119 wl_1_119 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7340 wl_0_99 wl_1_99 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8096 wl_0_33 wl_1_33 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8085 wl_0_44 wl_1_44 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8074 wl_0_55 wl_1_55 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7362 wl_0_124 wl_1_124 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7384 wl_0_119 wl_1_119 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7373 wl_0_118 wl_1_118 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7395 wl_0_125 wl_1_125 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6683 wl_0_75 wl_1_75 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6661 wl_0_79 wl_1_79 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6650 wl_0_80 wl_1_80 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6672 wl_0_86 wl_1_86 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6694 wl_0_66 wl_1_66 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5971 wl_0_70 wl_1_70 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5960 wl_0_74 wl_1_74 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5982 wl_0_69 wl_1_69 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5993 wl_0_72 wl_1_72 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3309 wl_0_33 wl_1_33 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2619 wl_0_26 wl_1_26 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2608 wl_0_30 wl_1_30 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1907 wl_0_32 wl_1_32 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1918 wl_0_31 wl_1_31 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1929 wl_0_32 wl_1_32 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5212 wl_0_125 wl_1_125 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5223 wl_0_114 wl_1_114 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5201 wl_0_105 wl_1_105 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5234 wl_0_103 wl_1_103 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5267 wl_0_108 wl_1_108 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5256 wl_0_104 wl_1_104 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5245 wl_0_97 wl_1_97 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4500 wl_0_78 wl_1_78 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4511 wl_0_81 wl_1_81 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4522 wl_0_94 wl_1_94 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5289 wl_0_109 wl_1_109 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5278 wl_0_100 wl_1_100 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3810 wl_0_45 wl_1_45 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4555 wl_0_81 wl_1_81 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4533 wl_0_85 wl_1_85 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4544 wl_0_92 wl_1_92 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3843 wl_0_14 wl_1_14 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3854 wl_0_3 wl_1_3 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3832 wl_0_25 wl_1_25 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3821 wl_0_34 wl_1_34 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4577 wl_0_83 wl_1_83 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4566 wl_0_84 wl_1_84 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4599 wl_0_85 wl_1_85 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4588 wl_0_86 wl_1_86 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3876 wl_0_32 wl_1_32 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3887 wl_0_31 wl_1_31 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3865 wl_0_31 wl_1_31 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3898 wl_0_32 wl_1_32 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7181 wl_0_109 wl_1_109 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7192 wl_0_98 wl_1_98 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7170 wl_0_98 wl_1_98 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6480 wl_0_82 wl_1_82 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6491 wl_0_85 wl_1_85 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5790 wl_0_115 wl_1_115 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3106 wl_0_55 wl_1_55 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2405 wl_0_9 wl_1_9 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3128 wl_0_56 wl_1_56 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3139 wl_0_56 wl_1_56 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3117 wl_0_60 wl_1_60 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2416 wl_0_14 wl_1_14 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2427 wl_0_10 wl_1_10 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2438 wl_0_4 wl_1_4 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2449 wl_0_3 wl_1_3 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1726 wl_0_43 wl_1_43 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1704 wl_0_47 wl_1_47 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1715 wl_0_54 wl_1_54 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1759 wl_0_40 wl_1_40 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1748 wl_0_51 wl_1_51 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1737 wl_0_62 wl_1_62 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5042 wl_0_123 wl_1_123 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5020 wl_0_122 wl_1_122 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5031 wl_0_119 wl_1_119 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5075 wl_0_127 wl_1_127 bl_0_14 bl_1_14 br_0_14
+ br_1_14 sky130_fd_bd_sram__openram_dp_cell_5075/a_38_n79# vdd_uq3198 gnd sky130_fd_bd_sram__openram_dp_cell_5075/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5053 wl_0_120 wl_1_120 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5064 wl_0_116 wl_1_116 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4330 wl_0_77 wl_1_77 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5097 wl_0_122 wl_1_122 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5086 wl_0_116 wl_1_116 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4341 wl_0_66 wl_1_66 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4352 wl_0_72 wl_1_72 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4363 wl_0_71 wl_1_71 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3640 wl_0_48 wl_1_48 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3651 wl_0_47 wl_1_47 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3662 wl_0_48 wl_1_48 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4374 wl_0_69 wl_1_69 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4385 wl_0_73 wl_1_73 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4396 wl_0_76 wl_1_76 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3695 wl_0_39 wl_1_39 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2950 wl_0_43 wl_1_43 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3684 wl_0_50 wl_1_50 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3673 wl_0_61 wl_1_61 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2972 wl_0_35 wl_1_35 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2961 wl_0_37 wl_1_37 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2983 wl_0_41 wl_1_41 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2994 wl_0_43 wl_1_43 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7906 wl_0_95 wl_1_95 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7917 wl_0_84 wl_1_84 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7939 wl_0_62 wl_1_62 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7928 wl_0_73 wl_1_73 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_419 wl_0_15 wl_1_15 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_408 wl_0_3 wl_1_3 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2213 wl_0_23 wl_1_23 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2202 wl_0_27 wl_1_27 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2224 wl_0_26 wl_1_26 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2235 wl_0_26 wl_1_26 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2246 wl_0_28 wl_1_28 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1501 wl_0_53 wl_1_53 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2279 wl_0_19 wl_1_19 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2257 wl_0_26 wl_1_26 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2268 wl_0_30 wl_1_30 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1534 wl_0_53 wl_1_53 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1512 wl_0_56 wl_1_56 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1545 wl_0_57 wl_1_57 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1523 wl_0_59 wl_1_59 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1567 wl_0_56 wl_1_56 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1578 wl_0_56 wl_1_56 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1556 wl_0_59 wl_1_59 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1589 wl_0_60 wl_1_60 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_920 wl_0_43 wl_1_43 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_942 wl_0_44 wl_1_44 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_931 wl_0_46 wl_1_46 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_975 wl_0_36 wl_1_36 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_964 wl_0_40 wl_1_40 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_953 wl_0_39 wl_1_39 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4171 wl_0_87 wl_1_87 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4160 wl_0_88 wl_1_88 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4182 wl_0_94 wl_1_94 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_997 wl_0_37 wl_1_37 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_986 wl_0_46 wl_1_46 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3470 wl_0_54 wl_1_54 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4193 wl_0_83 wl_1_83 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3481 wl_0_53 wl_1_53 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3492 wl_0_62 wl_1_62 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2780 wl_0_16 wl_1_16 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2791 wl_0_29 wl_1_29 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7725 wl_0_125 wl_1_125 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7714 wl_0_73 wl_1_73 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7703 wl_0_84 wl_1_84 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7736 wl_0_114 wl_1_114 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7747 wl_0_103 wl_1_103 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7758 wl_0_92 wl_1_92 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7769 wl_0_81 wl_1_81 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_216 wl_0_19 wl_1_19 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_238 wl_0_24 wl_1_24 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_227 wl_0_24 wl_1_24 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_205 wl_0_30 wl_1_30 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_249 wl_0_18 wl_1_18 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2021 wl_0_13 wl_1_13 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2010 wl_0_3 wl_1_3 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2054 wl_0_13 wl_1_13 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2043 wl_0_12 wl_1_12 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2032 wl_0_2 wl_1_2 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2065 wl_0_6 wl_1_6 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2076 wl_0_6 wl_1_6 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2098 wl_0_1 wl_1_1 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2087 wl_0_3 wl_1_3 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1331 wl_0_34 wl_1_34 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1353 wl_0_36 wl_1_36 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1342 wl_0_38 wl_1_38 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1320 wl_0_45 wl_1_45 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1386 wl_0_37 wl_1_37 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1375 wl_0_41 wl_1_41 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1364 wl_0_45 wl_1_45 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1397 wl_0_36 wl_1_36 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1 wl_0_0 wl_1_0 bl_0_63 bl_1_63 br_0_63 br_1_63
+ sky130_fd_bd_sram__openram_dp_cell_1/a_38_n79# vdd gnd sky130_fd_bd_sram__openram_dp_cell_1/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_750 wl_0_22 wl_1_22 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_772 wl_0_18 wl_1_18 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_761 wl_0_25 wl_1_25 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_783 wl_0_28 wl_1_28 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_794 wl_0_17 wl_1_17 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6309 wl_0_72 wl_1_72 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5608 wl_0_122 wl_1_122 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5619 wl_0_111 wl_1_111 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4907 wl_0_103 wl_1_103 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4929 wl_0_99 wl_1_99 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4918 wl_0_100 wl_1_100 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7500 wl_0_120 wl_1_120 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7511 wl_0_124 wl_1_124 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7533 wl_0_117 wl_1_117 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7522 wl_0_113 wl_1_113 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7566 wl_0_117 wl_1_117 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7544 wl_0_112 wl_1_112 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7555 wl_0_111 wl_1_111 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6821 wl_0_109 wl_1_109 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7577 wl_0_106 wl_1_106 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6810 wl_0_104 wl_1_104 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6832 wl_0_104 wl_1_104 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7588 wl_0_126 wl_1_126 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7599 wl_0_115 wl_1_115 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6865 wl_0_108 wl_1_108 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6843 wl_0_100 wl_1_100 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6854 wl_0_98 wl_1_98 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6898 wl_0_121 wl_1_121 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6887 wl_0_103 wl_1_103 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6876 wl_0_101 wl_1_101 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_40 wl_0_9 wl_1_9 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_51 wl_0_11 wl_1_11 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_73 wl_0_11 wl_1_11 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_62 wl_0_9 wl_1_9 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_84 wl_0_6 wl_1_6 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_95 wl_0_4 wl_1_4 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1161 wl_0_49 wl_1_49 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1150 wl_0_53 wl_1_53 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1194 wl_0_51 wl_1_51 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1172 wl_0_57 wl_1_57 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1183 wl_0_62 wl_1_62 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_591 wl_0_14 wl_1_14 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_580 wl_0_6 wl_1_6 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6106 wl_0_85 wl_1_85 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6117 wl_0_86 wl_1_86 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5416 wl_0_115 wl_1_115 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5405 wl_0_105 wl_1_105 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6139 wl_0_82 wl_1_82 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6128 wl_0_93 wl_1_93 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5449 wl_0_127 wl_1_127 bl_0_21 bl_1_21 br_0_21
+ br_1_21 sky130_fd_bd_sram__openram_dp_cell_5449/a_38_n79# vdd_uq2750 gnd sky130_fd_bd_sram__openram_dp_cell_5449/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5427 wl_0_123 wl_1_123 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5438 wl_0_121 wl_1_121 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4704 wl_0_92 wl_1_92 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4737 wl_0_65 wl_1_65 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4726 wl_0_72 wl_1_72 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4715 wl_0_81 wl_1_81 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4748 wl_0_84 wl_1_84 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4759 wl_0_73 wl_1_73 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8020 wl_0_109 wl_1_109 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8031 wl_0_98 wl_1_98 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8053 wl_0_76 wl_1_76 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8042 wl_0_87 wl_1_87 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7341 wl_0_110 wl_1_110 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7330 wl_0_109 wl_1_109 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8086 wl_0_43 wl_1_43 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8075 wl_0_54 wl_1_54 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8064 wl_0_65 wl_1_65 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7374 wl_0_127 wl_1_127 bl_0_54 bl_1_54 br_0_54
+ br_1_54 sky130_fd_bd_sram__openram_dp_cell_7374/a_38_n79# vdd_uq638 gnd sky130_fd_bd_sram__openram_dp_cell_7374/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7363 wl_0_123 wl_1_123 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7385 wl_0_118 wl_1_118 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7352 wl_0_118 wl_1_118 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8097 wl_0_32 wl_1_32 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6640 wl_0_82 wl_1_82 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7396 wl_0_124 wl_1_124 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6662 wl_0_80 wl_1_80 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6651 wl_0_79 wl_1_79 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6673 wl_0_85 wl_1_85 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6695 wl_0_65 wl_1_65 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5972 wl_0_69 wl_1_69 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5950 wl_0_71 wl_1_71 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5961 wl_0_73 wl_1_73 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6684 wl_0_74 wl_1_74 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5983 wl_0_68 wl_1_68 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5994 wl_0_69 wl_1_69 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2609 wl_0_29 wl_1_29 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1908 wl_0_31 wl_1_31 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1919 wl_0_32 wl_1_32 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5213 wl_0_124 wl_1_124 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5224 wl_0_113 wl_1_113 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5202 wl_0_104 wl_1_104 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5257 wl_0_103 wl_1_103 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5235 wl_0_102 wl_1_102 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5246 wl_0_101 wl_1_101 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4501 wl_0_77 wl_1_77 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4512 wl_0_93 wl_1_93 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5268 wl_0_110 wl_1_110 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5279 wl_0_99 wl_1_99 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3811 wl_0_44 wl_1_44 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3800 wl_0_55 wl_1_55 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4534 wl_0_84 wl_1_84 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4545 wl_0_91 wl_1_91 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4523 wl_0_93 wl_1_93 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4556 wl_0_94 wl_1_94 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3833 wl_0_24 wl_1_24 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3844 wl_0_13 wl_1_13 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3822 wl_0_33 wl_1_33 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4578 wl_0_82 wl_1_82 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4567 wl_0_83 wl_1_83 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4589 wl_0_85 wl_1_85 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3855 wl_0_2 wl_1_2 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3877 wl_0_31 wl_1_31 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3888 wl_0_32 wl_1_32 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3866 wl_0_32 wl_1_32 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3899 wl_0_31 wl_1_31 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7160 wl_0_111 wl_1_111 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7182 wl_0_108 wl_1_108 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7193 wl_0_97 wl_1_97 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7171 wl_0_97 wl_1_97 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6470 wl_0_75 wl_1_75 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6481 wl_0_81 wl_1_81 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5780 wl_0_125 wl_1_125 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6492 wl_0_84 wl_1_84 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5791 wl_0_114 wl_1_114 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3107 wl_0_60 wl_1_60 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3129 wl_0_55 wl_1_55 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3118 wl_0_59 wl_1_59 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2428 wl_0_14 wl_1_14 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2417 wl_0_13 wl_1_13 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2406 wl_0_8 wl_1_8 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2439 wl_0_3 wl_1_3 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1727 wl_0_42 wl_1_42 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1705 wl_0_48 wl_1_48 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1716 wl_0_53 wl_1_53 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1749 wl_0_50 wl_1_50 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1738 wl_0_61 wl_1_61 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5021 wl_0_126 wl_1_126 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5010 wl_0_124 wl_1_124 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5032 wl_0_118 wl_1_118 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5076 wl_0_126 wl_1_126 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5043 wl_0_122 wl_1_122 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5054 wl_0_119 wl_1_119 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5065 wl_0_115 wl_1_115 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4320 wl_0_66 wl_1_66 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4331 wl_0_76 wl_1_76 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5098 wl_0_121 wl_1_121 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5087 wl_0_115 wl_1_115 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4342 wl_0_65 wl_1_65 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4364 wl_0_70 wl_1_70 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4353 wl_0_71 wl_1_71 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3641 wl_0_47 wl_1_47 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3652 wl_0_48 wl_1_48 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3630 wl_0_56 wl_1_56 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4375 wl_0_68 wl_1_68 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4397 wl_0_68 wl_1_68 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4386 wl_0_72 wl_1_72 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3696 wl_0_38 wl_1_38 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2940 wl_0_41 wl_1_41 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2951 wl_0_42 wl_1_42 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3663 wl_0_47 wl_1_47 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3685 wl_0_49 wl_1_49 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3674 wl_0_60 wl_1_60 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2973 wl_0_36 wl_1_36 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2962 wl_0_36 wl_1_36 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2984 wl_0_40 wl_1_40 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2995 wl_0_42 wl_1_42 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7907 wl_0_94 wl_1_94 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7929 wl_0_72 wl_1_72 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7918 wl_0_83 wl_1_83 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_409 wl_0_2 wl_1_2 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2203 wl_0_26 wl_1_26 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2214 wl_0_22 wl_1_22 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2225 wl_0_25 wl_1_25 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2236 wl_0_25 wl_1_25 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2247 wl_0_27 wl_1_27 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1502 wl_0_52 wl_1_52 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2258 wl_0_25 wl_1_25 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2269 wl_0_29 wl_1_29 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1535 wl_0_52 wl_1_52 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1513 wl_0_55 wl_1_55 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1524 wl_0_58 wl_1_58 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1568 wl_0_55 wl_1_55 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1546 wl_0_56 wl_1_56 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1557 wl_0_58 wl_1_58 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1579 wl_0_55 wl_1_55 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_921 wl_0_42 wl_1_42 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_910 wl_0_43 wl_1_43 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_932 wl_0_46 wl_1_46 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_965 wl_0_34 wl_1_34 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_976 wl_0_35 wl_1_35 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_954 wl_0_38 wl_1_38 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_943 wl_0_43 wl_1_43 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4172 wl_0_86 wl_1_86 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4161 wl_0_87 wl_1_87 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4150 wl_0_89 wl_1_89 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3460 wl_0_34 wl_1_34 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_987 wl_0_45 wl_1_45 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_998 wl_0_46 wl_1_46 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3471 wl_0_53 wl_1_53 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4194 wl_0_82 wl_1_82 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4183 wl_0_93 wl_1_93 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3482 wl_0_52 wl_1_52 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3493 wl_0_61 wl_1_61 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2781 wl_0_15 wl_1_15 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2770 wl_0_26 wl_1_26 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2792 wl_0_28 wl_1_28 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7726 wl_0_124 wl_1_124 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7715 wl_0_72 wl_1_72 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7704 wl_0_83 wl_1_83 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7737 wl_0_113 wl_1_113 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7748 wl_0_102 wl_1_102 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7759 wl_0_91 wl_1_91 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_217 wl_0_18 wl_1_18 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_228 wl_0_26 wl_1_26 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_206 wl_0_29 wl_1_29 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_239 wl_0_23 wl_1_23 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2000 wl_0_9 wl_1_9 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2011 wl_0_2 wl_1_2 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2044 wl_0_14 wl_1_14 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2022 wl_0_12 wl_1_12 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2055 wl_0_12 wl_1_12 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2033 wl_0_1 wl_1_1 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1310 wl_0_48 wl_1_48 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2088 wl_0_2 wl_1_2 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2077 wl_0_5 wl_1_5 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2066 wl_0_5 wl_1_5 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1332 wl_0_33 wl_1_33 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1343 wl_0_37 wl_1_37 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1321 wl_0_44 wl_1_44 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2099 wl_0_0 wl_1_0 bl_0_22 bl_1_22 br_0_22 br_1_22
+ sky130_fd_bd_sram__openram_dp_cell_2099/a_38_n79# vdd_uq2686 gnd sky130_fd_bd_sram__openram_dp_cell_2099/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1354 wl_0_35 wl_1_35 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1376 wl_0_40 wl_1_40 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1365 wl_0_44 wl_1_44 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1398 wl_0_35 wl_1_35 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1387 wl_0_46 wl_1_46 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2 wl_0_3 wl_1_3 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_740 wl_0_24 wl_1_24 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_751 wl_0_30 wl_1_30 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_773 wl_0_17 wl_1_17 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_762 wl_0_24 wl_1_24 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_784 wl_0_27 wl_1_27 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_795 wl_0_24 wl_1_24 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3290 wl_0_35 wl_1_35 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5609 wl_0_121 wl_1_121 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4919 wl_0_102 wl_1_102 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4908 wl_0_102 wl_1_102 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7523 wl_0_127 wl_1_127 bl_0_59 bl_1_59 br_0_59
+ br_1_59 sky130_fd_bd_sram__openram_dp_cell_7523/a_38_n79# vdd_uq318 gnd sky130_fd_bd_sram__openram_dp_cell_7523/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7512 wl_0_123 wl_1_123 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7501 wl_0_119 wl_1_119 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7534 wl_0_116 wl_1_116 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7556 wl_0_127 wl_1_127 bl_0_56 bl_1_56 br_0_56
+ br_1_56 sky130_fd_bd_sram__openram_dp_cell_7556/a_38_n79# vdd_uq510 gnd sky130_fd_bd_sram__openram_dp_cell_7556/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7567 wl_0_116 wl_1_116 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7545 wl_0_111 wl_1_111 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6822 wl_0_108 wl_1_108 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6800 wl_0_106 wl_1_106 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6811 wl_0_103 wl_1_103 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7589 wl_0_125 wl_1_125 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6833 wl_0_106 wl_1_106 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7578 wl_0_105 wl_1_105 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6844 wl_0_104 wl_1_104 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6855 wl_0_97 wl_1_97 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6899 wl_0_120 wl_1_120 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6888 wl_0_102 wl_1_102 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6877 wl_0_100 wl_1_100 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6866 wl_0_98 wl_1_98 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_41 wl_0_14 wl_1_14 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_30 wl_0_3 wl_1_3 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_63 wl_0_14 wl_1_14 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_52 wl_0_10 wl_1_10 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_74 wl_0_10 wl_1_10 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_96 wl_0_3 wl_1_3 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_85 wl_0_5 wl_1_5 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1151 wl_0_51 wl_1_51 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1140 wl_0_54 wl_1_54 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1195 wl_0_50 wl_1_50 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1173 wl_0_56 wl_1_56 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1184 wl_0_61 wl_1_61 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1162 wl_0_62 wl_1_62 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_592 wl_0_13 wl_1_13 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_570 wl_0_12 wl_1_12 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_581 wl_0_9 wl_1_9 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6107 wl_0_84 wl_1_84 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6118 wl_0_85 wl_1_85 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5406 wl_0_104 wl_1_104 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6129 wl_0_92 wl_1_92 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5428 wl_0_122 wl_1_122 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5439 wl_0_120 wl_1_120 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5417 wl_0_114 wl_1_114 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4705 wl_0_91 wl_1_91 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4727 wl_0_71 wl_1_71 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4716 wl_0_80 wl_1_80 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4738 wl_0_94 wl_1_94 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4749 wl_0_83 wl_1_83 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8010 wl_0_119 wl_1_119 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8021 wl_0_108 wl_1_108 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8032 wl_0_97 wl_1_97 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8054 wl_0_75 wl_1_75 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8043 wl_0_86 wl_1_86 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7342 wl_0_109 wl_1_109 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7331 wl_0_108 wl_1_108 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7320 wl_0_99 wl_1_99 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8087 wl_0_42 wl_1_42 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8076 wl_0_53 wl_1_53 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8065 wl_0_64 wl_1_64 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7375 wl_0_126 wl_1_126 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7364 wl_0_125 wl_1_125 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7353 wl_0_117 wl_1_117 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8098 wl_0_31 wl_1_31 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6630 wl_0_92 wl_1_92 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7397 wl_0_123 wl_1_123 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7386 wl_0_117 wl_1_117 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6663 wl_0_79 wl_1_79 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6652 wl_0_80 wl_1_80 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6641 wl_0_81 wl_1_81 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6674 wl_0_84 wl_1_84 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5940 wl_0_66 wl_1_66 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5951 wl_0_70 wl_1_70 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5962 wl_0_72 wl_1_72 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6685 wl_0_73 wl_1_73 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6696 wl_0_80 wl_1_80 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5995 wl_0_68 wl_1_68 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5984 wl_0_67 wl_1_67 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5973 wl_0_68 wl_1_68 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1909 wl_0_32 wl_1_32 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5214 wl_0_123 wl_1_123 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5225 wl_0_112 wl_1_112 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5203 wl_0_103 wl_1_103 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5258 wl_0_102 wl_1_102 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5236 wl_0_101 wl_1_101 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5247 wl_0_100 wl_1_100 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4502 wl_0_76 wl_1_76 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4513 wl_0_83 wl_1_83 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5269 wl_0_109 wl_1_109 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3801 wl_0_54 wl_1_54 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4535 wl_0_83 wl_1_83 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4546 wl_0_90 wl_1_90 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4524 wl_0_94 wl_1_94 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3834 wl_0_23 wl_1_23 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3845 wl_0_12 wl_1_12 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3823 wl_0_32 wl_1_32 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3812 wl_0_43 wl_1_43 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4579 wl_0_81 wl_1_81 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4568 wl_0_82 wl_1_82 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4557 wl_0_93 wl_1_93 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3856 wl_0_1 wl_1_1 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3878 wl_0_32 wl_1_32 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3867 wl_0_31 wl_1_31 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3889 wl_0_31 wl_1_31 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7150 wl_0_111 wl_1_111 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7161 wl_0_112 wl_1_112 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7183 wl_0_107 wl_1_107 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7172 wl_0_101 wl_1_101 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7194 wl_0_98 wl_1_98 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6460 wl_0_72 wl_1_72 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6471 wl_0_74 wl_1_74 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6482 wl_0_94 wl_1_94 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5770 wl_0_70 wl_1_70 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6493 wl_0_83 wl_1_83 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5781 wl_0_124 wl_1_124 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5792 wl_0_113 wl_1_113 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3119 wl_0_58 wl_1_58 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3108 wl_0_59 wl_1_59 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2429 wl_0_13 wl_1_13 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2418 wl_0_12 wl_1_12 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2407 wl_0_7 wl_1_7 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1706 wl_0_47 wl_1_47 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1717 wl_0_52 wl_1_52 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1728 wl_0_41 wl_1_41 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1739 wl_0_60 wl_1_60 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5022 wl_0_125 wl_1_125 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5011 wl_0_123 wl_1_123 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5000 wl_0_121 wl_1_121 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5033 wl_0_117 wl_1_117 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5044 wl_0_121 wl_1_121 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5055 wl_0_120 wl_1_120 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5066 wl_0_114 wl_1_114 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4321 wl_0_65 wl_1_65 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4310 wl_0_76 wl_1_76 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5077 wl_0_125 wl_1_125 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5099 wl_0_120 wl_1_120 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5088 wl_0_114 wl_1_114 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3620 wl_0_50 wl_1_50 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4343 wl_0_66 wl_1_66 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4354 wl_0_70 wl_1_70 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4332 wl_0_75 wl_1_75 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3642 wl_0_40 wl_1_40 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3653 wl_0_47 wl_1_47 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3631 wl_0_55 wl_1_55 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4398 wl_0_65 wl_1_65 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4376 wl_0_67 wl_1_67 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4387 wl_0_71 wl_1_71 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4365 wl_0_78 wl_1_78 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2941 wl_0_40 wl_1_40 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2930 wl_0_41 wl_1_41 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3686 wl_0_48 wl_1_48 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3664 wl_0_48 wl_1_48 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3675 wl_0_59 wl_1_59 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2974 wl_0_35 wl_1_35 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2963 wl_0_35 wl_1_35 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3697 wl_0_37 wl_1_37 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2985 wl_0_39 wl_1_39 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2952 wl_0_46 wl_1_46 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2996 wl_0_46 wl_1_46 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6290 wl_0_67 wl_1_67 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7908 wl_0_93 wl_1_93 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7919 wl_0_82 wl_1_82 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2204 wl_0_25 wl_1_25 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2237 wl_0_24 wl_1_24 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2226 wl_0_24 wl_1_24 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2215 wl_0_21 wl_1_21 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2259 wl_0_24 wl_1_24 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2248 wl_0_26 wl_1_26 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1503 wl_0_51 wl_1_51 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1514 wl_0_54 wl_1_54 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1525 wl_0_57 wl_1_57 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1536 wl_0_51 wl_1_51 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1569 wl_0_54 wl_1_54 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1547 wl_0_55 wl_1_55 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1558 wl_0_57 wl_1_57 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_900 wl_0_37 wl_1_37 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_922 wl_0_41 wl_1_41 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_911 wl_0_42 wl_1_42 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_933 wl_0_45 wl_1_45 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_966 wl_0_33 wl_1_33 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_955 wl_0_37 wl_1_37 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_944 wl_0_42 wl_1_42 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4173 wl_0_85 wl_1_85 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4162 wl_0_86 wl_1_86 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4140 wl_0_88 wl_1_88 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4151 wl_0_88 wl_1_88 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3461 wl_0_33 wl_1_33 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_977 wl_0_34 wl_1_34 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3450 wl_0_44 wl_1_44 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_999 wl_0_45 wl_1_45 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_988 wl_0_46 wl_1_46 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4195 wl_0_81 wl_1_81 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4184 wl_0_92 wl_1_92 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2760 wl_0_20 wl_1_20 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3483 wl_0_51 wl_1_51 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3494 wl_0_60 wl_1_60 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3472 wl_0_62 wl_1_62 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2782 wl_0_14 wl_1_14 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2771 wl_0_25 wl_1_25 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2793 wl_0_27 wl_1_27 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7716 wl_0_71 wl_1_71 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7705 wl_0_82 wl_1_82 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7727 wl_0_123 wl_1_123 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7738 wl_0_112 wl_1_112 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7749 wl_0_101 wl_1_101 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_218 wl_0_17 wl_1_17 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_229 wl_0_25 wl_1_25 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_207 wl_0_28 wl_1_28 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2012 wl_0_14 wl_1_14 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2001 wl_0_8 wl_1_8 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2045 wl_0_13 wl_1_13 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2023 wl_0_11 wl_1_11 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2034 wl_0_0 wl_1_0 bl_0_27 bl_1_27 br_0_27 br_1_27
+ sky130_fd_bd_sram__openram_dp_cell_2034/a_38_n79# vdd_uq2366 gnd sky130_fd_bd_sram__openram_dp_cell_2034/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1300 wl_0_48 wl_1_48 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2056 wl_0_11 wl_1_11 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2089 wl_0_9 wl_1_9 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2078 wl_0_4 wl_1_4 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2067 wl_0_4 wl_1_4 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1333 wl_0_36 wl_1_36 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1344 wl_0_36 wl_1_36 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1322 wl_0_43 wl_1_43 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1311 wl_0_47 wl_1_47 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1355 wl_0_34 wl_1_34 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1377 wl_0_39 wl_1_39 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1366 wl_0_43 wl_1_43 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1399 wl_0_34 wl_1_34 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1388 wl_0_45 wl_1_45 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3 wl_0_6 wl_1_6 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_741 wl_0_23 wl_1_23 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_730 wl_0_29 wl_1_29 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_774 wl_0_21 wl_1_21 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_763 wl_0_23 wl_1_23 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_752 wl_0_29 wl_1_29 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_796 wl_0_17 wl_1_17 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_785 wl_0_26 wl_1_26 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3291 wl_0_34 wl_1_34 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3280 wl_0_45 wl_1_45 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2590 wl_0_25 wl_1_25 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4909 wl_0_101 wl_1_101 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7524 wl_0_126 wl_1_126 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7513 wl_0_122 wl_1_122 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7502 wl_0_120 wl_1_120 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7557 wl_0_126 wl_1_126 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7535 wl_0_115 wl_1_115 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7568 wl_0_115 wl_1_115 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7546 wl_0_112 wl_1_112 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6823 wl_0_107 wl_1_107 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6801 wl_0_105 wl_1_105 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6812 wl_0_102 wl_1_102 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6834 wl_0_105 wl_1_105 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6845 wl_0_105 wl_1_105 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7579 wl_0_104 wl_1_104 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6856 wl_0_97 wl_1_97 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6889 wl_0_108 wl_1_108 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6878 wl_0_99 wl_1_99 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6867 wl_0_97 wl_1_97 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_31 wl_0_2 wl_1_2 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_20 wl_0_2 wl_1_2 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_64 wl_0_13 wl_1_13 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_42 wl_0_13 wl_1_13 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_53 wl_0_9 wl_1_9 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_75 wl_0_9 wl_1_9 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_97 wl_0_2 wl_1_2 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_86 wl_0_4 wl_1_4 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1130 wl_0_49 wl_1_49 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1152 wl_0_50 wl_1_50 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1141 wl_0_62 wl_1_62 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1174 wl_0_55 wl_1_55 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1185 wl_0_60 wl_1_60 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1163 wl_0_61 wl_1_61 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1196 wl_0_55 wl_1_55 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_571 wl_0_11 wl_1_11 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_593 wl_0_12 wl_1_12 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_582 wl_0_8 wl_1_8 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_560 wl_0_6 wl_1_6 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6108 wl_0_83 wl_1_83 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5407 wl_0_103 wl_1_103 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6119 wl_0_84 wl_1_84 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5429 wl_0_121 wl_1_121 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5418 wl_0_113 wl_1_113 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4728 wl_0_70 wl_1_70 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4717 wl_0_79 wl_1_79 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4706 wl_0_90 wl_1_90 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4739 wl_0_93 wl_1_93 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8011 wl_0_118 wl_1_118 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8000 wl_0_1 wl_1_1 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8022 wl_0_107 wl_1_107 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8044 wl_0_85 wl_1_85 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8033 wl_0_96 wl_1_96 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7310 wl_0_109 wl_1_109 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7332 wl_0_107 wl_1_107 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7321 wl_0_98 wl_1_98 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8077 wl_0_52 wl_1_52 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8066 wl_0_63 wl_1_63 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8055 wl_0_74 wl_1_74 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7376 wl_0_125 wl_1_125 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7365 wl_0_124 wl_1_124 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7354 wl_0_116 wl_1_116 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7343 wl_0_98 wl_1_98 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8099 wl_0_30 wl_1_30 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8088 wl_0_41 wl_1_41 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6620 wl_0_89 wl_1_89 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6631 wl_0_91 wl_1_91 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7398 wl_0_122 wl_1_122 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7387 wl_0_116 wl_1_116 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6653 wl_0_79 wl_1_79 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6642 wl_0_81 wl_1_81 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6664 wl_0_94 wl_1_94 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5941 wl_0_65 wl_1_65 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5952 wl_0_69 wl_1_69 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6686 wl_0_72 wl_1_72 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5930 wl_0_76 wl_1_76 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5963 wl_0_78 wl_1_78 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6697 wl_0_79 wl_1_79 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6675 wl_0_83 wl_1_83 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5985 wl_0_66 wl_1_66 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5996 wl_0_67 wl_1_67 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5974 wl_0_67 wl_1_67 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_390 wl_0_19 wl_1_19 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5215 wl_0_122 wl_1_122 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5204 wl_0_102 wl_1_102 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5226 wl_0_111 wl_1_111 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5248 wl_0_99 wl_1_99 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5237 wl_0_100 wl_1_100 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4503 wl_0_75 wl_1_75 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5259 wl_0_101 wl_1_101 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3802 wl_0_53 wl_1_53 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4536 wl_0_82 wl_1_82 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4547 wl_0_89 wl_1_89 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4514 wl_0_92 wl_1_92 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4525 wl_0_93 wl_1_93 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3835 wl_0_22 wl_1_22 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3824 wl_0_31 wl_1_31 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3813 wl_0_42 wl_1_42 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4569 wl_0_81 wl_1_81 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4558 wl_0_92 wl_1_92 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3846 wl_0_11 wl_1_11 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3857 wl_0_0 wl_1_0 bl_0_15 bl_1_15 br_0_15 br_1_15
+ sky130_fd_bd_sram__openram_dp_cell_3857/a_38_n79# vdd_uq3134 gnd sky130_fd_bd_sram__openram_dp_cell_3857/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3868 wl_0_32 wl_1_32 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3879 wl_0_31 wl_1_31 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7151 wl_0_112 wl_1_112 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7140 wl_0_111 wl_1_111 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7162 wl_0_111 wl_1_111 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7184 wl_0_106 wl_1_106 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7173 wl_0_100 wl_1_100 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7195 wl_0_110 wl_1_110 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6450 wl_0_65 wl_1_65 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6461 wl_0_71 wl_1_71 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6472 wl_0_73 wl_1_73 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5771 wl_0_69 wl_1_69 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5760 wl_0_80 wl_1_80 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6494 wl_0_82 wl_1_82 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6483 wl_0_93 wl_1_93 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5782 wl_0_123 wl_1_123 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5793 wl_0_112 wl_1_112 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3109 wl_0_58 wl_1_58 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2419 wl_0_11 wl_1_11 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2408 wl_0_6 wl_1_6 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1718 wl_0_51 wl_1_51 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1707 wl_0_62 wl_1_62 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1729 wl_0_40 wl_1_40 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5023 wl_0_127 wl_1_127 bl_0_4 bl_1_4 br_0_4 br_1_4
+ sky130_fd_bd_sram__openram_dp_cell_5023/a_38_n79# vdd_uq3838 gnd sky130_fd_bd_sram__openram_dp_cell_5023/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5001 wl_0_123 wl_1_123 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5012 wl_0_122 wl_1_122 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5045 wl_0_120 wl_1_120 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5056 wl_0_120 wl_1_120 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5034 wl_0_116 wl_1_116 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5067 wl_0_113 wl_1_113 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4311 wl_0_75 wl_1_75 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4322 wl_0_80 wl_1_80 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4300 wl_0_86 wl_1_86 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5078 wl_0_124 wl_1_124 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5089 wl_0_113 wl_1_113 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3610 wl_0_60 wl_1_60 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4344 wl_0_65 wl_1_65 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4355 wl_0_69 wl_1_69 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4333 wl_0_74 wl_1_74 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3643 wl_0_39 wl_1_39 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3621 wl_0_49 wl_1_49 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3632 wl_0_54 wl_1_54 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4377 wl_0_66 wl_1_66 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4388 wl_0_70 wl_1_70 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4366 wl_0_77 wl_1_77 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2920 wl_0_38 wl_1_38 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2942 wl_0_39 wl_1_39 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2931 wl_0_42 wl_1_42 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3654 wl_0_48 wl_1_48 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3687 wl_0_47 wl_1_47 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3665 wl_0_47 wl_1_47 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3676 wl_0_58 wl_1_58 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4399 wl_0_67 wl_1_67 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2975 wl_0_34 wl_1_34 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2964 wl_0_34 wl_1_34 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3698 wl_0_36 wl_1_36 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2953 wl_0_45 wl_1_45 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2997 wl_0_37 wl_1_37 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2986 wl_0_38 wl_1_38 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6291 wl_0_66 wl_1_66 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6280 wl_0_77 wl_1_77 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5590 wl_0_111 wl_1_111 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7909 wl_0_92 wl_1_92 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2238 wl_0_23 wl_1_23 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2227 wl_0_23 wl_1_23 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2205 wl_0_24 wl_1_24 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2216 wl_0_20 wl_1_20 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2249 wl_0_25 wl_1_25 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1504 wl_0_50 wl_1_50 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1515 wl_0_53 wl_1_53 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1526 wl_0_61 wl_1_61 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1537 wl_0_50 wl_1_50 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1548 wl_0_54 wl_1_54 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1559 wl_0_56 wl_1_56 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_901 wl_0_36 wl_1_36 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_923 wl_0_40 wl_1_40 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_912 wl_0_41 wl_1_41 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4130 wl_0_94 wl_1_94 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_956 wl_0_36 wl_1_36 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_967 wl_0_37 wl_1_37 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_945 wl_0_41 wl_1_41 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_934 wl_0_44 wl_1_44 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4163 wl_0_85 wl_1_85 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4141 wl_0_87 wl_1_87 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4152 wl_0_87 wl_1_87 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_978 wl_0_33 wl_1_33 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3440 wl_0_40 wl_1_40 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3462 wl_0_44 wl_1_44 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3451 wl_0_43 wl_1_43 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_989 wl_0_45 wl_1_45 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4174 wl_0_84 wl_1_84 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4185 wl_0_91 wl_1_91 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4196 wl_0_92 wl_1_92 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2750 wl_0_17 wl_1_17 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3484 wl_0_50 wl_1_50 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3495 wl_0_59 wl_1_59 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3473 wl_0_61 wl_1_61 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2772 wl_0_24 wl_1_24 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2761 wl_0_19 wl_1_19 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2783 wl_0_16 wl_1_16 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2794 wl_0_26 wl_1_26 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7717 wl_0_70 wl_1_70 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7706 wl_0_81 wl_1_81 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7728 wl_0_122 wl_1_122 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7739 wl_0_111 wl_1_111 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_208 wl_0_27 wl_1_27 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_219 wl_0_28 wl_1_28 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2002 wl_0_7 wl_1_7 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2013 wl_0_13 wl_1_13 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2046 wl_0_12 wl_1_12 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2024 wl_0_10 wl_1_10 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2035 wl_0_5 wl_1_5 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1301 wl_0_47 wl_1_47 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2057 wl_0_14 wl_1_14 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2079 wl_0_3 wl_1_3 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2068 wl_0_3 wl_1_3 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1323 wl_0_42 wl_1_42 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1334 wl_0_46 wl_1_46 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1312 wl_0_62 wl_1_62 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1356 wl_0_33 wl_1_33 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1345 wl_0_35 wl_1_35 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1367 wl_0_42 wl_1_42 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1378 wl_0_38 wl_1_38 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1389 wl_0_44 wl_1_44 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4 wl_0_5 wl_1_5 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_742 wl_0_22 wl_1_22 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_720 wl_0_19 wl_1_19 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_731 wl_0_30 wl_1_30 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_764 wl_0_22 wl_1_22 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_775 wl_0_20 wl_1_20 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_753 wl_0_28 wl_1_28 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_797 wl_0_23 wl_1_23 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_786 wl_0_25 wl_1_25 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3270 wl_0_55 wl_1_55 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3292 wl_0_33 wl_1_33 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3281 wl_0_44 wl_1_44 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2591 wl_0_24 wl_1_24 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2580 wl_0_8 wl_1_8 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1890 wl_0_14 wl_1_14 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7525 wl_0_125 wl_1_125 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7514 wl_0_121 wl_1_121 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7503 wl_0_119 wl_1_119 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7558 wl_0_125 wl_1_125 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7536 wl_0_114 wl_1_114 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7547 wl_0_111 wl_1_111 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6813 wl_0_107 wl_1_107 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6802 wl_0_104 wl_1_104 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7569 wl_0_114 wl_1_114 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6824 wl_0_110 wl_1_110 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6835 wl_0_103 wl_1_103 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6846 wl_0_104 wl_1_104 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6868 wl_0_107 wl_1_107 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6857 wl_0_103 wl_1_103 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6879 wl_0_98 wl_1_98 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_32 wl_0_1 wl_1_1 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_21 wl_0_0 wl_1_0 bl_0_58 bl_1_58 br_0_58 br_1_58
+ sky130_fd_bd_sram__openram_dp_cell_21/a_38_n79# vdd_uq382 gnd sky130_fd_bd_sram__openram_dp_cell_21/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_10 wl_0_0 wl_1_0 bl_0_61 bl_1_61 br_0_61 br_1_61
+ sky130_fd_bd_sram__openram_dp_cell_10/a_38_n79# vdd_uq190 gnd sky130_fd_bd_sram__openram_dp_cell_10/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_54 wl_0_11 wl_1_11 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_43 wl_0_12 wl_1_12 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_65 wl_0_8 wl_1_8 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_76 wl_0_14 wl_1_14 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_98 wl_0_1 wl_1_1 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_87 wl_0_3 wl_1_3 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1131 wl_0_52 wl_1_52 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1120 wl_0_53 wl_1_53 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1142 wl_0_61 wl_1_61 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1153 wl_0_49 wl_1_49 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1175 wl_0_54 wl_1_54 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1164 wl_0_60 wl_1_60 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1186 wl_0_59 wl_1_59 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1197 wl_0_56 wl_1_56 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_550 wl_0_7 wl_1_7 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_572 wl_0_10 wl_1_10 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_561 wl_0_5 wl_1_5 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_583 wl_0_5 wl_1_5 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_594 wl_0_14 wl_1_14 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6109 wl_0_94 wl_1_94 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5419 wl_0_114 wl_1_114 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5408 wl_0_102 wl_1_102 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4729 wl_0_69 wl_1_69 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4718 wl_0_80 wl_1_80 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4707 wl_0_89 wl_1_89 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8001 wl_0_0 wl_1_0 bl_0_32 bl_1_32 br_0_32 br_1_32
+ sky130_fd_bd_sram__openram_dp_cell_8001/a_38_n79# vdd_uq2046 gnd sky130_fd_bd_sram__openram_dp_cell_8001/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8012 wl_0_117 wl_1_117 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8023 wl_0_106 wl_1_106 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7300 wl_0_105 wl_1_105 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8045 wl_0_84 wl_1_84 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8034 wl_0_95 wl_1_95 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7311 wl_0_108 wl_1_108 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7333 wl_0_106 wl_1_106 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7322 wl_0_97 wl_1_97 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8078 wl_0_51 wl_1_51 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8067 wl_0_62 wl_1_62 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8056 wl_0_73 wl_1_73 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7366 wl_0_123 wl_1_123 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7355 wl_0_115 wl_1_115 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7344 wl_0_110 wl_1_110 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8089 wl_0_40 wl_1_40 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6610 wl_0_86 wl_1_86 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6621 wl_0_88 wl_1_88 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7377 wl_0_124 wl_1_124 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7399 wl_0_121 wl_1_121 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7388 wl_0_115 wl_1_115 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5920 wl_0_66 wl_1_66 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6654 wl_0_80 wl_1_80 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6632 wl_0_90 wl_1_90 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6665 wl_0_93 wl_1_93 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6643 wl_0_94 wl_1_94 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5953 wl_0_68 wl_1_68 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6687 wl_0_71 wl_1_71 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5942 wl_0_75 wl_1_75 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5931 wl_0_75 wl_1_75 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6698 wl_0_80 wl_1_80 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6676 wl_0_82 wl_1_82 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5986 wl_0_65 wl_1_65 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5975 wl_0_66 wl_1_66 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5964 wl_0_77 wl_1_77 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5997 wl_0_66 wl_1_66 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_391 wl_0_18 wl_1_18 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_380 wl_0_27 wl_1_27 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5216 wl_0_121 wl_1_121 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5205 wl_0_101 wl_1_101 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5227 wl_0_110 wl_1_110 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5238 wl_0_99 wl_1_99 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5249 wl_0_98 wl_1_98 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4504 wl_0_74 wl_1_74 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4537 wl_0_81 wl_1_81 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4515 wl_0_91 wl_1_91 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4526 wl_0_92 wl_1_92 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3836 wl_0_21 wl_1_21 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3825 wl_0_30 wl_1_30 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3814 wl_0_41 wl_1_41 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3803 wl_0_52 wl_1_52 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4548 wl_0_88 wl_1_88 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4559 wl_0_91 wl_1_91 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3847 wl_0_10 wl_1_10 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3869 wl_0_31 wl_1_31 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3858 wl_0_32 wl_1_32 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7141 wl_0_112 wl_1_112 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7130 wl_0_105 wl_1_105 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7152 wl_0_111 wl_1_111 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7163 wl_0_105 wl_1_105 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7174 wl_0_99 wl_1_99 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6440 wl_0_78 wl_1_78 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7196 wl_0_109 wl_1_109 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7185 wl_0_105 wl_1_105 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6451 wl_0_72 wl_1_72 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6473 wl_0_72 wl_1_72 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6462 wl_0_74 wl_1_74 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5761 wl_0_79 wl_1_79 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6495 wl_0_81 wl_1_81 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5750 wl_0_90 wl_1_90 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6484 wl_0_92 wl_1_92 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5783 wl_0_122 wl_1_122 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5794 wl_0_111 wl_1_111 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5772 wl_0_68 wl_1_68 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2409 wl_0_5 wl_1_5 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1708 wl_0_61 wl_1_61 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1719 wl_0_50 wl_1_50 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5013 wl_0_127 wl_1_127 bl_0_5 bl_1_5 br_0_5 br_1_5
+ sky130_fd_bd_sram__openram_dp_cell_5013/a_38_n79# vdd_uq3774 gnd sky130_fd_bd_sram__openram_dp_cell_5013/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5024 wl_0_126 wl_1_126 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5002 wl_0_124 wl_1_124 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5046 wl_0_119 wl_1_119 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5057 wl_0_119 wl_1_119 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5035 wl_0_115 wl_1_115 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4312 wl_0_74 wl_1_74 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4301 wl_0_85 wl_1_85 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5079 wl_0_123 wl_1_123 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5068 wl_0_114 wl_1_114 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3600 wl_0_54 wl_1_54 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3611 wl_0_59 wl_1_59 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4334 wl_0_73 wl_1_73 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4345 wl_0_78 wl_1_78 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4323 wl_0_79 wl_1_79 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3644 wl_0_38 wl_1_38 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3633 wl_0_53 wl_1_53 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3622 wl_0_54 wl_1_54 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4378 wl_0_69 wl_1_69 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4389 wl_0_69 wl_1_69 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4367 wl_0_76 wl_1_76 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4356 wl_0_78 wl_1_78 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2921 wl_0_37 wl_1_37 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2910 wl_0_39 wl_1_39 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2932 wl_0_46 wl_1_46 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3655 wl_0_47 wl_1_47 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3666 wl_0_48 wl_1_48 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3677 wl_0_57 wl_1_57 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2976 wl_0_33 wl_1_33 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2965 wl_0_33 wl_1_33 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3699 wl_0_35 wl_1_35 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2943 wl_0_38 wl_1_38 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2954 wl_0_44 wl_1_44 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3688 wl_0_46 wl_1_46 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2998 wl_0_36 wl_1_36 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2987 wl_0_37 wl_1_37 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6281 wl_0_76 wl_1_76 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6270 wl_0_87 wl_1_87 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5580 wl_0_114 wl_1_114 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6292 wl_0_65 wl_1_65 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5591 wl_0_112 wl_1_112 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4890 wl_0_102 wl_1_102 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2206 wl_0_23 wl_1_23 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2228 wl_0_22 wl_1_22 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2217 wl_0_18 wl_1_18 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2239 wl_0_22 wl_1_22 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1505 wl_0_49 wl_1_49 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1516 wl_0_52 wl_1_52 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1538 wl_0_49 wl_1_49 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1549 wl_0_53 wl_1_53 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1527 wl_0_60 wl_1_60 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_913 wl_0_35 wl_1_35 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_902 wl_0_40 wl_1_40 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_924 wl_0_39 wl_1_39 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4120 wl_0_88 wl_1_88 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_957 wl_0_35 wl_1_35 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_935 wl_0_43 wl_1_43 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_946 wl_0_46 wl_1_46 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4164 wl_0_84 wl_1_84 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4142 wl_0_86 wl_1_86 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4153 wl_0_86 wl_1_86 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4131 wl_0_93 wl_1_93 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_968 wl_0_36 wl_1_36 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3441 wl_0_39 wl_1_39 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_979 wl_0_40 wl_1_40 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3430 wl_0_42 wl_1_42 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3452 wl_0_42 wl_1_42 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4175 wl_0_83 wl_1_83 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4186 wl_0_90 wl_1_90 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4197 wl_0_91 wl_1_91 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2751 wl_0_29 wl_1_29 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2740 wl_0_30 wl_1_30 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3463 wl_0_43 wl_1_43 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3485 wl_0_49 wl_1_49 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3474 wl_0_60 wl_1_60 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2773 wl_0_23 wl_1_23 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2762 wl_0_18 wl_1_18 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2784 wl_0_15 wl_1_15 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3496 wl_0_54 wl_1_54 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2795 wl_0_25 wl_1_25 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7707 wl_0_80 wl_1_80 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7729 wl_0_121 wl_1_121 bl_0_47 bl_1_47 br_0_47
+ br_1_47 bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7718 wl_0_69 wl_1_69 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_209 wl_0_26 wl_1_26 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2003 wl_0_6 wl_1_6 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2014 wl_0_12 wl_1_12 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2025 wl_0_9 wl_1_9 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2036 wl_0_4 wl_1_4 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2058 wl_0_13 wl_1_13 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2047 wl_0_11 wl_1_11 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2069 wl_0_2 wl_1_2 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1324 wl_0_41 wl_1_41 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1335 wl_0_45 wl_1_45 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1302 wl_0_48 wl_1_48 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1313 wl_0_61 wl_1_61 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1346 wl_0_34 wl_1_34 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1368 wl_0_41 wl_1_41 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1357 wl_0_46 wl_1_46 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1379 wl_0_37 wl_1_37 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5 wl_0_6 wl_1_6 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_721 wl_0_19 wl_1_19 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_710 wl_0_25 wl_1_25 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_732 wl_0_29 wl_1_29 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_765 wl_0_21 wl_1_21 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_743 wl_0_21 wl_1_21 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_754 wl_0_27 wl_1_27 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_798 wl_0_22 wl_1_22 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_776 wl_0_19 wl_1_19 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_787 wl_0_24 wl_1_24 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3260 wl_0_47 wl_1_47 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3282 wl_0_43 wl_1_43 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3293 wl_0_48 wl_1_48 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3271 wl_0_54 wl_1_54 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2592 wl_0_19 wl_1_19 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2570 wl_0_11 wl_1_11 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2581 wl_0_7 wl_1_7 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1891 wl_0_13 wl_1_13 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1880 wl_0_24 wl_1_24 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7504 wl_0_120 wl_1_120 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7515 wl_0_120 wl_1_120 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7526 wl_0_124 wl_1_124 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7559 wl_0_124 wl_1_124 bl_0_56 bl_1_56 br_0_56
+ br_1_56 bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7537 wl_0_113 wl_1_113 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7548 wl_0_112 wl_1_112 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6814 wl_0_106 wl_1_106 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6803 wl_0_103 wl_1_103 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6825 wl_0_109 wl_1_109 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6847 wl_0_103 wl_1_103 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6836 wl_0_102 wl_1_102 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6869 wl_0_106 wl_1_106 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6858 wl_0_102 wl_1_102 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_22 wl_0_6 wl_1_6 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_11 wl_0_4 wl_1_4 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_55 wl_0_14 wl_1_14 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_44 wl_0_11 wl_1_11 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_66 wl_0_8 wl_1_8 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_33 wl_0_0 wl_1_0 bl_0_57 bl_1_57 br_0_57 br_1_57
+ sky130_fd_bd_sram__openram_dp_cell_33/a_38_n79# vdd_uq446 gnd sky130_fd_bd_sram__openram_dp_cell_33/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1110 wl_0_56 wl_1_56 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_77 wl_0_13 wl_1_13 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_99 wl_0_0 wl_1_0 bl_0_59 bl_1_59 br_0_59 br_1_59
+ sky130_fd_bd_sram__openram_dp_cell_99/a_38_n79# vdd_uq318 gnd sky130_fd_bd_sram__openram_dp_cell_99/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_88 wl_0_2 wl_1_2 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1121 wl_0_52 wl_1_52 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1143 wl_0_60 wl_1_60 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1132 wl_0_62 wl_1_62 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1154 wl_0_50 wl_1_50 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1176 wl_0_53 wl_1_53 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1165 wl_0_59 wl_1_59 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1198 wl_0_55 wl_1_55 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1187 wl_0_58 wl_1_58 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_540 wl_0_2 wl_1_2 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_573 wl_0_14 wl_1_14 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_551 wl_0_6 wl_1_6 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_562 wl_0_4 wl_1_4 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_584 wl_0_4 wl_1_4 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_595 wl_0_13 wl_1_13 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3090 wl_0_57 wl_1_57 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5409 wl_0_127 wl_1_127 bl_0_17 bl_1_17 br_0_17
+ br_1_17 sky130_fd_bd_sram__openram_dp_cell_5409/a_38_n79# vdd_uq3006 gnd sky130_fd_bd_sram__openram_dp_cell_5409/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4719 wl_0_79 wl_1_79 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4708 wl_0_88 wl_1_88 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8002 wl_0_127 wl_1_127 bl_0_31 bl_1_31 br_0_31
+ br_1_31 sky130_fd_bd_sram__openram_dp_cell_8002/a_38_n79# vdd_uq2110 gnd sky130_fd_bd_sram__openram_dp_cell_8002/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8013 wl_0_116 wl_1_116 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8024 wl_0_105 wl_1_105 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8035 wl_0_94 wl_1_94 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7312 wl_0_107 wl_1_107 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7323 wl_0_106 wl_1_106 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7301 wl_0_104 wl_1_104 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8068 wl_0_61 wl_1_61 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8057 wl_0_72 wl_1_72 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8046 wl_0_83 wl_1_83 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7345 wl_0_123 wl_1_123 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7367 wl_0_122 wl_1_122 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7356 wl_0_114 wl_1_114 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7334 wl_0_105 wl_1_105 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8079 wl_0_50 wl_1_50 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6611 wl_0_85 wl_1_85 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6600 wl_0_86 wl_1_86 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6622 wl_0_87 wl_1_87 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7378 wl_0_123 wl_1_123 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7389 wl_0_114 wl_1_114 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5910 wl_0_76 wl_1_76 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6655 wl_0_79 wl_1_79 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6633 wl_0_89 wl_1_89 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6644 wl_0_93 wl_1_93 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5921 wl_0_65 wl_1_65 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5954 wl_0_67 wl_1_67 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6688 wl_0_70 wl_1_70 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5932 wl_0_74 wl_1_74 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5943 wl_0_78 wl_1_78 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6677 wl_0_81 wl_1_81 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6666 wl_0_92 wl_1_92 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5976 wl_0_65 wl_1_65 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5987 wl_0_71 wl_1_71 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5965 wl_0_76 wl_1_76 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6699 wl_0_79 wl_1_79 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5998 wl_0_65 wl_1_65 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7890 wl_0_111 wl_1_111 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_370 wl_0_22 wl_1_22 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_392 wl_0_17 wl_1_17 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_381 wl_0_26 wl_1_26 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5206 wl_0_100 wl_1_100 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5217 wl_0_120 wl_1_120 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5228 wl_0_109 wl_1_109 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5239 wl_0_98 wl_1_98 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4505 wl_0_73 wl_1_73 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4516 wl_0_84 wl_1_84 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4538 wl_0_92 wl_1_92 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4527 wl_0_91 wl_1_91 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3826 wl_0_32 wl_1_32 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3815 wl_0_40 wl_1_40 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3804 wl_0_51 wl_1_51 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4549 wl_0_87 wl_1_87 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3837 wl_0_20 wl_1_20 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3848 wl_0_9 wl_1_9 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3859 wl_0_31 wl_1_31 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7120 wl_0_115 wl_1_115 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7142 wl_0_111 wl_1_111 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7131 wl_0_104 wl_1_104 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7153 wl_0_112 wl_1_112 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7164 wl_0_104 wl_1_104 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7175 wl_0_98 wl_1_98 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6430 wl_0_73 wl_1_73 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7197 wl_0_108 wl_1_108 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7186 wl_0_104 wl_1_104 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6452 wl_0_71 wl_1_71 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6463 wl_0_73 wl_1_73 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6441 wl_0_77 wl_1_77 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5740 wl_0_100 wl_1_100 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6474 wl_0_71 wl_1_71 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5762 wl_0_78 wl_1_78 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5751 wl_0_89 wl_1_89 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6496 wl_0_90 wl_1_90 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6485 wl_0_91 wl_1_91 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5784 wl_0_121 wl_1_121 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5795 wl_0_110 wl_1_110 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5773 wl_0_67 wl_1_67 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1709 wl_0_60 wl_1_60 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5003 wl_0_127 wl_1_127 bl_0_2 bl_1_2 br_0_2 br_1_2
+ sky130_fd_bd_sram__openram_dp_cell_5003/a_38_n79# vdd_uq3966 gnd sky130_fd_bd_sram__openram_dp_cell_5003/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5014 wl_0_126 wl_1_126 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5025 wl_0_125 wl_1_125 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5058 wl_0_119 wl_1_119 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5047 wl_0_118 wl_1_118 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5036 wl_0_114 wl_1_114 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4313 wl_0_73 wl_1_73 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4302 wl_0_84 wl_1_84 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5069 wl_0_113 wl_1_113 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3601 wl_0_53 wl_1_53 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4335 wl_0_72 wl_1_72 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4346 wl_0_77 wl_1_77 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4324 wl_0_80 wl_1_80 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2900 wl_0_34 wl_1_34 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3634 wl_0_52 wl_1_52 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3623 wl_0_53 wl_1_53 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3612 wl_0_58 wl_1_58 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4379 wl_0_68 wl_1_68 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4368 wl_0_75 wl_1_75 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4357 wl_0_77 wl_1_77 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2922 wl_0_36 wl_1_36 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3645 wl_0_37 wl_1_37 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2911 wl_0_38 wl_1_38 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2933 wl_0_45 wl_1_45 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3656 wl_0_48 wl_1_48 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3667 wl_0_47 wl_1_47 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3678 wl_0_56 wl_1_56 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2944 wl_0_36 wl_1_36 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2966 wl_0_41 wl_1_41 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2955 wl_0_43 wl_1_43 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3689 wl_0_45 wl_1_45 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2988 wl_0_36 wl_1_36 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2999 wl_0_35 wl_1_35 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2977 wl_0_46 wl_1_46 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6282 wl_0_75 wl_1_75 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6260 wl_0_80 wl_1_80 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6271 wl_0_86 wl_1_86 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5570 wl_0_124 wl_1_124 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6293 wl_0_79 wl_1_79 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5581 wl_0_113 wl_1_113 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5592 wl_0_111 wl_1_111 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4891 wl_0_101 wl_1_101 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4880 wl_0_97 wl_1_97 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2207 wl_0_22 wl_1_22 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2229 wl_0_21 wl_1_21 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2218 wl_0_17 wl_1_17 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1517 wl_0_51 wl_1_51 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1506 wl_0_62 wl_1_62 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1528 wl_0_59 wl_1_59 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1539 wl_0_62 wl_1_62 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_914 wl_0_35 wl_1_35 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_903 wl_0_39 wl_1_39 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4110 wl_0_81 wl_1_81 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4121 wl_0_87 wl_1_87 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_925 wl_0_38 wl_1_38 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_936 wl_0_42 wl_1_42 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_947 wl_0_45 wl_1_45 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_958 wl_0_46 wl_1_46 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4143 wl_0_85 wl_1_85 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4154 wl_0_85 wl_1_85 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4132 wl_0_92 wl_1_92 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_969 wl_0_35 wl_1_35 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3420 wl_0_37 wl_1_37 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3431 wl_0_41 wl_1_41 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3453 wl_0_41 wl_1_41 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3442 wl_0_42 wl_1_42 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4176 wl_0_82 wl_1_82 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4165 wl_0_83 wl_1_83 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4187 wl_0_89 wl_1_89 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2730 wl_0_21 wl_1_21 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2741 wl_0_25 wl_1_25 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3464 wl_0_46 wl_1_46 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3486 wl_0_52 wl_1_52 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3475 wl_0_59 wl_1_59 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4198 wl_0_90 wl_1_90 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2774 wl_0_22 wl_1_22 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2763 wl_0_17 wl_1_17 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2752 wl_0_28 wl_1_28 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3497 wl_0_53 wl_1_53 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2796 wl_0_24 wl_1_24 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2785 wl_0_16 wl_1_16 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6090 wl_0_94 wl_1_94 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7708 wl_0_79 wl_1_79 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7719 wl_0_68 wl_1_68 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2015 wl_0_11 wl_1_11 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2004 wl_0_9 wl_1_9 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2026 wl_0_8 wl_1_8 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2037 wl_0_3 wl_1_3 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2059 wl_0_12 wl_1_12 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2048 wl_0_10 wl_1_10 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1325 wl_0_40 wl_1_40 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1303 wl_0_47 wl_1_47 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1314 wl_0_60 wl_1_60 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1347 wl_0_33 wl_1_33 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1336 wl_0_44 wl_1_44 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1358 wl_0_45 wl_1_45 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1369 wl_0_40 wl_1_40 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6 wl_0_5 wl_1_5 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_722 wl_0_18 wl_1_18 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_711 wl_0_24 wl_1_24 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_700 wl_0_25 wl_1_25 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_733 wl_0_28 wl_1_28 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_766 wl_0_20 wl_1_20 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_744 wl_0_20 wl_1_20 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_755 wl_0_26 wl_1_26 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_777 wl_0_18 wl_1_18 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_788 wl_0_23 wl_1_23 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_799 wl_0_30 wl_1_30 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3261 wl_0_48 wl_1_48 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3250 wl_0_47 wl_1_47 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3283 wl_0_42 wl_1_42 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3294 wl_0_47 wl_1_47 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3272 wl_0_53 wl_1_53 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2571 wl_0_14 wl_1_14 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2560 wl_0_3 wl_1_3 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2593 wl_0_28 wl_1_28 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2582 wl_0_30 wl_1_30 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1881 wl_0_23 wl_1_23 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1870 wl_0_32 wl_1_32 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1892 wl_0_12 wl_1_12 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7505 wl_0_119 wl_1_119 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7516 wl_0_119 wl_1_119 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7527 wl_0_123 wl_1_123 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7538 wl_0_120 wl_1_120 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7549 wl_0_111 wl_1_111 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6804 wl_0_110 wl_1_110 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6826 wl_0_108 wl_1_108 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6815 wl_0_108 wl_1_108 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6837 wl_0_101 wl_1_101 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6848 wl_0_102 wl_1_102 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6859 wl_0_101 wl_1_101 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_12 wl_0_3 wl_1_3 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_23 wl_0_5 wl_1_5 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_56 wl_0_13 wl_1_13 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_45 wl_0_10 wl_1_10 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_34 wl_0_1 wl_1_1 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1100 wl_0_54 wl_1_54 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_78 wl_0_12 wl_1_12 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_67 wl_0_8 wl_1_8 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_89 wl_0_1 wl_1_1 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1122 wl_0_51 wl_1_51 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1111 wl_0_55 wl_1_55 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1133 wl_0_61 wl_1_61 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1177 wl_0_52 wl_1_52 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1144 wl_0_59 wl_1_59 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1155 wl_0_62 wl_1_62 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1166 wl_0_62 wl_1_62 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1199 wl_0_54 wl_1_54 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1188 wl_0_57 wl_1_57 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_530 wl_0_12 wl_1_12 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_541 wl_0_1 wl_1_1 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_574 wl_0_14 wl_1_14 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_563 wl_0_5 wl_1_5 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_552 wl_0_5 wl_1_5 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_596 wl_0_12 wl_1_12 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_585 wl_0_3 wl_1_3 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3091 wl_0_56 wl_1_56 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3080 wl_0_58 wl_1_58 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2390 wl_0_14 wl_1_14 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4709 wl_0_87 wl_1_87 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8003 wl_0_126 wl_1_126 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8014 wl_0_115 wl_1_115 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8025 wl_0_104 wl_1_104 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7313 wl_0_106 wl_1_106 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7324 wl_0_105 wl_1_105 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7302 wl_0_103 wl_1_103 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8069 wl_0_60 wl_1_60 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8058 wl_0_71 wl_1_71 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8047 wl_0_82 wl_1_82 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8036 wl_0_93 wl_1_93 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7346 wl_0_122 wl_1_122 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7357 wl_0_113 wl_1_113 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7335 wl_0_104 wl_1_104 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6612 wl_0_84 wl_1_84 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6601 wl_0_85 wl_1_85 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7379 wl_0_122 wl_1_122 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7368 wl_0_121 wl_1_121 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5900 wl_0_66 wl_1_66 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6645 wl_0_67 wl_1_67 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5911 wl_0_75 wl_1_75 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6656 wl_0_80 wl_1_80 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6623 wl_0_86 wl_1_86 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6634 wl_0_88 wl_1_88 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6689 wl_0_69 wl_1_69 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5922 wl_0_70 wl_1_70 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5933 wl_0_73 wl_1_73 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5944 wl_0_77 wl_1_77 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6678 wl_0_80 wl_1_80 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6667 wl_0_91 wl_1_91 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5977 wl_0_74 wl_1_74 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5966 wl_0_75 wl_1_75 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5955 wl_0_78 wl_1_78 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5988 wl_0_70 wl_1_70 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5999 wl_0_71 wl_1_71 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7880 wl_0_121 wl_1_121 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7891 wl_0_110 wl_1_110 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_371 wl_0_21 wl_1_21 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_360 wl_0_18 wl_1_18 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_382 wl_0_25 wl_1_25 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_393 wl_0_16 wl_1_16 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5207 wl_0_99 wl_1_99 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5218 wl_0_119 wl_1_119 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5229 wl_0_108 wl_1_108 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4506 wl_0_72 wl_1_72 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4517 wl_0_83 wl_1_83 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4528 wl_0_90 wl_1_90 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3827 wl_0_31 wl_1_31 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3816 wl_0_39 wl_1_39 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3805 wl_0_50 wl_1_50 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4539 wl_0_91 wl_1_91 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3838 wl_0_19 wl_1_19 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3849 wl_0_8 wl_1_8 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7110 wl_0_125 wl_1_125 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7121 wl_0_114 wl_1_114 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7132 wl_0_103 wl_1_103 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7154 wl_0_111 wl_1_111 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7143 wl_0_112 wl_1_112 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7165 wl_0_103 wl_1_103 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6431 wl_0_70 wl_1_70 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6420 wl_0_77 wl_1_77 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7198 wl_0_107 wl_1_107 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7187 wl_0_103 wl_1_103 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7176 wl_0_97 wl_1_97 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6464 wl_0_72 wl_1_72 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6442 wl_0_76 wl_1_76 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6453 wl_0_78 wl_1_78 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5730 wl_0_110 wl_1_110 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5741 wl_0_99 wl_1_99 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6475 wl_0_70 wl_1_70 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5752 wl_0_88 wl_1_88 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6497 wl_0_89 wl_1_89 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6486 wl_0_90 wl_1_90 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5785 wl_0_120 wl_1_120 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5796 wl_0_109 wl_1_109 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5774 wl_0_66 wl_1_66 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5763 wl_0_77 wl_1_77 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_190 wl_0_14 wl_1_14 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5004 wl_0_126 wl_1_126 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5015 wl_0_121 wl_1_121 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5026 wl_0_124 wl_1_124 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5048 wl_0_117 wl_1_117 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5037 wl_0_113 wl_1_113 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4303 wl_0_83 wl_1_83 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5059 wl_0_119 wl_1_119 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3602 wl_0_52 wl_1_52 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4336 wl_0_71 wl_1_71 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4314 wl_0_72 wl_1_72 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4325 wl_0_80 wl_1_80 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3635 wl_0_51 wl_1_51 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3613 wl_0_57 wl_1_57 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3624 wl_0_62 wl_1_62 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4369 wl_0_74 wl_1_74 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4347 wl_0_76 wl_1_76 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4358 wl_0_76 wl_1_76 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2901 wl_0_33 wl_1_33 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3646 wl_0_36 wl_1_36 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2923 wl_0_37 wl_1_37 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2912 wl_0_43 wl_1_43 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3657 wl_0_47 wl_1_47 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3668 wl_0_48 wl_1_48 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2945 wl_0_35 wl_1_35 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2967 wl_0_40 wl_1_40 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2956 wl_0_42 wl_1_42 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2934 wl_0_46 wl_1_46 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3679 wl_0_55 wl_1_55 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2989 wl_0_35 wl_1_35 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2978 wl_0_46 wl_1_46 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6250 wl_0_71 wl_1_71 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6261 wl_0_80 wl_1_80 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6272 wl_0_85 wl_1_85 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5571 wl_0_123 wl_1_123 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5560 wl_0_117 wl_1_117 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6283 wl_0_74 wl_1_74 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6294 wl_0_80 wl_1_80 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5582 wl_0_114 wl_1_114 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5593 wl_0_112 wl_1_112 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4870 wl_0_107 wl_1_107 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4881 wl_0_106 wl_1_106 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4892 wl_0_100 wl_1_100 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2208 wl_0_21 wl_1_21 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2219 wl_0_28 wl_1_28 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1507 wl_0_61 wl_1_61 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1518 wl_0_50 wl_1_50 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1529 wl_0_58 wl_1_58 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_915 wl_0_34 wl_1_34 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_904 wl_0_38 wl_1_38 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4100 wl_0_84 wl_1_84 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4111 wl_0_94 wl_1_94 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_926 wl_0_37 wl_1_37 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3410 wl_0_40 wl_1_40 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_937 wl_0_41 wl_1_41 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_948 wl_0_44 wl_1_44 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4122 wl_0_86 wl_1_86 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4155 wl_0_89 wl_1_89 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4133 wl_0_91 wl_1_91 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4144 wl_0_94 wl_1_94 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3421 wl_0_36 wl_1_36 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3432 wl_0_40 wl_1_40 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3443 wl_0_41 wl_1_41 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_959 wl_0_45 wl_1_45 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4177 wl_0_81 wl_1_81 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4166 wl_0_82 wl_1_82 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4188 wl_0_88 wl_1_88 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2742 wl_0_24 wl_1_24 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2731 wl_0_20 wl_1_20 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2720 wl_0_20 wl_1_20 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3465 wl_0_38 wl_1_38 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3454 wl_0_40 wl_1_40 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3476 wl_0_58 wl_1_58 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4199 wl_0_89 wl_1_89 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2753 wl_0_21 wl_1_21 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2775 wl_0_21 wl_1_21 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2764 wl_0_16 wl_1_16 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3498 wl_0_52 wl_1_52 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3487 wl_0_51 wl_1_51 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2797 wl_0_23 wl_1_23 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2786 wl_0_15 wl_1_15 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6080 wl_0_85 wl_1_85 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6091 wl_0_93 wl_1_93 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5390 wl_0_101 wl_1_101 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7709 wl_0_78 wl_1_78 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2016 wl_0_10 wl_1_10 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2005 wl_0_8 wl_1_8 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2027 wl_0_7 wl_1_7 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2049 wl_0_14 wl_1_14 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2038 wl_0_2 wl_1_2 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1326 wl_0_39 wl_1_39 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1304 wl_0_48 wl_1_48 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1315 wl_0_59 wl_1_59 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1348 wl_0_35 wl_1_35 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1359 wl_0_44 wl_1_44 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1337 wl_0_43 wl_1_43 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7 wl_0_4 wl_1_4 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_723 wl_0_17 wl_1_17 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_712 wl_0_23 wl_1_23 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_701 wl_0_24 wl_1_24 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_745 wl_0_19 wl_1_19 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_756 wl_0_25 wl_1_25 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_734 wl_0_27 wl_1_27 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_789 wl_0_22 wl_1_22 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_767 wl_0_19 wl_1_19 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_778 wl_0_17 wl_1_17 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3240 wl_0_41 wl_1_41 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3251 wl_0_48 wl_1_48 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2550 wl_0_7 wl_1_7 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3284 wl_0_41 wl_1_41 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3295 wl_0_48 wl_1_48 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3262 wl_0_47 wl_1_47 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3273 wl_0_52 wl_1_52 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2572 wl_0_13 wl_1_13 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2561 wl_0_2 wl_1_2 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2583 wl_0_29 wl_1_29 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1882 wl_0_22 wl_1_22 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2594 wl_0_27 wl_1_27 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1871 wl_0_31 wl_1_31 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1860 wl_0_42 wl_1_42 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1893 wl_0_11 wl_1_11 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7506 wl_0_120 wl_1_120 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7528 wl_0_122 wl_1_122 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7539 wl_0_119 wl_1_119 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7517 wl_0_118 wl_1_118 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6805 wl_0_109 wl_1_109 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6827 wl_0_107 wl_1_107 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6816 wl_0_107 wl_1_107 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6838 wl_0_100 wl_1_100 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6849 wl_0_101 wl_1_101 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_13 wl_0_2 wl_1_2 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_35 wl_0_14 wl_1_14 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_57 wl_0_12 wl_1_12 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_46 wl_0_9 wl_1_9 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_24 wl_0_4 wl_1_4 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1101 wl_0_50 wl_1_50 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_79 wl_0_11 wl_1_11 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_68 wl_0_7 wl_1_7 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1123 wl_0_54 wl_1_54 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1134 wl_0_60 wl_1_60 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1112 wl_0_61 wl_1_61 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1145 wl_0_58 wl_1_58 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1156 wl_0_61 wl_1_61 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1167 wl_0_61 wl_1_61 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1178 wl_0_51 wl_1_51 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1189 wl_0_56 wl_1_56 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_520 wl_0_13 wl_1_13 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_531 wl_0_11 wl_1_11 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_575 wl_0_13 wl_1_13 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_542 wl_0_0 wl_1_0 bl_0_46 bl_1_46 br_0_46 br_1_46
+ sky130_fd_bd_sram__openram_dp_cell_542/a_38_n79# vdd_uq1150 gnd sky130_fd_bd_sram__openram_dp_cell_542/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_564 wl_0_4 wl_1_4 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_553 wl_0_4 wl_1_4 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_597 wl_0_11 wl_1_11 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_586 wl_0_2 wl_1_2 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3070 wl_0_61 wl_1_61 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3092 wl_0_55 wl_1_55 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3081 wl_0_57 wl_1_57 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2380 wl_0_16 wl_1_16 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2391 wl_0_13 wl_1_13 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1690 wl_0_47 wl_1_47 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8004 wl_0_125 wl_1_125 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8015 wl_0_114 wl_1_114 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8026 wl_0_103 wl_1_103 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7314 wl_0_105 wl_1_105 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7303 wl_0_102 wl_1_102 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8059 wl_0_70 wl_1_70 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8048 wl_0_81 wl_1_81 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8037 wl_0_92 wl_1_92 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7358 wl_0_125 wl_1_125 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7347 wl_0_121 wl_1_121 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7336 wl_0_103 wl_1_103 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7325 wl_0_102 wl_1_102 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6613 wl_0_83 wl_1_83 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6602 wl_0_94 wl_1_94 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7369 wl_0_114 wl_1_114 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5901 wl_0_65 wl_1_65 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6646 wl_0_66 wl_1_66 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6624 wl_0_85 wl_1_85 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6635 wl_0_87 wl_1_87 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5923 wl_0_69 wl_1_69 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5934 wl_0_72 wl_1_72 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5912 wl_0_74 wl_1_74 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5945 wl_0_76 wl_1_76 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6657 wl_0_79 wl_1_79 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6679 wl_0_79 wl_1_79 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6668 wl_0_90 wl_1_90 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5978 wl_0_73 wl_1_73 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5967 wl_0_74 wl_1_74 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5956 wl_0_77 wl_1_77 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5989 wl_0_69 wl_1_69 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7870 wl_0_64 wl_1_64 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7881 wl_0_120 wl_1_120 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7892 wl_0_109 wl_1_109 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_350 wl_0_21 wl_1_21 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_372 wl_0_20 wl_1_20 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_361 wl_0_17 wl_1_17 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_383 wl_0_24 wl_1_24 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_394 wl_0_15 wl_1_15 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5219 wl_0_118 wl_1_118 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5208 wl_0_98 wl_1_98 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4507 wl_0_71 wl_1_71 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4518 wl_0_82 wl_1_82 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4529 wl_0_89 wl_1_89 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3817 wl_0_38 wl_1_38 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3806 wl_0_49 wl_1_49 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3839 wl_0_18 wl_1_18 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3828 wl_0_29 wl_1_29 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7111 wl_0_124 wl_1_124 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7122 wl_0_113 wl_1_113 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7100 wl_0_104 wl_1_104 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7133 wl_0_102 wl_1_102 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7144 wl_0_111 wl_1_111 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7155 wl_0_112 wl_1_112 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7166 wl_0_102 wl_1_102 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6410 wl_0_72 wl_1_72 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6421 wl_0_76 wl_1_76 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5720 wl_0_120 wl_1_120 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7199 wl_0_106 wl_1_106 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7188 wl_0_102 wl_1_102 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7177 wl_0_101 wl_1_101 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6432 wl_0_69 wl_1_69 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6443 wl_0_75 wl_1_75 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6454 wl_0_77 wl_1_77 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5731 wl_0_109 wl_1_109 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5742 wl_0_98 wl_1_98 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6476 wl_0_69 wl_1_69 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6465 wl_0_71 wl_1_71 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5753 wl_0_87 wl_1_87 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6487 wl_0_89 wl_1_89 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6498 wl_0_94 wl_1_94 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5786 wl_0_119 wl_1_119 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5775 wl_0_65 wl_1_65 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5764 wl_0_76 wl_1_76 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5797 wl_0_108 wl_1_108 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_191 wl_0_13 wl_1_13 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_180 wl_0_0 wl_1_0 bl_0_50 bl_1_50 br_0_50 br_1_50
+ sky130_fd_bd_sram__openram_dp_cell_180/a_38_n79# vdd_uq894 gnd sky130_fd_bd_sram__openram_dp_cell_180/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5005 wl_0_125 wl_1_125 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5038 wl_0_127 wl_1_127 bl_0_3 bl_1_3 br_0_3 br_1_3
+ sky130_fd_bd_sram__openram_dp_cell_5038/a_38_n79# vdd_uq3902 gnd sky130_fd_bd_sram__openram_dp_cell_5038/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5016 wl_0_124 wl_1_124 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5027 wl_0_123 wl_1_123 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5049 wl_0_116 wl_1_116 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4304 wl_0_82 wl_1_82 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4326 wl_0_69 wl_1_69 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4337 wl_0_70 wl_1_70 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4315 wl_0_71 wl_1_71 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3603 wl_0_51 wl_1_51 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3614 wl_0_56 wl_1_56 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3625 wl_0_61 wl_1_61 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4359 wl_0_75 wl_1_75 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4348 wl_0_78 wl_1_78 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2913 wl_0_35 wl_1_35 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2924 wl_0_36 wl_1_36 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3647 wl_0_35 wl_1_35 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2902 wl_0_40 wl_1_40 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3669 wl_0_47 wl_1_47 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3658 wl_0_48 wl_1_48 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3636 wl_0_50 wl_1_50 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2946 wl_0_34 wl_1_34 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2957 wl_0_41 wl_1_41 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2935 wl_0_45 wl_1_45 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2968 wl_0_39 wl_1_39 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2979 wl_0_45 wl_1_45 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6251 wl_0_70 wl_1_70 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6262 wl_0_79 wl_1_79 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6240 wl_0_81 wl_1_81 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6273 wl_0_84 wl_1_84 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5550 wl_0_127 wl_1_127 bl_0_27 bl_1_27 br_0_27
+ br_1_27 sky130_fd_bd_sram__openram_dp_cell_5550/a_38_n79# vdd_uq2366 gnd sky130_fd_bd_sram__openram_dp_cell_5550/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5561 wl_0_116 wl_1_116 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6284 wl_0_73 wl_1_73 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6295 wl_0_79 wl_1_79 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5572 wl_0_122 wl_1_122 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5583 wl_0_113 wl_1_113 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5594 wl_0_111 wl_1_111 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4882 wl_0_110 wl_1_110 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4871 wl_0_106 wl_1_106 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4893 wl_0_99 wl_1_99 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4860 wl_0_99 wl_1_99 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2209 wl_0_20 wl_1_20 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1508 wl_0_60 wl_1_60 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1519 wl_0_49 wl_1_49 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_905 wl_0_37 wl_1_37 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4101 wl_0_83 wl_1_83 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4112 wl_0_93 wl_1_93 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_916 wl_0_33 wl_1_33 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_927 wl_0_36 wl_1_36 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_938 wl_0_40 wl_1_40 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3400 wl_0_43 wl_1_43 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_949 wl_0_43 wl_1_43 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4123 wl_0_85 wl_1_85 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4145 wl_0_93 wl_1_93 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4134 wl_0_94 wl_1_94 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3422 wl_0_35 wl_1_35 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3411 wl_0_39 wl_1_39 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3444 wl_0_40 wl_1_40 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3433 wl_0_39 wl_1_39 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4167 wl_0_81 wl_1_81 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4156 wl_0_88 wl_1_88 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4178 wl_0_92 wl_1_92 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2732 wl_0_19 wl_1_19 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2721 wl_0_19 wl_1_19 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2710 wl_0_28 wl_1_28 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3466 wl_0_37 wl_1_37 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3455 wl_0_39 wl_1_39 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3477 wl_0_57 wl_1_57 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4189 wl_0_87 wl_1_87 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2743 wl_0_23 wl_1_23 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2754 wl_0_20 wl_1_20 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2765 wl_0_15 wl_1_15 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3488 wl_0_50 wl_1_50 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3499 wl_0_51 wl_1_51 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2798 wl_0_22 wl_1_22 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2776 wl_0_20 wl_1_20 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2787 wl_0_16 wl_1_16 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6070 wl_0_83 wl_1_83 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6081 wl_0_94 wl_1_94 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6092 wl_0_92 wl_1_92 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5380 wl_0_104 wl_1_104 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5391 wl_0_100 wl_1_100 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4690 wl_0_80 wl_1_80 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2017 wl_0_9 wl_1_9 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2006 wl_0_7 wl_1_7 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2028 wl_0_6 wl_1_6 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2039 wl_0_1 wl_1_1 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1305 wl_0_48 wl_1_48 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1316 wl_0_58 wl_1_58 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1349 wl_0_34 wl_1_34 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1327 wl_0_38 wl_1_38 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1338 wl_0_42 wl_1_42 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8 wl_0_2 wl_1_2 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_713 wl_0_22 wl_1_22 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_724 wl_0_18 wl_1_18 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_702 wl_0_25 wl_1_25 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_746 wl_0_18 wl_1_18 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_757 wl_0_24 wl_1_24 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_735 wl_0_26 wl_1_26 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_779 wl_0_21 wl_1_21 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_768 wl_0_18 wl_1_18 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3241 wl_0_40 wl_1_40 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3252 wl_0_47 wl_1_47 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3230 wl_0_51 wl_1_51 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2540 wl_0_12 wl_1_12 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3285 wl_0_40 wl_1_40 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3274 wl_0_51 wl_1_51 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3263 wl_0_62 wl_1_62 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2584 wl_0_17 wl_1_17 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2573 wl_0_12 wl_1_12 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2551 wl_0_6 wl_1_6 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2562 wl_0_1 wl_1_1 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3296 wl_0_47 wl_1_47 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2595 wl_0_26 wl_1_26 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1872 wl_0_30 wl_1_30 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1861 wl_0_41 wl_1_41 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1850 wl_0_52 wl_1_52 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1883 wl_0_21 wl_1_21 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1894 wl_0_10 wl_1_10 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7507 wl_0_119 wl_1_119 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7529 wl_0_121 wl_1_121 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7518 wl_0_117 wl_1_117 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6806 wl_0_108 wl_1_108 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6828 wl_0_106 wl_1_106 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6817 wl_0_106 wl_1_106 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6839 wl_0_99 wl_1_99 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_14 wl_0_1 wl_1_1 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_36 wl_0_13 wl_1_13 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_47 wl_0_12 wl_1_12 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_25 wl_0_3 wl_1_3 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_58 wl_0_11 wl_1_11 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_69 wl_0_7 wl_1_7 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1124 wl_0_53 wl_1_53 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1102 wl_0_53 wl_1_53 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1113 wl_0_60 wl_1_60 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1146 wl_0_57 wl_1_57 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1135 wl_0_59 wl_1_59 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1157 wl_0_60 wl_1_60 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1168 wl_0_60 wl_1_60 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1179 wl_0_50 wl_1_50 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_521 wl_0_12 wl_1_12 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_532 wl_0_10 wl_1_10 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_510 wl_0_3 wl_1_3 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_543 wl_0_11 wl_1_11 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_565 wl_0_3 wl_1_3 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_554 wl_0_3 wl_1_3 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_587 wl_0_11 wl_1_11 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_576 wl_0_12 wl_1_12 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_598 wl_0_10 wl_1_10 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3060 wl_0_49 wl_1_49 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3093 wl_0_54 wl_1_54 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3082 wl_0_56 wl_1_56 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3071 wl_0_62 wl_1_62 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2381 wl_0_15 wl_1_15 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2392 wl_0_12 wl_1_12 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2370 wl_0_9 wl_1_9 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1680 wl_0_57 wl_1_57 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1691 wl_0_48 wl_1_48 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8005 wl_0_124 wl_1_124 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8016 wl_0_113 wl_1_113 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7315 wl_0_104 wl_1_104 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8027 wl_0_102 wl_1_102 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7304 wl_0_101 wl_1_101 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8049 wl_0_80 wl_1_80 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8038 wl_0_91 wl_1_91 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7348 wl_0_116 wl_1_116 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7337 wl_0_102 wl_1_102 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7326 wl_0_101 wl_1_101 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6603 wl_0_93 wl_1_93 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7359 wl_0_127 wl_1_127 bl_0_49 bl_1_49 br_0_49
+ br_1_49 sky130_fd_bd_sram__openram_dp_cell_7359/a_38_n79# vdd_uq958 gnd sky130_fd_bd_sram__openram_dp_cell_7359/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6647 wl_0_65 wl_1_65 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5902 wl_0_66 wl_1_66 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6614 wl_0_82 wl_1_82 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6625 wl_0_84 wl_1_84 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6636 wl_0_86 wl_1_86 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5924 wl_0_68 wl_1_68 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5935 wl_0_71 wl_1_71 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5913 wl_0_73 wl_1_73 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6658 wl_0_80 wl_1_80 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6669 wl_0_89 wl_1_89 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5968 wl_0_73 wl_1_73 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5946 wl_0_75 wl_1_75 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5957 wl_0_77 wl_1_77 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5979 wl_0_72 wl_1_72 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7871 wl_0_63 wl_1_63 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7860 wl_0_64 wl_1_64 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7882 wl_0_119 wl_1_119 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7893 wl_0_108 wl_1_108 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_340 wl_0_22 wl_1_22 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_351 wl_0_20 wl_1_20 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_373 wl_0_19 wl_1_19 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_362 wl_0_30 wl_1_30 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_395 wl_0_14 wl_1_14 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_384 wl_0_23 wl_1_23 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5209 wl_0_97 wl_1_97 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4519 wl_0_81 wl_1_81 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4508 wl_0_88 wl_1_88 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3818 wl_0_37 wl_1_37 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3807 wl_0_48 wl_1_48 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3829 wl_0_28 wl_1_28 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7112 wl_0_123 wl_1_123 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7123 wl_0_112 wl_1_112 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7101 wl_0_103 wl_1_103 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7156 wl_0_112 wl_1_112 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7145 wl_0_112 wl_1_112 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7134 wl_0_101 wl_1_101 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6400 wl_0_66 wl_1_66 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6411 wl_0_71 wl_1_71 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6422 wl_0_75 wl_1_75 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7189 wl_0_101 wl_1_101 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7167 wl_0_101 wl_1_101 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7178 wl_0_100 wl_1_100 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6455 wl_0_65 wl_1_65 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6433 wl_0_67 wl_1_67 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6444 wl_0_74 wl_1_74 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5710 wl_0_95 wl_1_95 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5721 wl_0_119 wl_1_119 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5732 wl_0_108 wl_1_108 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5743 wl_0_97 wl_1_97 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6466 wl_0_70 wl_1_70 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6477 wl_0_86 wl_1_86 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6488 wl_0_88 wl_1_88 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5787 wl_0_118 wl_1_118 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5765 wl_0_75 wl_1_75 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5754 wl_0_86 wl_1_86 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6499 wl_0_93 wl_1_93 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5776 wl_0_96 wl_1_96 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5798 wl_0_107 wl_1_107 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7690 wl_0_97 wl_1_97 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_170 wl_0_14 wl_1_14 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_181 wl_0_3 wl_1_3 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_192 wl_0_12 wl_1_12 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5006 wl_0_124 wl_1_124 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5039 wl_0_126 wl_1_126 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5028 wl_0_122 wl_1_122 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5017 wl_0_121 wl_1_121 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4327 wl_0_68 wl_1_68 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4316 wl_0_70 wl_1_70 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4305 wl_0_81 wl_1_81 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3604 wl_0_50 wl_1_50 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3615 wl_0_55 wl_1_55 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3626 wl_0_60 wl_1_60 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4338 wl_0_69 wl_1_69 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4349 wl_0_75 wl_1_75 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3648 wl_0_34 wl_1_34 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2903 wl_0_39 wl_1_39 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2914 wl_0_42 wl_1_42 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3659 wl_0_47 wl_1_47 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3637 wl_0_49 wl_1_49 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2947 wl_0_33 wl_1_33 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2925 wl_0_35 wl_1_35 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2936 wl_0_38 wl_1_38 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2958 wl_0_40 wl_1_40 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2969 wl_0_38 wl_1_38 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6230 wl_0_91 wl_1_91 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6252 wl_0_69 wl_1_69 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6241 wl_0_80 wl_1_80 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6263 wl_0_94 wl_1_94 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5551 wl_0_126 wl_1_126 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5540 wl_0_120 wl_1_120 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5562 wl_0_115 wl_1_115 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6285 wl_0_72 wl_1_72 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6296 wl_0_79 wl_1_79 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6274 wl_0_83 wl_1_83 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5584 wl_0_127 wl_1_127 bl_0_25 bl_1_25 br_0_25
+ br_1_25 sky130_fd_bd_sram__openram_dp_cell_5584/a_38_n79# vdd_uq2494 gnd sky130_fd_bd_sram__openram_dp_cell_5584/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5573 wl_0_121 wl_1_121 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5595 wl_0_112 wl_1_112 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4850 wl_0_102 wl_1_102 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4883 wl_0_109 wl_1_109 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4872 wl_0_105 wl_1_105 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4861 wl_0_98 wl_1_98 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4894 wl_0_98 wl_1_98 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1509 wl_0_59 wl_1_59 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_906 wl_0_36 wl_1_36 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4102 wl_0_82 wl_1_82 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_928 wl_0_35 wl_1_35 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_939 wl_0_39 wl_1_39 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3401 wl_0_42 wl_1_42 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_917 wl_0_46 wl_1_46 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4124 wl_0_84 wl_1_84 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4113 wl_0_92 wl_1_92 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4146 wl_0_92 wl_1_92 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4135 wl_0_93 wl_1_93 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3423 wl_0_34 wl_1_34 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3412 wl_0_38 wl_1_38 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3434 wl_0_38 wl_1_38 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4157 wl_0_87 wl_1_87 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4168 wl_0_90 wl_1_90 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4179 wl_0_91 wl_1_91 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2700 wl_0_23 wl_1_23 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2733 wl_0_18 wl_1_18 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2722 wl_0_18 wl_1_18 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2711 wl_0_26 wl_1_26 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3467 wl_0_38 wl_1_38 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3456 wl_0_38 wl_1_38 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3445 wl_0_39 wl_1_39 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2744 wl_0_22 wl_1_22 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2755 wl_0_19 wl_1_19 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2766 wl_0_30 wl_1_30 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3489 wl_0_49 wl_1_49 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3478 wl_0_56 wl_1_56 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2799 wl_0_21 wl_1_21 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2777 wl_0_19 wl_1_19 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2788 wl_0_15 wl_1_15 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6060 wl_0_89 wl_1_89 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6071 wl_0_94 wl_1_94 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5370 wl_0_105 wl_1_105 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6093 wl_0_91 wl_1_91 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6082 wl_0_93 wl_1_93 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5381 wl_0_103 wl_1_103 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5392 wl_0_99 wl_1_99 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4691 wl_0_79 wl_1_79 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4680 wl_0_84 wl_1_84 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3990 wl_0_78 wl_1_78 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2018 wl_0_8 wl_1_8 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2007 wl_0_6 wl_1_6 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2029 wl_0_5 wl_1_5 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1306 wl_0_47 wl_1_47 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1317 wl_0_57 wl_1_57 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1328 wl_0_37 wl_1_37 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1339 wl_0_41 wl_1_41 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_9 wl_0_1 wl_1_1 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_714 wl_0_21 wl_1_21 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_703 wl_0_23 wl_1_23 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_747 wl_0_19 wl_1_19 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_725 wl_0_17 wl_1_17 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_736 wl_0_28 wl_1_28 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_769 wl_0_17 wl_1_17 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_758 wl_0_23 wl_1_23 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3242 wl_0_39 wl_1_39 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3231 wl_0_50 wl_1_50 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3220 wl_0_61 wl_1_61 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2530 wl_0_13 wl_1_13 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2541 wl_0_11 wl_1_11 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3286 wl_0_39 wl_1_39 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3253 wl_0_48 wl_1_48 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3275 wl_0_50 wl_1_50 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3264 wl_0_61 wl_1_61 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2574 wl_0_11 wl_1_11 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2563 wl_0_0 wl_1_0 bl_0_3 bl_1_3 br_0_3 br_1_3
+ sky130_fd_bd_sram__openram_dp_cell_2563/a_38_n79# vdd_uq3902 gnd sky130_fd_bd_sram__openram_dp_cell_2563/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2552 wl_0_5 wl_1_5 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3297 wl_0_48 wl_1_48 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2585 wl_0_19 wl_1_19 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2596 wl_0_25 wl_1_25 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1862 wl_0_40 wl_1_40 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1851 wl_0_51 wl_1_51 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1840 wl_0_62 wl_1_62 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1884 wl_0_20 wl_1_20 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1895 wl_0_9 wl_1_9 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1873 wl_0_29 wl_1_29 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7508 wl_0_127 wl_1_127 bl_0_60 bl_1_60 br_0_60
+ br_1_60 sky130_fd_bd_sram__openram_dp_cell_7508/a_38_n79# vdd_uq254 gnd sky130_fd_bd_sram__openram_dp_cell_7508/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7519 wl_0_116 wl_1_116 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6807 wl_0_107 wl_1_107 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6818 wl_0_105 wl_1_105 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6829 wl_0_100 wl_1_100 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_48 wl_0_14 wl_1_14 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_37 wl_0_12 wl_1_12 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_15 wl_0_0 wl_1_0 bl_0_62 bl_1_62 br_0_62 br_1_62
+ sky130_fd_bd_sram__openram_dp_cell_15/a_38_n79# vdd_uq99 gnd sky130_fd_bd_sram__openram_dp_cell_15/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_26 wl_0_2 wl_1_2 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_59 wl_0_10 wl_1_10 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1125 wl_0_52 wl_1_52 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1114 wl_0_59 wl_1_59 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1103 wl_0_62 wl_1_62 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1147 wl_0_56 wl_1_56 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1136 wl_0_58 wl_1_58 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1158 wl_0_59 wl_1_59 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1169 wl_0_59 wl_1_59 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_500 wl_0_11 wl_1_11 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_522 wl_0_8 wl_1_8 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_511 wl_0_2 wl_1_2 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_555 wl_0_11 wl_1_11 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_544 wl_0_10 wl_1_10 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_533 wl_0_9 wl_1_9 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_566 wl_0_2 wl_1_2 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_577 wl_0_11 wl_1_11 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_588 wl_0_10 wl_1_10 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_599 wl_0_9 wl_1_9 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3050 wl_0_50 wl_1_50 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3061 wl_0_51 wl_1_51 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3094 wl_0_53 wl_1_53 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3083 wl_0_55 wl_1_55 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3072 wl_0_61 wl_1_61 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2360 wl_0_17 wl_1_17 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2382 wl_0_16 wl_1_16 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2371 wl_0_8 wl_1_8 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2393 wl_0_11 wl_1_11 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1670 wl_0_51 wl_1_51 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1681 wl_0_56 wl_1_56 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1692 wl_0_47 wl_1_47 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8006 wl_0_123 wl_1_123 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8017 wl_0_112 wl_1_112 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8028 wl_0_101 wl_1_101 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7305 wl_0_100 wl_1_100 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8039 wl_0_90 wl_1_90 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7349 wl_0_115 wl_1_115 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7316 wl_0_103 wl_1_103 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7338 wl_0_101 wl_1_101 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7327 wl_0_99 wl_1_99 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6604 wl_0_92 wl_1_92 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6615 wl_0_81 wl_1_81 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6626 wl_0_83 wl_1_83 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6637 wl_0_85 wl_1_85 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5903 wl_0_65 wl_1_65 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5936 wl_0_70 wl_1_70 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5914 wl_0_72 wl_1_72 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5925 wl_0_78 wl_1_78 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6648 wl_0_80 wl_1_80 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6659 wl_0_79 wl_1_79 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5969 wl_0_72 wl_1_72 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5947 wl_0_74 wl_1_74 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5958 wl_0_76 wl_1_76 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7861 wl_0_63 wl_1_63 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7850 wl_0_64 wl_1_64 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7883 wl_0_118 wl_1_118 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7894 wl_0_107 wl_1_107 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7872 wl_0_64 wl_1_64 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_330 wl_0_18 wl_1_18 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_352 wl_0_19 wl_1_19 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_374 wl_0_18 wl_1_18 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_363 wl_0_29 wl_1_29 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_341 wl_0_30 wl_1_30 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_385 wl_0_22 wl_1_22 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_396 wl_0_13 wl_1_13 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2190 wl_0_21 wl_1_21 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4509 wl_0_87 wl_1_87 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3808 wl_0_47 wl_1_47 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3819 wl_0_36 wl_1_36 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7113 wl_0_122 wl_1_122 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7124 wl_0_111 wl_1_111 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7102 wl_0_102 wl_1_102 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7157 wl_0_111 wl_1_111 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7146 wl_0_111 wl_1_111 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7135 wl_0_100 wl_1_100 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6401 wl_0_65 wl_1_65 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6412 wl_0_70 wl_1_70 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7168 wl_0_100 wl_1_100 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7179 wl_0_99 wl_1_99 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6434 wl_0_65 wl_1_65 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6445 wl_0_73 wl_1_73 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6423 wl_0_74 wl_1_74 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5711 wl_0_96 wl_1_96 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5700 wl_0_95 wl_1_95 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5722 wl_0_118 wl_1_118 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5733 wl_0_107 wl_1_107 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6456 wl_0_78 wl_1_78 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6467 wl_0_78 wl_1_78 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6478 wl_0_85 wl_1_85 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6489 wl_0_87 wl_1_87 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5744 wl_0_96 wl_1_96 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5766 wl_0_74 wl_1_74 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5755 wl_0_85 wl_1_85 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5777 wl_0_95 wl_1_95 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5788 wl_0_117 wl_1_117 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5799 wl_0_106 wl_1_106 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7680 wl_0_107 wl_1_107 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7691 wl_0_96 wl_1_96 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6990 wl_0_123 wl_1_123 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_171 wl_0_13 wl_1_13 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_160 wl_0_6 wl_1_6 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_182 wl_0_2 wl_1_2 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_193 wl_0_11 wl_1_11 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5018 wl_0_127 wl_1_127 bl_0_6 bl_1_6 br_0_6 br_1_6
+ sky130_fd_bd_sram__openram_dp_cell_5018/a_38_n79# vdd_uq3710 gnd sky130_fd_bd_sram__openram_dp_cell_5018/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5007 wl_0_123 wl_1_123 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5029 wl_0_121 wl_1_121 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4328 wl_0_67 wl_1_67 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4317 wl_0_69 wl_1_69 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4306 wl_0_80 wl_1_80 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3605 wl_0_49 wl_1_49 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3616 wl_0_54 wl_1_54 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4339 wl_0_68 wl_1_68 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3649 wl_0_33 wl_1_33 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2915 wl_0_34 wl_1_34 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2904 wl_0_38 wl_1_38 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3638 wl_0_42 wl_1_42 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3627 wl_0_59 wl_1_59 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2926 wl_0_34 wl_1_34 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2948 wl_0_37 wl_1_37 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2937 wl_0_37 wl_1_37 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2959 wl_0_39 wl_1_39 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6220 wl_0_93 wl_1_93 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6253 wl_0_68 wl_1_68 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6242 wl_0_79 wl_1_79 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6231 wl_0_90 wl_1_90 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6264 wl_0_93 wl_1_93 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5552 wl_0_125 wl_1_125 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5541 wl_0_119 wl_1_119 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5530 wl_0_113 wl_1_113 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6286 wl_0_71 wl_1_71 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6297 wl_0_80 wl_1_80 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6275 wl_0_82 wl_1_82 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5585 wl_0_126 wl_1_126 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5574 wl_0_120 wl_1_120 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5563 wl_0_114 wl_1_114 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4840 wl_0_110 wl_1_110 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5596 wl_0_111 wl_1_111 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4884 wl_0_108 wl_1_108 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4873 wl_0_104 wl_1_104 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4851 wl_0_101 wl_1_101 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4862 wl_0_97 wl_1_97 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4895 wl_0_97 wl_1_97 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4103 wl_0_81 wl_1_81 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_929 wl_0_34 wl_1_34 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_918 wl_0_45 wl_1_45 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_907 wl_0_46 wl_1_46 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4125 wl_0_83 wl_1_83 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4136 wl_0_92 wl_1_92 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4114 wl_0_94 wl_1_94 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3424 wl_0_33 wl_1_33 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3413 wl_0_37 wl_1_37 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3435 wl_0_37 wl_1_37 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3402 wl_0_41 wl_1_41 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4169 wl_0_89 wl_1_89 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4158 wl_0_90 wl_1_90 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4147 wl_0_91 wl_1_91 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2701 wl_0_22 wl_1_22 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2712 wl_0_25 wl_1_25 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2723 wl_0_30 wl_1_30 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3468 wl_0_37 wl_1_37 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3457 wl_0_37 wl_1_37 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3446 wl_0_46 wl_1_46 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2745 wl_0_21 wl_1_21 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2756 wl_0_18 wl_1_18 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2734 wl_0_17 wl_1_17 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3479 wl_0_55 wl_1_55 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2778 wl_0_18 wl_1_18 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2789 wl_0_16 wl_1_16 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2767 wl_0_29 wl_1_29 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6061 wl_0_84 wl_1_84 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6050 wl_0_88 wl_1_88 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6072 wl_0_93 wl_1_93 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5360 wl_0_105 wl_1_105 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6094 wl_0_90 wl_1_90 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6083 wl_0_92 wl_1_92 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5371 wl_0_104 wl_1_104 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5382 wl_0_102 wl_1_102 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5393 wl_0_98 wl_1_98 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4692 wl_0_80 wl_1_80 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4681 wl_0_83 wl_1_83 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4670 wl_0_94 wl_1_94 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3980 wl_0_76 wl_1_76 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3991 wl_0_77 wl_1_77 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2019 wl_0_7 wl_1_7 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2008 wl_0_5 wl_1_5 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1307 wl_0_47 wl_1_47 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1329 wl_0_36 wl_1_36 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1318 wl_0_56 wl_1_56 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_704 wl_0_22 wl_1_22 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_715 wl_0_20 wl_1_20 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_748 wl_0_18 wl_1_18 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_726 wl_0_24 wl_1_24 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_737 wl_0_27 wl_1_27 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_759 wl_0_22 wl_1_22 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3243 wl_0_38 wl_1_38 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3232 wl_0_49 wl_1_49 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3210 wl_0_52 wl_1_52 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3221 wl_0_60 wl_1_60 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2520 wl_0_14 wl_1_14 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2531 wl_0_12 wl_1_12 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3254 wl_0_47 wl_1_47 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3276 wl_0_49 wl_1_49 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3265 wl_0_60 wl_1_60 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2575 wl_0_10 wl_1_10 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2564 wl_0_8 wl_1_8 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2542 wl_0_6 wl_1_6 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2553 wl_0_4 wl_1_4 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1830 wl_0_5 wl_1_5 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3287 wl_0_38 wl_1_38 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3298 wl_0_47 wl_1_47 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2586 wl_0_29 wl_1_29 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2597 wl_0_30 wl_1_30 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1863 wl_0_39 wl_1_39 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1852 wl_0_50 wl_1_50 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1841 wl_0_61 wl_1_61 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1885 wl_0_19 wl_1_19 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1896 wl_0_8 wl_1_8 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1874 wl_0_28 wl_1_28 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5190 wl_0_114 wl_1_114 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7509 wl_0_126 wl_1_126 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6808 wl_0_106 wl_1_106 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6819 wl_0_104 wl_1_104 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_38 wl_0_11 wl_1_11 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_16 wl_0_6 wl_1_6 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_27 wl_0_6 wl_1_6 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_49 wl_0_13 wl_1_13 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1115 wl_0_58 wl_1_58 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1104 wl_0_62 wl_1_62 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1126 wl_0_51 wl_1_51 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1148 wl_0_55 wl_1_55 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1137 wl_0_57 wl_1_57 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1159 wl_0_58 wl_1_58 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_512 wl_0_14 wl_1_14 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_501 wl_0_10 wl_1_10 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_523 wl_0_7 wl_1_7 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_545 wl_0_12 wl_1_12 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_556 wl_0_10 wl_1_10 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_534 wl_0_8 wl_1_8 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_589 wl_0_9 wl_1_9 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_578 wl_0_7 wl_1_7 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_567 wl_0_2 wl_1_2 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3051 wl_0_49 wl_1_49 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3040 wl_0_56 wl_1_56 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3062 wl_0_54 wl_1_54 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3084 wl_0_54 wl_1_54 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3073 wl_0_60 wl_1_60 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2361 wl_0_16 wl_1_16 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2383 wl_0_15 wl_1_15 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2372 wl_0_7 wl_1_7 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2350 wl_0_27 wl_1_27 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3095 wl_0_52 wl_1_52 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2394 wl_0_10 wl_1_10 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1671 wl_0_50 wl_1_50 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1660 wl_0_61 wl_1_61 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1693 wl_0_48 wl_1_48 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1682 wl_0_55 wl_1_55 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8007 wl_0_122 wl_1_122 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8018 wl_0_111 wl_1_111 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7306 wl_0_99 wl_1_99 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8029 wl_0_100 wl_1_100 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7317 wl_0_102 wl_1_102 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7339 wl_0_100 wl_1_100 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7328 wl_0_97 wl_1_97 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6627 wl_0_82 wl_1_82 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6638 wl_0_84 wl_1_84 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6616 wl_0_84 wl_1_84 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6605 wl_0_91 wl_1_91 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5915 wl_0_71 wl_1_71 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5904 wl_0_74 wl_1_74 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5926 wl_0_77 wl_1_77 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6649 wl_0_79 wl_1_79 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5937 wl_0_69 wl_1_69 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5948 wl_0_73 wl_1_73 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5959 wl_0_75 wl_1_75 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7862 wl_0_64 wl_1_64 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7851 wl_0_63 wl_1_63 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7840 wl_0_64 wl_1_64 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7884 wl_0_117 wl_1_117 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7895 wl_0_106 wl_1_106 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7873 wl_0_63 wl_1_63 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_331 wl_0_17 wl_1_17 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_320 wl_0_28 wl_1_28 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_353 wl_0_18 wl_1_18 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_364 wl_0_28 wl_1_28 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_342 wl_0_29 wl_1_29 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_386 wl_0_21 wl_1_21 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_375 wl_0_17 wl_1_17 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_397 wl_0_12 wl_1_12 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2191 wl_0_20 wl_1_20 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2180 wl_0_28 wl_1_28 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1490 wl_0_46 wl_1_46 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3809 wl_0_46 wl_1_46 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7114 wl_0_121 wl_1_121 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7103 wl_0_101 wl_1_101 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7147 wl_0_112 wl_1_112 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7125 wl_0_110 wl_1_110 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7136 wl_0_99 wl_1_99 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6402 wl_0_68 wl_1_68 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6413 wl_0_69 wl_1_69 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7158 wl_0_111 wl_1_111 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7169 wl_0_99 wl_1_99 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6435 wl_0_69 wl_1_69 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6446 wl_0_69 wl_1_69 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6424 wl_0_73 wl_1_73 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5701 wl_0_96 wl_1_96 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5723 wl_0_117 wl_1_117 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5734 wl_0_106 wl_1_106 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6457 wl_0_77 wl_1_77 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6468 wl_0_77 wl_1_77 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6479 wl_0_83 wl_1_83 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5712 wl_0_95 wl_1_95 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5778 wl_0_127 wl_1_127 bl_0_15 bl_1_15 br_0_15
+ br_1_15 sky130_fd_bd_sram__openram_dp_cell_5778/a_38_n79# vdd_uq3134 gnd sky130_fd_bd_sram__openram_dp_cell_5778/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5767 wl_0_73 wl_1_73 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5756 wl_0_84 wl_1_84 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5745 wl_0_95 wl_1_95 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5789 wl_0_116 wl_1_116 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7670 wl_0_117 wl_1_117 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7681 wl_0_106 wl_1_106 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7692 wl_0_95 wl_1_95 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6991 wl_0_122 wl_1_122 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6980 wl_0_120 wl_1_120 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_172 wl_0_12 wl_1_12 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_150 wl_0_4 wl_1_4 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_161 wl_0_5 wl_1_5 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_194 wl_0_14 wl_1_14 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_183 wl_0_1 wl_1_1 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5019 wl_0_123 wl_1_123 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5008 wl_0_122 wl_1_122 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4318 wl_0_68 wl_1_68 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4307 wl_0_79 wl_1_79 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3617 wl_0_53 wl_1_53 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3606 wl_0_56 wl_1_56 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4329 wl_0_78 wl_1_78 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2905 wl_0_37 wl_1_37 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3639 wl_0_41 wl_1_41 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3628 wl_0_58 wl_1_58 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2916 wl_0_33 wl_1_33 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2927 wl_0_33 wl_1_33 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2938 wl_0_34 wl_1_34 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2949 wl_0_44 wl_1_44 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6210 wl_0_83 wl_1_83 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6221 wl_0_92 wl_1_92 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6254 wl_0_67 wl_1_67 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6243 wl_0_78 wl_1_78 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6232 wl_0_89 wl_1_89 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5520 wl_0_123 wl_1_123 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5553 wl_0_124 wl_1_124 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5531 wl_0_120 wl_1_120 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5542 wl_0_118 wl_1_118 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6287 wl_0_70 wl_1_70 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6276 wl_0_81 wl_1_81 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6265 wl_0_92 wl_1_92 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5586 wl_0_125 wl_1_125 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5575 wl_0_119 wl_1_119 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5564 wl_0_113 wl_1_113 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4841 wl_0_109 wl_1_109 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4830 wl_0_102 wl_1_102 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6298 wl_0_79 wl_1_79 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5597 wl_0_112 wl_1_112 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4863 wl_0_106 wl_1_106 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4874 wl_0_103 wl_1_103 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4852 wl_0_100 wl_1_100 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4885 wl_0_107 wl_1_107 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4896 wl_0_108 wl_1_108 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8190 wl_0_64 wl_1_64 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_919 wl_0_44 wl_1_44 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_908 wl_0_45 wl_1_45 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4126 wl_0_82 wl_1_82 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4104 wl_0_86 wl_1_86 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4137 wl_0_91 wl_1_91 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4115 wl_0_93 wl_1_93 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3414 wl_0_36 wl_1_36 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3403 wl_0_40 wl_1_40 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3425 wl_0_45 wl_1_45 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4159 wl_0_89 wl_1_89 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4148 wl_0_90 wl_1_90 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2702 wl_0_21 wl_1_21 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2724 wl_0_27 wl_1_27 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2713 wl_0_30 wl_1_30 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3436 wl_0_36 wl_1_36 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3458 wl_0_36 wl_1_36 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3447 wl_0_45 wl_1_45 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2757 wl_0_23 wl_1_23 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2746 wl_0_20 wl_1_20 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2735 wl_0_26 wl_1_26 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3469 wl_0_36 wl_1_36 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2779 wl_0_17 wl_1_17 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2768 wl_0_28 wl_1_28 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6040 wl_0_78 wl_1_78 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6062 wl_0_83 wl_1_83 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6051 wl_0_87 wl_1_87 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5350 wl_0_108 wl_1_108 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5361 wl_0_104 wl_1_104 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6095 wl_0_89 wl_1_89 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6073 wl_0_92 wl_1_92 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6084 wl_0_91 wl_1_91 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5372 wl_0_103 wl_1_103 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5383 wl_0_101 wl_1_101 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5394 wl_0_97 wl_1_97 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4682 wl_0_82 wl_1_82 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4660 wl_0_82 wl_1_82 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4671 wl_0_93 wl_1_93 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3970 wl_0_73 wl_1_73 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3981 wl_0_75 wl_1_75 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4693 wl_0_79 wl_1_79 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3992 wl_0_76 wl_1_76 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2009 wl_0_4 wl_1_4 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1308 wl_0_48 wl_1_48 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1319 wl_0_46 wl_1_46 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_705 wl_0_21 wl_1_21 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_716 wl_0_19 wl_1_19 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_727 wl_0_23 wl_1_23 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_738 wl_0_26 wl_1_26 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3200 wl_0_49 wl_1_49 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_749 wl_0_17 wl_1_17 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3233 wl_0_48 wl_1_48 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3211 wl_0_51 wl_1_51 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3222 wl_0_59 wl_1_59 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2521 wl_0_14 wl_1_14 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2532 wl_0_10 wl_1_10 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2510 wl_0_3 wl_1_3 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3244 wl_0_37 wl_1_37 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3255 wl_0_48 wl_1_48 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3277 wl_0_48 wl_1_48 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3266 wl_0_59 wl_1_59 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1820 wl_0_15 wl_1_15 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2543 wl_0_8 wl_1_8 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2565 wl_0_7 wl_1_7 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2554 wl_0_3 wl_1_3 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3288 wl_0_37 wl_1_37 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3299 wl_0_48 wl_1_48 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2598 wl_0_18 wl_1_18 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2576 wl_0_9 wl_1_9 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1831 wl_0_4 wl_1_4 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2587 wl_0_28 wl_1_28 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1853 wl_0_49 wl_1_49 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1842 wl_0_60 wl_1_60 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1886 wl_0_18 wl_1_18 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1897 wl_0_7 wl_1_7 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1875 wl_0_32 wl_1_32 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1864 wl_0_38 wl_1_38 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5180 wl_0_124 wl_1_124 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5191 wl_0_113 wl_1_113 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4490 wl_0_66 wl_1_66 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6809 wl_0_105 wl_1_105 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_28 wl_0_5 wl_1_5 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_17 wl_0_5 wl_1_5 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_39 wl_0_10 wl_1_10 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1116 wl_0_57 wl_1_57 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1105 wl_0_61 wl_1_61 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1127 wl_0_50 wl_1_50 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1149 wl_0_54 wl_1_54 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1138 wl_0_56 wl_1_56 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_513 wl_0_13 wl_1_13 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_502 wl_0_9 wl_1_9 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_546 wl_0_11 wl_1_11 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_524 wl_0_11 wl_1_11 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_557 wl_0_9 wl_1_9 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_535 wl_0_7 wl_1_7 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_568 wl_0_14 wl_1_14 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_579 wl_0_10 wl_1_10 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3030 wl_0_41 wl_1_41 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3041 wl_0_55 wl_1_55 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2340 wl_0_2 wl_1_2 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3052 wl_0_52 wl_1_52 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3063 wl_0_53 wl_1_53 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3085 wl_0_53 wl_1_53 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3074 wl_0_59 wl_1_59 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2362 wl_0_15 wl_1_15 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2373 wl_0_6 wl_1_6 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2351 wl_0_26 wl_1_26 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3096 wl_0_51 wl_1_51 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2384 wl_0_16 wl_1_16 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2395 wl_0_9 wl_1_9 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1672 wl_0_49 wl_1_49 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1650 wl_0_55 wl_1_55 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1661 wl_0_60 wl_1_60 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1694 wl_0_47 wl_1_47 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1683 wl_0_48 wl_1_48 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8008 wl_0_121 wl_1_121 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8019 wl_0_110 wl_1_110 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7329 wl_0_110 wl_1_110 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7318 wl_0_101 wl_1_101 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7307 wl_0_98 wl_1_98 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6617 wl_0_83 wl_1_83 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6606 wl_0_90 wl_1_90 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6628 wl_0_94 wl_1_94 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5916 wl_0_70 wl_1_70 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5905 wl_0_73 wl_1_73 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5927 wl_0_76 wl_1_76 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6639 wl_0_83 wl_1_83 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5938 wl_0_68 wl_1_68 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5949 wl_0_72 wl_1_72 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7852 wl_0_64 wl_1_64 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7841 wl_0_63 wl_1_63 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7830 wl_0_64 wl_1_64 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7874 wl_0_127 wl_1_127 bl_0_32 bl_1_32 br_0_32
+ br_1_32 sky130_fd_bd_sram__openram_dp_cell_7874/a_38_n79# vdd_uq2046 gnd sky130_fd_bd_sram__openram_dp_cell_7874/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7885 wl_0_116 wl_1_116 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7896 wl_0_105 wl_1_105 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7863 wl_0_63 wl_1_63 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_310 wl_0_26 wl_1_26 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_321 wl_0_27 wl_1_27 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_354 wl_0_17 wl_1_17 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_365 wl_0_27 wl_1_27 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_343 wl_0_28 wl_1_28 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_332 wl_0_30 wl_1_30 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_387 wl_0_20 wl_1_20 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_398 wl_0_11 wl_1_11 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_376 wl_0_30 wl_1_30 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2170 wl_0_24 wl_1_24 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2181 wl_0_30 wl_1_30 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2192 wl_0_19 wl_1_19 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1480 wl_0_33 wl_1_33 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1491 wl_0_45 wl_1_45 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7115 wl_0_120 wl_1_120 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7104 wl_0_100 wl_1_100 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7148 wl_0_111 wl_1_111 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7126 wl_0_109 wl_1_109 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7137 wl_0_98 wl_1_98 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6403 wl_0_77 wl_1_77 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7159 wl_0_112 wl_1_112 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6436 wl_0_68 wl_1_68 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6414 wl_0_68 wl_1_68 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6425 wl_0_72 wl_1_72 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5702 wl_0_95 wl_1_95 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5713 wl_0_127 wl_1_127 bl_0_16 bl_1_16 br_0_16
+ br_1_16 sky130_fd_bd_sram__openram_dp_cell_5713/a_38_n79# vdd_uq3070 gnd sky130_fd_bd_sram__openram_dp_cell_5713/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5724 wl_0_116 wl_1_116 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5735 wl_0_105 wl_1_105 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6447 wl_0_68 wl_1_68 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6458 wl_0_76 wl_1_76 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6469 wl_0_76 wl_1_76 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5768 wl_0_72 wl_1_72 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5757 wl_0_83 wl_1_83 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5746 wl_0_94 wl_1_94 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5779 wl_0_126 wl_1_126 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7660 wl_0_127 wl_1_127 bl_0_48 bl_1_48 br_0_48
+ br_1_48 sky130_fd_bd_sram__openram_dp_cell_7660/a_38_n79# vdd_uq999 gnd sky130_fd_bd_sram__openram_dp_cell_7660/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7671 wl_0_116 wl_1_116 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7682 wl_0_105 wl_1_105 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7693 wl_0_94 wl_1_94 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6992 wl_0_121 wl_1_121 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6970 wl_0_120 wl_1_120 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6981 wl_0_119 wl_1_119 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_140 wl_0_14 wl_1_14 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_173 wl_0_11 wl_1_11 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_162 wl_0_4 wl_1_4 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_151 wl_0_3 wl_1_3 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_184 wl_0_0 wl_1_0 bl_0_49 bl_1_49 br_0_49 br_1_49
+ sky130_fd_bd_sram__openram_dp_cell_184/a_38_n79# vdd_uq958 gnd sky130_fd_bd_sram__openram_dp_cell_184/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_195 wl_0_24 wl_1_24 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5009 wl_0_125 wl_1_125 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4319 wl_0_67 wl_1_67 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4308 wl_0_78 wl_1_78 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3607 wl_0_55 wl_1_55 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2906 wl_0_36 wl_1_36 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3618 wl_0_52 wl_1_52 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3629 wl_0_57 wl_1_57 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2939 wl_0_33 wl_1_33 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2917 wl_0_41 wl_1_41 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2928 wl_0_44 wl_1_44 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6211 wl_0_82 wl_1_82 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6200 wl_0_85 wl_1_85 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5510 wl_0_116 wl_1_116 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6255 wl_0_66 wl_1_66 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6244 wl_0_77 wl_1_77 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6233 wl_0_88 wl_1_88 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6222 wl_0_91 wl_1_91 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5521 wl_0_122 wl_1_122 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5532 wl_0_119 wl_1_119 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5543 wl_0_117 wl_1_117 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6288 wl_0_69 wl_1_69 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6277 wl_0_80 wl_1_80 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6266 wl_0_91 wl_1_91 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5554 wl_0_123 wl_1_123 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5576 wl_0_118 wl_1_118 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5565 wl_0_116 wl_1_116 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4831 wl_0_101 wl_1_101 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4820 wl_0_98 wl_1_98 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6299 wl_0_80 wl_1_80 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5587 wl_0_124 wl_1_124 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5598 wl_0_111 wl_1_111 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4842 wl_0_108 wl_1_108 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4864 wl_0_105 wl_1_105 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4875 wl_0_102 wl_1_102 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4853 wl_0_99 wl_1_99 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4897 wl_0_107 wl_1_107 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4886 wl_0_106 wl_1_106 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8180 wl_0_64 wl_1_64 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8191 wl_0_63 wl_1_63 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7490 wl_0_125 wl_1_125 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_909 wl_0_44 wl_1_44 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4127 wl_0_81 wl_1_81 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4105 wl_0_85 wl_1_85 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4116 wl_0_92 wl_1_92 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3415 wl_0_35 wl_1_35 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3426 wl_0_44 wl_1_44 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3404 wl_0_46 wl_1_46 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4138 wl_0_90 wl_1_90 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4149 wl_0_90 wl_1_90 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2703 wl_0_20 wl_1_20 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2714 wl_0_29 wl_1_29 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3437 wl_0_35 wl_1_35 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3459 wl_0_35 wl_1_35 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3448 wl_0_46 wl_1_46 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2747 wl_0_24 wl_1_24 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2736 wl_0_17 wl_1_17 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2725 wl_0_26 wl_1_26 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2758 wl_0_22 wl_1_22 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2769 wl_0_27 wl_1_27 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6030 wl_0_77 wl_1_77 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6063 wl_0_82 wl_1_82 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6041 wl_0_84 wl_1_84 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6052 wl_0_86 wl_1_86 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5351 wl_0_107 wl_1_107 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5340 wl_0_100 wl_1_100 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6096 wl_0_88 wl_1_88 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6085 wl_0_90 wl_1_90 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6074 wl_0_91 wl_1_91 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5362 wl_0_103 wl_1_103 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5373 wl_0_102 wl_1_102 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5395 wl_0_102 wl_1_102 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5384 wl_0_100 wl_1_100 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4650 wl_0_86 wl_1_86 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4683 wl_0_81 wl_1_81 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4661 wl_0_81 wl_1_81 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4672 wl_0_92 wl_1_92 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3960 wl_0_72 wl_1_72 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3971 wl_0_72 wl_1_72 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4694 wl_0_80 wl_1_80 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3982 wl_0_74 wl_1_74 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3993 wl_0_75 wl_1_75 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1309 wl_0_47 wl_1_47 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_706 wl_0_29 wl_1_29 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_717 wl_0_18 wl_1_18 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_739 wl_0_25 wl_1_25 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_728 wl_0_30 wl_1_30 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3234 wl_0_47 wl_1_47 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3212 wl_0_50 wl_1_50 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3223 wl_0_58 wl_1_58 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3201 wl_0_62 wl_1_62 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2522 wl_0_13 wl_1_13 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2511 wl_0_2 wl_1_2 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2500 wl_0_5 wl_1_5 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3245 wl_0_36 wl_1_36 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3256 wl_0_47 wl_1_47 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3267 wl_0_58 wl_1_58 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1821 wl_0_14 wl_1_14 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2533 wl_0_14 wl_1_14 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2544 wl_0_7 wl_1_7 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2566 wl_0_7 wl_1_7 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2555 wl_0_2 wl_1_2 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1810 wl_0_25 wl_1_25 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3289 wl_0_36 wl_1_36 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3278 wl_0_47 wl_1_47 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2599 wl_0_17 wl_1_17 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2577 wl_0_8 wl_1_8 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1832 wl_0_3 wl_1_3 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2588 wl_0_27 wl_1_27 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1854 wl_0_48 wl_1_48 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1843 wl_0_59 wl_1_59 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1887 wl_0_17 wl_1_17 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1876 wl_0_31 wl_1_31 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1865 wl_0_37 wl_1_37 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1898 wl_0_6 wl_1_6 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5181 wl_0_123 wl_1_123 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5170 wl_0_111 wl_1_111 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5192 wl_0_112 wl_1_112 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4491 wl_0_65 wl_1_65 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4480 wl_0_76 wl_1_76 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3790 wl_0_0 wl_1_0 bl_0_16 bl_1_16 br_0_16 br_1_16
+ sky130_fd_bd_sram__openram_dp_cell_3790/a_38_n79# vdd_uq3070 gnd sky130_fd_bd_sram__openram_dp_cell_3790/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_29 wl_0_4 wl_1_4 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_18 wl_0_4 wl_1_4 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1106 wl_0_60 wl_1_60 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1128 wl_0_49 wl_1_49 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1117 wl_0_56 wl_1_56 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1139 wl_0_55 wl_1_55 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_514 wl_0_12 wl_1_12 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_503 wl_0_8 wl_1_8 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_525 wl_0_14 wl_1_14 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_547 wl_0_10 wl_1_10 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_536 wl_0_6 wl_1_6 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_569 wl_0_13 wl_1_13 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_558 wl_0_8 wl_1_8 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3031 wl_0_40 wl_1_40 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3020 wl_0_43 wl_1_43 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3042 wl_0_54 wl_1_54 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2330 wl_0_12 wl_1_12 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3064 wl_0_50 wl_1_50 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3053 wl_0_52 wl_1_52 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3075 wl_0_58 wl_1_58 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2363 wl_0_14 wl_1_14 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2341 wl_0_1 wl_1_1 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2374 wl_0_5 wl_1_5 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2352 wl_0_25 wl_1_25 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3097 wl_0_50 wl_1_50 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3086 wl_0_52 wl_1_52 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2385 wl_0_16 wl_1_16 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2396 wl_0_8 wl_1_8 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1651 wl_0_54 wl_1_54 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1640 wl_0_57 wl_1_57 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1662 wl_0_59 wl_1_59 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1684 wl_0_47 wl_1_47 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1695 wl_0_48 wl_1_48 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1673 wl_0_52 wl_1_52 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8009 wl_0_120 wl_1_120 bl_0_31 bl_1_31 br_0_31
+ br_1_31 bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7319 wl_0_100 wl_1_100 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7308 wl_0_97 wl_1_97 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6618 wl_0_82 wl_1_82 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6607 wl_0_89 wl_1_89 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6629 wl_0_93 wl_1_93 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5917 wl_0_69 wl_1_69 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5906 wl_0_72 wl_1_72 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5939 wl_0_67 wl_1_67 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5928 wl_0_78 wl_1_78 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7853 wl_0_63 wl_1_63 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7842 wl_0_64 wl_1_64 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7831 wl_0_63 wl_1_63 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7820 wl_0_64 wl_1_64 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7875 wl_0_126 wl_1_126 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7886 wl_0_115 wl_1_115 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7864 wl_0_64 wl_1_64 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7897 wl_0_104 wl_1_104 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_300 wl_0_20 wl_1_20 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_311 wl_0_25 wl_1_25 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_322 wl_0_26 wl_1_26 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_355 wl_0_21 wl_1_21 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_344 wl_0_27 wl_1_27 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_333 wl_0_29 wl_1_29 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_388 wl_0_16 wl_1_16 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_399 wl_0_10 wl_1_10 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_366 wl_0_26 wl_1_26 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_377 wl_0_30 wl_1_30 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2171 wl_0_23 wl_1_23 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2182 wl_0_29 wl_1_29 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2160 wl_0_29 wl_1_29 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2193 wl_0_18 wl_1_18 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1470 wl_0_41 wl_1_41 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1481 wl_0_40 wl_1_40 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1492 wl_0_44 wl_1_44 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7105 wl_0_99 wl_1_99 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7116 wl_0_119 wl_1_119 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7127 wl_0_108 wl_1_108 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7138 wl_0_97 wl_1_97 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6404 wl_0_76 wl_1_76 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7149 wl_0_112 wl_1_112 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6437 wl_0_67 wl_1_67 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6415 wl_0_67 wl_1_67 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6426 wl_0_71 wl_1_71 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5714 wl_0_126 wl_1_126 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5725 wl_0_115 wl_1_115 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6448 wl_0_67 wl_1_67 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6459 wl_0_75 wl_1_75 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5703 wl_0_96 wl_1_96 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5736 wl_0_104 wl_1_104 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5769 wl_0_71 wl_1_71 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5758 wl_0_82 wl_1_82 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5747 wl_0_93 wl_1_93 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7661 wl_0_126 wl_1_126 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7650 wl_0_96 wl_1_96 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7672 wl_0_115 wl_1_115 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7683 wl_0_104 wl_1_104 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7694 wl_0_93 wl_1_93 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6982 wl_0_127 wl_1_127 bl_0_37 bl_1_37 br_0_37
+ br_1_37 sky130_fd_bd_sram__openram_dp_cell_6982/a_38_n79# vdd_uq1726 gnd sky130_fd_bd_sram__openram_dp_cell_6982/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6960 wl_0_123 wl_1_123 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6993 wl_0_120 wl_1_120 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6971 wl_0_119 wl_1_119 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_130 wl_0_11 wl_1_11 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_141 wl_0_13 wl_1_13 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_152 wl_0_2 wl_1_2 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_163 wl_0_3 wl_1_3 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_174 wl_0_10 wl_1_10 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_185 wl_0_8 wl_1_8 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_196 wl_0_23 wl_1_23 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4309 wl_0_77 wl_1_77 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3608 wl_0_62 wl_1_62 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3619 wl_0_51 wl_1_51 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2907 wl_0_35 wl_1_35 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2918 wl_0_40 wl_1_40 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2929 wl_0_43 wl_1_43 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6212 wl_0_81 wl_1_81 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6201 wl_0_84 wl_1_84 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5500 wl_0_126 wl_1_126 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6245 wl_0_76 wl_1_76 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6223 wl_0_80 wl_1_80 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6234 wl_0_87 wl_1_87 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5533 wl_0_127 wl_1_127 bl_0_28 bl_1_28 br_0_28
+ br_1_28 sky130_fd_bd_sram__openram_dp_cell_5533/a_38_n79# vdd_uq2302 gnd sky130_fd_bd_sram__openram_dp_cell_5533/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5522 wl_0_121 wl_1_121 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5511 wl_0_115 wl_1_115 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5544 wl_0_116 wl_1_116 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6256 wl_0_65 wl_1_65 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6278 wl_0_79 wl_1_79 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6267 wl_0_90 wl_1_90 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5555 wl_0_122 wl_1_122 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5577 wl_0_117 wl_1_117 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5566 wl_0_115 wl_1_115 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4821 wl_0_110 wl_1_110 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4832 wl_0_100 wl_1_100 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4810 wl_0_97 wl_1_97 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6289 wl_0_68 wl_1_68 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5588 wl_0_123 wl_1_123 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5599 wl_0_112 wl_1_112 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4843 wl_0_107 wl_1_107 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4854 wl_0_106 wl_1_106 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4865 wl_0_98 wl_1_98 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4887 wl_0_105 wl_1_105 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4898 wl_0_104 wl_1_104 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4876 wl_0_101 wl_1_101 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8181 wl_0_63 wl_1_63 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8170 wl_0_64 wl_1_64 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7480 wl_0_126 wl_1_126 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7491 wl_0_124 wl_1_124 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6790 wl_0_106 wl_1_106 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4106 wl_0_84 wl_1_84 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4117 wl_0_91 wl_1_91 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4128 wl_0_91 wl_1_91 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3416 wl_0_34 wl_1_34 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3405 wl_0_45 wl_1_45 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4139 wl_0_89 wl_1_89 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2704 wl_0_27 wl_1_27 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2715 wl_0_28 wl_1_28 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3438 wl_0_34 wl_1_34 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3427 wl_0_43 wl_1_43 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3449 wl_0_45 wl_1_45 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2748 wl_0_19 wl_1_19 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2726 wl_0_25 wl_1_25 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2737 wl_0_26 wl_1_26 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2759 wl_0_21 wl_1_21 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6020 wl_0_70 wl_1_70 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6031 wl_0_78 wl_1_78 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6042 wl_0_83 wl_1_83 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6053 wl_0_85 wl_1_85 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5330 wl_0_110 wl_1_110 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5352 wl_0_106 wl_1_106 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5341 wl_0_99 wl_1_99 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6064 wl_0_81 wl_1_81 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6086 wl_0_82 wl_1_82 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6097 wl_0_87 wl_1_87 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6075 wl_0_90 wl_1_90 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5374 wl_0_110 wl_1_110 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5363 wl_0_102 wl_1_102 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5385 wl_0_99 wl_1_99 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4640 wl_0_88 wl_1_88 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5396 wl_0_101 wl_1_101 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4651 wl_0_85 wl_1_85 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4662 wl_0_90 wl_1_90 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4673 wl_0_91 wl_1_91 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3961 wl_0_71 wl_1_71 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3972 wl_0_71 wl_1_71 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3950 wl_0_73 wl_1_73 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4695 wl_0_79 wl_1_79 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4684 wl_0_82 wl_1_82 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3994 wl_0_74 wl_1_74 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3983 wl_0_78 wl_1_78 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_718 wl_0_17 wl_1_17 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_707 wl_0_28 wl_1_28 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_729 wl_0_30 wl_1_30 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3213 wl_0_49 wl_1_49 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3224 wl_0_57 wl_1_57 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3202 wl_0_61 wl_1_61 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2512 wl_0_11 wl_1_11 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2523 wl_0_12 wl_1_12 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2501 wl_0_6 wl_1_6 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3246 wl_0_35 wl_1_35 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3235 wl_0_46 wl_1_46 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3257 wl_0_48 wl_1_48 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3268 wl_0_57 wl_1_57 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2534 wl_0_9 wl_1_9 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2545 wl_0_8 wl_1_8 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2556 wl_0_1 wl_1_1 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1811 wl_0_24 wl_1_24 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1800 wl_0_33 wl_1_33 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3279 wl_0_46 wl_1_46 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2567 wl_0_14 wl_1_14 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1822 wl_0_13 wl_1_13 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2578 wl_0_10 wl_1_10 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1833 wl_0_2 wl_1_2 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2589 wl_0_26 wl_1_26 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1844 wl_0_58 wl_1_58 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1888 wl_0_16 wl_1_16 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1877 wl_0_27 wl_1_27 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1866 wl_0_36 wl_1_36 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1855 wl_0_47 wl_1_47 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1899 wl_0_5 wl_1_5 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5160 wl_0_111 wl_1_111 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5182 wl_0_122 wl_1_122 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5171 wl_0_112 wl_1_112 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5193 wl_0_111 wl_1_111 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4492 wl_0_70 wl_1_70 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4470 wl_0_75 wl_1_75 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4481 wl_0_75 wl_1_75 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3780 wl_0_10 wl_1_10 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3791 wl_0_32 wl_1_32 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_19 wl_0_3 wl_1_3 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1107 wl_0_59 wl_1_59 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1129 wl_0_50 wl_1_50 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1118 wl_0_55 wl_1_55 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_504 wl_0_7 wl_1_7 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_526 wl_0_13 wl_1_13 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_515 wl_0_11 wl_1_11 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_537 wl_0_5 wl_1_5 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_548 wl_0_9 wl_1_9 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_559 wl_0_7 wl_1_7 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3010 wl_0_38 wl_1_38 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3032 wl_0_39 wl_1_39 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3021 wl_0_42 wl_1_42 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2320 wl_0_20 wl_1_20 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2331 wl_0_11 wl_1_11 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3065 wl_0_49 wl_1_49 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3043 wl_0_53 wl_1_53 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3054 wl_0_55 wl_1_55 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3076 wl_0_62 wl_1_62 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2353 wl_0_24 wl_1_24 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2364 wl_0_13 wl_1_13 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2342 wl_0_0 wl_1_0 bl_0_23 bl_1_23 br_0_23 br_1_23
+ sky130_fd_bd_sram__openram_dp_cell_2342/a_38_n79# vdd_uq2622 gnd sky130_fd_bd_sram__openram_dp_cell_2342/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3098 wl_0_49 wl_1_49 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3087 wl_0_51 wl_1_51 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2386 wl_0_15 wl_1_15 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2397 wl_0_7 wl_1_7 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2375 wl_0_4 wl_1_4 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1652 wl_0_53 wl_1_53 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1641 wl_0_56 wl_1_56 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1630 wl_0_57 wl_1_57 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1663 wl_0_58 wl_1_58 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1696 wl_0_47 wl_1_47 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1685 wl_0_48 wl_1_48 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1674 wl_0_51 wl_1_51 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7309 wl_0_110 wl_1_110 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6619 wl_0_81 wl_1_81 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6608 wl_0_88 wl_1_88 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5918 wl_0_68 wl_1_68 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5907 wl_0_71 wl_1_71 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5929 wl_0_77 wl_1_77 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7810 wl_0_96 wl_1_96 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7843 wl_0_63 wl_1_63 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7832 wl_0_64 wl_1_64 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7821 wl_0_63 wl_1_63 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7876 wl_0_125 wl_1_125 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7887 wl_0_114 wl_1_114 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7865 wl_0_63 wl_1_63 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7854 wl_0_64 wl_1_64 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7898 wl_0_103 wl_1_103 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_301 wl_0_19 wl_1_19 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_312 wl_0_24 wl_1_24 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_356 wl_0_20 wl_1_20 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_323 wl_0_25 wl_1_25 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_345 wl_0_26 wl_1_26 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_334 wl_0_28 wl_1_28 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_389 wl_0_15 wl_1_15 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_367 wl_0_25 wl_1_25 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_378 wl_0_29 wl_1_29 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2150 wl_0_24 wl_1_24 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2172 wl_0_22 wl_1_22 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2161 wl_0_30 wl_1_30 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2194 wl_0_17 wl_1_17 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2183 wl_0_28 wl_1_28 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1471 wl_0_40 wl_1_40 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1460 wl_0_43 wl_1_43 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1482 wl_0_39 wl_1_39 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1493 wl_0_43 wl_1_43 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_890 wl_0_1 wl_1_1 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7106 wl_0_98 wl_1_98 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7117 wl_0_118 wl_1_118 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7139 wl_0_112 wl_1_112 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7128 wl_0_107 wl_1_107 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6416 wl_0_66 wl_1_66 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6427 wl_0_70 wl_1_70 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6405 wl_0_75 wl_1_75 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5715 wl_0_125 wl_1_125 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5726 wl_0_114 wl_1_114 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6438 wl_0_66 wl_1_66 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6449 wl_0_66 wl_1_66 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5704 wl_0_95 wl_1_95 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5737 wl_0_103 wl_1_103 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5759 wl_0_81 wl_1_81 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5748 wl_0_92 wl_1_92 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7640 wl_0_96 wl_1_96 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7651 wl_0_95 wl_1_95 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7662 wl_0_125 wl_1_125 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7673 wl_0_114 wl_1_114 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6950 wl_0_114 wl_1_114 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7684 wl_0_103 wl_1_103 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7695 wl_0_92 wl_1_92 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6983 wl_0_126 wl_1_126 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6961 wl_0_122 wl_1_122 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6972 wl_0_118 wl_1_118 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6994 wl_0_119 wl_1_119 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_131 wl_0_10 wl_1_10 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_120 wl_0_1 wl_1_1 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_142 wl_0_12 wl_1_12 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_153 wl_0_1 wl_1_1 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_164 wl_0_2 wl_1_2 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_197 wl_0_22 wl_1_22 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_175 wl_0_9 wl_1_9 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_186 wl_0_7 wl_1_7 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1290 wl_0_38 wl_1_38 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3609 wl_0_61 wl_1_61 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2908 wl_0_34 wl_1_34 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2919 wl_0_39 wl_1_39 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6202 wl_0_83 wl_1_83 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5501 wl_0_125 wl_1_125 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6246 wl_0_75 wl_1_75 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6224 wl_0_79 wl_1_79 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6235 wl_0_86 wl_1_86 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6213 wl_0_90 wl_1_90 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5534 wl_0_126 wl_1_126 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5523 wl_0_120 wl_1_120 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5512 wl_0_114 wl_1_114 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6279 wl_0_78 wl_1_78 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6257 wl_0_80 wl_1_80 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6268 wl_0_89 wl_1_89 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5567 wl_0_127 wl_1_127 bl_0_26 bl_1_26 br_0_26
+ br_1_26 sky130_fd_bd_sram__openram_dp_cell_5567/a_38_n79# vdd_uq2430 gnd sky130_fd_bd_sram__openram_dp_cell_5567/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5556 wl_0_121 wl_1_121 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5545 wl_0_115 wl_1_115 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4822 wl_0_110 wl_1_110 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4811 wl_0_103 wl_1_103 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4800 wl_0_99 wl_1_99 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5578 wl_0_116 wl_1_116 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5589 wl_0_112 wl_1_112 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4844 wl_0_106 wl_1_106 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4855 wl_0_104 wl_1_104 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4833 wl_0_99 wl_1_99 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4866 wl_0_97 wl_1_97 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4899 wl_0_103 wl_1_103 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4888 wl_0_104 wl_1_104 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4877 wl_0_100 wl_1_100 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8171 wl_0_63 wl_1_63 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8160 wl_0_64 wl_1_64 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7470 wl_0_125 wl_1_125 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8182 wl_0_64 wl_1_64 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7481 wl_0_125 wl_1_125 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7492 wl_0_123 wl_1_123 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6791 wl_0_105 wl_1_105 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6780 wl_0_99 wl_1_99 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4107 wl_0_83 wl_1_83 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4118 wl_0_90 wl_1_90 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3417 wl_0_33 wl_1_33 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3406 wl_0_44 wl_1_44 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4129 wl_0_90 wl_1_90 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2705 wl_0_26 wl_1_26 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3439 wl_0_33 wl_1_33 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3428 wl_0_42 wl_1_42 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2727 wl_0_24 wl_1_24 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2738 wl_0_25 wl_1_25 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2716 wl_0_27 wl_1_27 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2749 wl_0_18 wl_1_18 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6010 wl_0_65 wl_1_65 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6021 wl_0_66 wl_1_66 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6032 wl_0_77 wl_1_77 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6043 wl_0_82 wl_1_82 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6054 wl_0_84 wl_1_84 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5331 wl_0_109 wl_1_109 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5320 wl_0_101 wl_1_101 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5342 wl_0_98 wl_1_98 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6087 wl_0_81 wl_1_81 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6065 wl_0_88 wl_1_88 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6076 wl_0_89 wl_1_89 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5353 wl_0_110 wl_1_110 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5375 wl_0_109 wl_1_109 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5364 wl_0_101 wl_1_101 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5386 wl_0_98 wl_1_98 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4630 wl_0_88 wl_1_88 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4641 wl_0_87 wl_1_87 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6098 wl_0_94 wl_1_94 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5397 wl_0_100 wl_1_100 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4652 wl_0_84 wl_1_84 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4663 wl_0_89 wl_1_89 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4674 wl_0_90 wl_1_90 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3962 wl_0_70 wl_1_70 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3951 wl_0_72 wl_1_72 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3940 wl_0_78 wl_1_78 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4696 wl_0_80 wl_1_80 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4685 wl_0_81 wl_1_81 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3973 wl_0_70 wl_1_70 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3995 wl_0_73 wl_1_73 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3984 wl_0_77 wl_1_77 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_719 wl_0_20 wl_1_20 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_708 wl_0_27 wl_1_27 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3225 wl_0_56 wl_1_56 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3203 wl_0_59 wl_1_59 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3214 wl_0_60 wl_1_60 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2513 wl_0_10 wl_1_10 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2502 wl_0_5 wl_1_5 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3247 wl_0_34 wl_1_34 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3236 wl_0_45 wl_1_45 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3258 wl_0_47 wl_1_47 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2535 wl_0_14 wl_1_14 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2524 wl_0_11 wl_1_11 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2546 wl_0_8 wl_1_8 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2557 wl_0_0 wl_1_0 bl_0_4 bl_1_4 br_0_4 br_1_4
+ sky130_fd_bd_sram__openram_dp_cell_2557/a_38_n79# vdd_uq3838 gnd sky130_fd_bd_sram__openram_dp_cell_2557/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1812 wl_0_23 wl_1_23 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1801 wl_0_32 wl_1_32 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3269 wl_0_56 wl_1_56 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2568 wl_0_13 wl_1_13 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1823 wl_0_12 wl_1_12 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2579 wl_0_9 wl_1_9 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1834 wl_0_1 wl_1_1 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1845 wl_0_57 wl_1_57 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1878 wl_0_26 wl_1_26 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1867 wl_0_35 wl_1_35 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1856 wl_0_46 wl_1_46 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1889 wl_0_15 wl_1_15 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5150 wl_0_120 wl_1_120 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5183 wl_0_121 wl_1_121 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5172 wl_0_111 wl_1_111 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5161 wl_0_112 wl_1_112 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5194 wl_0_110 wl_1_110 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4460 wl_0_66 wl_1_66 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4482 wl_0_74 wl_1_74 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4471 wl_0_76 wl_1_76 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3770 wl_0_20 wl_1_20 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3781 wl_0_9 wl_1_9 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4493 wl_0_69 wl_1_69 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3792 wl_0_31 wl_1_31 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1119 wl_0_54 wl_1_54 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1108 wl_0_58 wl_1_58 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_505 wl_0_6 wl_1_6 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_527 wl_0_12 wl_1_12 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_516 wl_0_10 wl_1_10 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_538 wl_0_4 wl_1_4 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3000 wl_0_34 wl_1_34 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_549 wl_0_8 wl_1_8 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3011 wl_0_37 wl_1_37 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3033 wl_0_38 wl_1_38 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3022 wl_0_41 wl_1_41 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2321 wl_0_19 wl_1_19 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2310 wl_0_15 wl_1_15 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3066 wl_0_51 wl_1_51 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3044 wl_0_52 wl_1_52 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3055 wl_0_54 wl_1_54 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2354 wl_0_23 wl_1_23 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2343 wl_0_16 wl_1_16 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2365 wl_0_12 wl_1_12 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2332 wl_0_10 wl_1_10 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1620 wl_0_49 wl_1_49 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3088 wl_0_50 wl_1_50 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3077 wl_0_61 wl_1_61 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3099 wl_0_62 wl_1_62 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2387 wl_0_12 wl_1_12 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2398 wl_0_6 wl_1_6 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2376 wl_0_3 wl_1_3 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1653 wl_0_52 wl_1_52 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1642 wl_0_55 wl_1_55 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1631 wl_0_56 wl_1_56 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1686 wl_0_47 wl_1_47 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1664 wl_0_57 wl_1_57 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1675 wl_0_62 wl_1_62 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1697 wl_0_48 wl_1_48 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4290 wl_0_80 wl_1_80 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6609 wl_0_87 wl_1_87 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5908 wl_0_78 wl_1_78 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5919 wl_0_67 wl_1_67 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7800 wl_0_96 wl_1_96 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7811 wl_0_95 wl_1_95 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7844 wl_0_64 wl_1_64 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7833 wl_0_63 wl_1_63 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7822 wl_0_64 wl_1_64 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7877 wl_0_124 wl_1_124 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7866 wl_0_64 wl_1_64 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7855 wl_0_63 wl_1_63 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7888 wl_0_113 wl_1_113 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7899 wl_0_102 wl_1_102 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_302 wl_0_18 wl_1_18 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_313 wl_0_23 wl_1_23 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_324 wl_0_24 wl_1_24 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_346 wl_0_25 wl_1_25 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_335 wl_0_27 wl_1_27 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_357 wl_0_19 wl_1_19 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_368 wl_0_24 wl_1_24 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_379 wl_0_28 wl_1_28 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2140 wl_0_21 wl_1_21 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2151 wl_0_23 wl_1_23 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2173 wl_0_21 wl_1_21 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2162 wl_0_30 wl_1_30 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2184 wl_0_27 wl_1_27 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2195 wl_0_27 wl_1_27 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1461 wl_0_42 wl_1_42 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1450 wl_0_45 wl_1_45 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1483 wl_0_38 wl_1_38 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1472 wl_0_39 wl_1_39 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1494 wl_0_42 wl_1_42 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_880 wl_0_11 wl_1_11 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_891 wl_0_0 wl_1_0 bl_0_40 bl_1_40 br_0_40 br_1_40
+ sky130_fd_bd_sram__openram_dp_cell_891/a_38_n79# vdd_uq1534 gnd sky130_fd_bd_sram__openram_dp_cell_891/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7118 wl_0_117 wl_1_117 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7129 wl_0_106 wl_1_106 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7107 wl_0_97 wl_1_97 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6428 wl_0_65 wl_1_65 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6417 wl_0_68 wl_1_68 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6406 wl_0_74 wl_1_74 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5716 wl_0_124 wl_1_124 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6439 wl_0_67 wl_1_67 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5705 wl_0_96 wl_1_96 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5727 wl_0_113 wl_1_113 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5738 wl_0_102 wl_1_102 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5749 wl_0_91 wl_1_91 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7630 wl_0_96 wl_1_96 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7641 wl_0_95 wl_1_95 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7652 wl_0_96 wl_1_96 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7663 wl_0_124 wl_1_124 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6940 wl_0_120 wl_1_120 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7674 wl_0_113 wl_1_113 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7685 wl_0_102 wl_1_102 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6984 wl_0_125 wl_1_125 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6962 wl_0_121 wl_1_121 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6973 wl_0_117 wl_1_117 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6951 wl_0_113 wl_1_113 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7696 wl_0_91 wl_1_91 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6995 wl_0_118 wl_1_118 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_110 wl_0_8 wl_1_8 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_121 wl_0_0 wl_1_0 bl_0_52 bl_1_52 br_0_52 br_1_52
+ sky130_fd_bd_sram__openram_dp_cell_121/a_38_n79# vdd_uq766 gnd sky130_fd_bd_sram__openram_dp_cell_121/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_143 wl_0_11 wl_1_11 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_132 wl_0_9 wl_1_9 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_154 wl_0_0 wl_1_0 bl_0_54 bl_1_54 br_0_54 br_1_54
+ sky130_fd_bd_sram__openram_dp_cell_154/a_38_n79# vdd_uq638 gnd sky130_fd_bd_sram__openram_dp_cell_154/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_198 wl_0_21 wl_1_21 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_176 wl_0_8 wl_1_8 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_187 wl_0_6 wl_1_6 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_165 wl_0_1 wl_1_1 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1280 wl_0_48 wl_1_48 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1291 wl_0_37 wl_1_37 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2909 wl_0_33 wl_1_33 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6203 wl_0_82 wl_1_82 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6225 wl_0_80 wl_1_80 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6236 wl_0_85 wl_1_85 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6214 wl_0_89 wl_1_89 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5502 wl_0_124 wl_1_124 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5524 wl_0_119 wl_1_119 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5513 wl_0_113 wl_1_113 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6247 wl_0_74 wl_1_74 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6258 wl_0_79 wl_1_79 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6269 wl_0_88 wl_1_88 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5568 wl_0_126 wl_1_126 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5535 wl_0_125 wl_1_125 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5557 wl_0_120 wl_1_120 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5546 wl_0_114 wl_1_114 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4823 wl_0_109 wl_1_109 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4812 wl_0_102 wl_1_102 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4801 wl_0_98 wl_1_98 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5579 wl_0_115 wl_1_115 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4834 wl_0_109 wl_1_109 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4845 wl_0_105 wl_1_105 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4856 wl_0_98 wl_1_98 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4867 wl_0_110 wl_1_110 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4889 wl_0_103 wl_1_103 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4878 wl_0_99 wl_1_99 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8172 wl_0_64 wl_1_64 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8161 wl_0_63 wl_1_63 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8150 wl_0_64 wl_1_64 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7460 wl_0_116 wl_1_116 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8183 wl_0_63 wl_1_63 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7482 wl_0_124 wl_1_124 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7493 wl_0_122 wl_1_122 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7471 wl_0_122 wl_1_122 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6770 wl_0_109 wl_1_109 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6792 wl_0_104 wl_1_104 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6781 wl_0_98 wl_1_98 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4108 wl_0_82 wl_1_82 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4119 wl_0_89 wl_1_89 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3407 wl_0_43 wl_1_43 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2706 wl_0_25 wl_1_25 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3418 wl_0_39 wl_1_39 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3429 wl_0_41 wl_1_41 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2728 wl_0_23 wl_1_23 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2739 wl_0_24 wl_1_24 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2717 wl_0_23 wl_1_23 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6011 wl_0_67 wl_1_67 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6000 wl_0_70 wl_1_70 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6022 wl_0_65 wl_1_65 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6033 wl_0_76 wl_1_76 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6044 wl_0_81 wl_1_81 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5332 wl_0_108 wl_1_108 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5310 wl_0_101 wl_1_101 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5321 wl_0_100 wl_1_100 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5343 wl_0_97 wl_1_97 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6055 wl_0_83 wl_1_83 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6088 wl_0_86 wl_1_86 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6077 wl_0_88 wl_1_88 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6066 wl_0_87 wl_1_87 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5365 wl_0_110 wl_1_110 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5354 wl_0_109 wl_1_109 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5376 wl_0_108 wl_1_108 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4631 wl_0_87 wl_1_87 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6099 wl_0_93 wl_1_93 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4620 wl_0_94 wl_1_94 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5398 wl_0_99 wl_1_99 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5387 wl_0_97 wl_1_97 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3930 wl_0_66 wl_1_66 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4653 wl_0_83 wl_1_83 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4664 wl_0_88 wl_1_88 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4642 wl_0_94 wl_1_94 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3963 wl_0_69 wl_1_69 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3952 wl_0_71 wl_1_71 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3941 wl_0_77 wl_1_77 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4697 wl_0_79 wl_1_79 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4675 wl_0_89 wl_1_89 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4686 wl_0_94 wl_1_94 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3974 wl_0_69 wl_1_69 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3996 wl_0_72 wl_1_72 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3985 wl_0_76 wl_1_76 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7290 wl_0_108 wl_1_108 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_709 wl_0_26 wl_1_26 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3204 wl_0_58 wl_1_58 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3215 wl_0_59 wl_1_59 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2514 wl_0_9 wl_1_9 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2503 wl_0_4 wl_1_4 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3248 wl_0_33 wl_1_33 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3237 wl_0_44 wl_1_44 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3259 wl_0_48 wl_1_48 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3226 wl_0_55 wl_1_55 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2536 wl_0_11 wl_1_11 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2525 wl_0_10 wl_1_10 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2547 wl_0_7 wl_1_7 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1802 wl_0_31 wl_1_31 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1813 wl_0_22 wl_1_22 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1824 wl_0_11 wl_1_11 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2569 wl_0_12 wl_1_12 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2558 wl_0_8 wl_1_8 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1835 wl_0_0 wl_1_0 bl_0_48 bl_1_48 br_0_48 br_1_48
+ sky130_fd_bd_sram__openram_dp_cell_1835/a_38_n79# vdd_uq999 gnd sky130_fd_bd_sram__openram_dp_cell_1835/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1879 wl_0_25 wl_1_25 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1868 wl_0_34 wl_1_34 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1857 wl_0_45 wl_1_45 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1846 wl_0_56 wl_1_56 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5151 wl_0_119 wl_1_119 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5140 wl_0_113 wl_1_113 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5184 wl_0_120 wl_1_120 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5173 wl_0_112 wl_1_112 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5162 wl_0_111 wl_1_111 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5195 wl_0_109 wl_1_109 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4461 wl_0_65 wl_1_65 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4483 wl_0_73 wl_1_73 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4450 wl_0_76 wl_1_76 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4472 wl_0_78 wl_1_78 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3771 wl_0_19 wl_1_19 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3760 wl_0_30 wl_1_30 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4494 wl_0_74 wl_1_74 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3782 wl_0_8 wl_1_8 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3793 wl_0_62 wl_1_62 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1109 wl_0_57 wl_1_57 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_528 wl_0_14 wl_1_14 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_517 wl_0_1 wl_1_1 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_506 wl_0_5 wl_1_5 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_539 wl_0_3 wl_1_3 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3001 wl_0_33 wl_1_33 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3012 wl_0_36 wl_1_36 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3023 wl_0_40 wl_1_40 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2300 wl_0_19 wl_1_19 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2322 wl_0_18 wl_1_18 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2311 wl_0_29 wl_1_29 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3067 wl_0_50 wl_1_50 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3045 wl_0_51 wl_1_51 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3056 wl_0_53 wl_1_53 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3034 wl_0_62 wl_1_62 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2355 wl_0_22 wl_1_22 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2344 wl_0_15 wl_1_15 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2333 wl_0_9 wl_1_9 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3089 wl_0_49 wl_1_49 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3078 wl_0_60 wl_1_60 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1610 wl_0_59 wl_1_59 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2366 wl_0_16 wl_1_16 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2388 wl_0_11 wl_1_11 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2377 wl_0_2 wl_1_2 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2399 wl_0_5 wl_1_5 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1654 wl_0_51 wl_1_51 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1632 wl_0_55 wl_1_55 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1621 wl_0_62 wl_1_62 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1643 wl_0_62 wl_1_62 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1687 wl_0_48 wl_1_48 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1665 wl_0_56 wl_1_56 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1676 wl_0_61 wl_1_61 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1698 wl_0_47 wl_1_47 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4291 wl_0_79 wl_1_79 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4280 wl_0_80 wl_1_80 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3590 wl_0_58 wl_1_58 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5909 wl_0_77 wl_1_77 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7801 wl_0_95 wl_1_95 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7834 wl_0_64 wl_1_64 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7823 wl_0_63 wl_1_63 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7812 wl_0_64 wl_1_64 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7878 wl_0_123 wl_1_123 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7867 wl_0_63 wl_1_63 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7856 wl_0_64 wl_1_64 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7845 wl_0_63 wl_1_63 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7889 wl_0_112 wl_1_112 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_303 wl_0_17 wl_1_17 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_314 wl_0_22 wl_1_22 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_325 wl_0_23 wl_1_23 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_347 wl_0_24 wl_1_24 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_336 wl_0_26 wl_1_26 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_358 wl_0_18 wl_1_18 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_369 wl_0_23 wl_1_23 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2130 wl_0_0 wl_1_0 bl_0_19 bl_1_19 br_0_19 br_1_19
+ sky130_fd_bd_sram__openram_dp_cell_2130/a_38_n79# vdd_uq2878 gnd sky130_fd_bd_sram__openram_dp_cell_2130/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2152 wl_0_22 wl_1_22 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2141 wl_0_20 wl_1_20 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2163 wl_0_29 wl_1_29 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2174 wl_0_20 wl_1_20 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2185 wl_0_26 wl_1_26 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2196 wl_0_26 wl_1_26 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1440 wl_0_40 wl_1_40 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1462 wl_0_41 wl_1_41 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1451 wl_0_44 wl_1_44 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1484 wl_0_37 wl_1_37 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1473 wl_0_38 wl_1_38 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1495 wl_0_41 wl_1_41 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_892 wl_0_16 wl_1_16 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_881 wl_0_10 wl_1_10 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_870 wl_0_7 wl_1_7 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7108 wl_0_127 wl_1_127 bl_0_39 bl_1_39 br_0_39
+ br_1_39 sky130_fd_bd_sram__openram_dp_cell_7108/a_38_n79# vdd_uq1598 gnd sky130_fd_bd_sram__openram_dp_cell_7108/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7119 wl_0_116 wl_1_116 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6418 wl_0_66 wl_1_66 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6407 wl_0_73 wl_1_73 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5717 wl_0_123 wl_1_123 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6429 wl_0_74 wl_1_74 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5706 wl_0_95 wl_1_95 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5728 wl_0_112 wl_1_112 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5739 wl_0_101 wl_1_101 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7620 wl_0_112 wl_1_112 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7631 wl_0_95 wl_1_95 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7642 wl_0_96 wl_1_96 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7664 wl_0_123 wl_1_123 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6941 wl_0_119 wl_1_119 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6930 wl_0_116 wl_1_116 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7675 wl_0_112 wl_1_112 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7686 wl_0_101 wl_1_101 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7653 wl_0_95 wl_1_95 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6963 wl_0_127 wl_1_127 bl_0_38 bl_1_38 br_0_38
+ br_1_38 sky130_fd_bd_sram__openram_dp_cell_6963/a_38_n79# vdd_uq1662 gnd sky130_fd_bd_sram__openram_dp_cell_6963/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6952 wl_0_125 wl_1_125 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6974 wl_0_116 wl_1_116 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7697 wl_0_90 wl_1_90 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6985 wl_0_124 wl_1_124 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6996 wl_0_117 wl_1_117 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_111 wl_0_14 wl_1_14 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_100 wl_0_7 wl_1_7 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_122 wl_0_7 wl_1_7 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_155 wl_0_11 wl_1_11 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_144 wl_0_10 wl_1_10 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_133 wl_0_8 wl_1_8 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_177 wl_0_7 wl_1_7 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_166 wl_0_0 wl_1_0 bl_0_51 bl_1_51 br_0_51 br_1_51
+ sky130_fd_bd_sram__openram_dp_cell_166/a_38_n79# vdd_uq830 gnd sky130_fd_bd_sram__openram_dp_cell_166/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_188 wl_0_5 wl_1_5 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_199 wl_0_20 wl_1_20 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1270 wl_0_58 wl_1_58 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1292 wl_0_36 wl_1_36 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1281 wl_0_47 wl_1_47 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6226 wl_0_79 wl_1_79 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6204 wl_0_81 wl_1_81 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6237 wl_0_84 wl_1_84 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6215 wl_0_88 wl_1_88 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5503 wl_0_123 wl_1_123 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5514 wl_0_122 wl_1_122 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5525 wl_0_118 wl_1_118 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6248 wl_0_73 wl_1_73 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6259 wl_0_80 wl_1_80 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5536 wl_0_124 wl_1_124 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5558 wl_0_119 wl_1_119 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5547 wl_0_113 wl_1_113 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4813 wl_0_101 wl_1_101 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4802 wl_0_97 wl_1_97 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5569 wl_0_125 wl_1_125 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4824 wl_0_108 wl_1_108 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4835 wl_0_108 wl_1_108 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4846 wl_0_104 wl_1_104 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4857 wl_0_97 wl_1_97 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4868 wl_0_109 wl_1_109 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4879 wl_0_98 wl_1_98 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8162 wl_0_64 wl_1_64 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8151 wl_0_63 wl_1_63 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8140 wl_0_64 wl_1_64 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7450 wl_0_117 wl_1_117 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7461 wl_0_115 wl_1_115 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8184 wl_0_64 wl_1_64 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8173 wl_0_63 wl_1_63 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7483 wl_0_123 wl_1_123 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7494 wl_0_121 wl_1_121 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7472 wl_0_121 wl_1_121 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6771 wl_0_108 wl_1_108 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6760 wl_0_106 wl_1_106 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6782 wl_0_97 wl_1_97 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6793 wl_0_103 wl_1_103 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4109 wl_0_81 wl_1_81 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3408 wl_0_42 wl_1_42 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3419 wl_0_38 wl_1_38 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2707 wl_0_24 wl_1_24 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2729 wl_0_22 wl_1_22 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2718 wl_0_22 wl_1_22 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6001 wl_0_69 wl_1_69 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5300 wl_0_107 wl_1_107 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6034 wl_0_75 wl_1_75 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6012 wl_0_78 wl_1_78 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6023 wl_0_78 wl_1_78 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6045 wl_0_93 wl_1_93 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5333 wl_0_107 wl_1_107 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5311 wl_0_100 wl_1_100 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5322 wl_0_99 wl_1_99 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6056 wl_0_82 wl_1_82 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6067 wl_0_86 wl_1_86 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6078 wl_0_87 wl_1_87 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5366 wl_0_109 wl_1_109 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5355 wl_0_108 wl_1_108 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5344 wl_0_104 wl_1_104 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6089 wl_0_85 wl_1_85 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4632 wl_0_86 wl_1_86 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4610 wl_0_90 wl_1_90 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4621 wl_0_93 wl_1_93 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5377 wl_0_107 wl_1_107 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5388 wl_0_106 wl_1_106 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5399 wl_0_98 wl_1_98 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3920 wl_0_76 wl_1_76 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4654 wl_0_82 wl_1_82 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4665 wl_0_87 wl_1_87 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4643 wl_0_93 wl_1_93 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3931 wl_0_65 wl_1_65 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3953 wl_0_70 wl_1_70 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3942 wl_0_76 wl_1_76 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4698 wl_0_80 wl_1_80 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4676 wl_0_88 wl_1_88 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4687 wl_0_93 wl_1_93 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3964 wl_0_68 wl_1_68 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3975 wl_0_68 wl_1_68 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3997 wl_0_71 wl_1_71 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3986 wl_0_75 wl_1_75 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7280 wl_0_108 wl_1_108 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7291 wl_0_107 wl_1_107 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6590 wl_0_88 wl_1_88 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3216 wl_0_48 wl_1_48 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3205 wl_0_57 wl_1_57 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2504 wl_0_6 wl_1_6 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3238 wl_0_43 wl_1_43 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3249 wl_0_48 wl_1_48 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3227 wl_0_54 wl_1_54 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2526 wl_0_14 wl_1_14 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2515 wl_0_13 wl_1_13 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2537 wl_0_10 wl_1_10 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2548 wl_0_5 wl_1_5 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1803 wl_0_30 wl_1_30 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1814 wl_0_21 wl_1_21 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1825 wl_0_10 wl_1_10 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2559 wl_0_7 wl_1_7 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1836 wl_0_32 wl_1_32 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1869 wl_0_33 wl_1_33 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1858 wl_0_44 wl_1_44 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1847 wl_0_55 wl_1_55 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5130 wl_0_123 wl_1_123 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5141 wl_0_116 wl_1_116 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5185 wl_0_119 wl_1_119 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5152 wl_0_118 wl_1_118 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5174 wl_0_111 wl_1_111 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5163 wl_0_112 wl_1_112 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4440 wl_0_72 wl_1_72 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5196 wl_0_108 wl_1_108 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4462 wl_0_74 wl_1_74 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4451 wl_0_75 wl_1_75 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4473 wl_0_77 wl_1_77 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3772 wl_0_18 wl_1_18 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3761 wl_0_29 wl_1_29 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3750 wl_0_40 wl_1_40 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4484 wl_0_72 wl_1_72 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4495 wl_0_73 wl_1_73 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3783 wl_0_7 wl_1_7 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3794 wl_0_61 wl_1_61 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_507 wl_0_14 wl_1_14 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_529 wl_0_13 wl_1_13 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_518 wl_0_0 wl_1_0 bl_0_42 bl_1_42 br_0_42 br_1_42
+ sky130_fd_bd_sram__openram_dp_cell_518/a_38_n79# vdd_uq1406 gnd sky130_fd_bd_sram__openram_dp_cell_518/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3013 wl_0_35 wl_1_35 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3024 wl_0_39 wl_1_39 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3002 wl_0_46 wl_1_46 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2301 wl_0_16 wl_1_16 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2312 wl_0_28 wl_1_28 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3046 wl_0_50 wl_1_50 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3057 wl_0_52 wl_1_52 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3035 wl_0_61 wl_1_61 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2356 wl_0_21 wl_1_21 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2323 wl_0_16 wl_1_16 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2345 wl_0_16 wl_1_16 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2334 wl_0_8 wl_1_8 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3068 wl_0_49 wl_1_49 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1600 wl_0_49 wl_1_49 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1611 wl_0_58 wl_1_58 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3079 wl_0_59 wl_1_59 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2367 wl_0_15 wl_1_15 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2389 wl_0_10 wl_1_10 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2378 wl_0_1 wl_1_1 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1633 wl_0_54 wl_1_54 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1622 wl_0_61 wl_1_61 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1644 wl_0_61 wl_1_61 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1655 wl_0_50 wl_1_50 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1666 wl_0_55 wl_1_55 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1677 wl_0_60 wl_1_60 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1688 wl_0_47 wl_1_47 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1699 wl_0_48 wl_1_48 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4270 wl_0_68 wl_1_68 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4281 wl_0_79 wl_1_79 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3580 wl_0_56 wl_1_56 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4292 wl_0_94 wl_1_94 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3591 wl_0_57 wl_1_57 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2890 wl_0_44 wl_1_44 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7802 wl_0_96 wl_1_96 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7835 wl_0_63 wl_1_63 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7824 wl_0_64 wl_1_64 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7813 wl_0_63 wl_1_63 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7868 wl_0_64 wl_1_64 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7857 wl_0_63 wl_1_63 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7846 wl_0_64 wl_1_64 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7879 wl_0_122 wl_1_122 bl_0_32 bl_1_32 br_0_32
+ br_1_32 bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_304 wl_0_22 wl_1_22 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_326 wl_0_22 wl_1_22 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_315 wl_0_21 wl_1_21 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_337 wl_0_25 wl_1_25 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_359 wl_0_17 wl_1_17 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_348 wl_0_23 wl_1_23 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2131 wl_0_14 wl_1_14 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2120 wl_0_7 wl_1_7 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2153 wl_0_21 wl_1_21 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2142 wl_0_19 wl_1_19 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2164 wl_0_30 wl_1_30 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2175 wl_0_19 wl_1_19 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2186 wl_0_25 wl_1_25 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2197 wl_0_25 wl_1_25 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1452 wl_0_37 wl_1_37 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1441 wl_0_39 wl_1_39 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1430 wl_0_46 wl_1_46 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1485 wl_0_33 wl_1_33 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1474 wl_0_37 wl_1_37 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1463 wl_0_39 wl_1_39 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1496 wl_0_45 wl_1_45 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_860 wl_0_14 wl_1_14 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_893 wl_0_15 wl_1_15 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_882 wl_0_9 wl_1_9 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_871 wl_0_6 wl_1_6 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7109 wl_0_126 wl_1_126 bl_0_39 bl_1_39 br_0_39
+ br_1_39 bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6408 wl_0_70 wl_1_70 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6419 wl_0_78 wl_1_78 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5707 wl_0_96 wl_1_96 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5718 wl_0_122 wl_1_122 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5729 wl_0_111 wl_1_111 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7610 wl_0_104 wl_1_104 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7621 wl_0_111 wl_1_111 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7632 wl_0_96 wl_1_96 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7643 wl_0_95 wl_1_95 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7665 wl_0_122 wl_1_122 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6920 wl_0_118 wl_1_118 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6931 wl_0_115 wl_1_115 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7676 wl_0_111 wl_1_111 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7654 wl_0_96 wl_1_96 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6953 wl_0_127 wl_1_127 bl_0_33 bl_1_33 br_0_33
+ br_1_33 sky130_fd_bd_sram__openram_dp_cell_6953/a_38_n79# vdd_uq1982 gnd sky130_fd_bd_sram__openram_dp_cell_6953/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6964 wl_0_126 wl_1_126 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6942 wl_0_118 wl_1_118 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6975 wl_0_115 wl_1_115 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7687 wl_0_100 wl_1_100 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7698 wl_0_89 wl_1_89 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6986 wl_0_123 wl_1_123 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6997 wl_0_116 wl_1_116 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_112 wl_0_13 wl_1_13 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_101 wl_0_8 wl_1_8 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_145 wl_0_9 wl_1_9 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_134 wl_0_7 wl_1_7 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_123 wl_0_6 wl_1_6 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_156 wl_0_10 wl_1_10 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_178 wl_0_6 wl_1_6 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_189 wl_0_4 wl_1_4 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_167 wl_0_3 wl_1_3 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1260 wl_0_34 wl_1_34 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1271 wl_0_57 wl_1_57 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1293 wl_0_35 wl_1_35 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1282 wl_0_46 wl_1_46 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_690 wl_0_30 wl_1_30 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6216 wl_0_87 wl_1_87 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6205 wl_0_88 wl_1_88 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6227 wl_0_94 wl_1_94 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5504 wl_0_122 wl_1_122 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5515 wl_0_121 wl_1_121 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6249 wl_0_72 wl_1_72 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6238 wl_0_83 wl_1_83 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5537 wl_0_123 wl_1_123 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5559 wl_0_118 wl_1_118 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5548 wl_0_118 wl_1_118 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5526 wl_0_117 wl_1_117 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4803 wl_0_100 wl_1_100 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4814 wl_0_100 wl_1_100 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4825 wl_0_107 wl_1_107 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4836 wl_0_107 wl_1_107 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4847 wl_0_103 wl_1_103 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4869 wl_0_108 wl_1_108 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4858 wl_0_103 wl_1_103 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8163 wl_0_63 wl_1_63 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8152 wl_0_64 wl_1_64 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8141 wl_0_63 wl_1_63 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8130 wl_0_64 wl_1_64 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7451 wl_0_116 wl_1_116 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7440 wl_0_114 wl_1_114 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8185 wl_0_63 wl_1_63 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8174 wl_0_64 wl_1_64 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7473 wl_0_127 wl_1_127 bl_0_57 bl_1_57 br_0_57
+ br_1_57 sky130_fd_bd_sram__openram_dp_cell_7473/a_38_n79# vdd_uq446 gnd sky130_fd_bd_sram__openram_dp_cell_7473/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7484 wl_0_122 wl_1_122 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7462 wl_0_113 wl_1_113 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6750 wl_0_97 wl_1_97 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7495 wl_0_122 wl_1_122 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6783 wl_0_109 wl_1_109 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6772 wl_0_107 wl_1_107 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6761 wl_0_105 wl_1_105 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6794 wl_0_102 wl_1_102 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1090 wl_0_51 wl_1_51 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3409 wl_0_41 wl_1_41 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2719 wl_0_21 wl_1_21 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2708 wl_0_30 wl_1_30 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6002 wl_0_68 wl_1_68 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6035 wl_0_76 wl_1_76 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6013 wl_0_77 wl_1_77 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6024 wl_0_77 wl_1_77 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5301 wl_0_110 wl_1_110 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5334 wl_0_106 wl_1_106 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5312 wl_0_99 wl_1_99 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5323 wl_0_98 wl_1_98 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6057 wl_0_81 wl_1_81 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6068 wl_0_85 wl_1_85 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6079 wl_0_86 wl_1_86 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6046 wl_0_92 wl_1_92 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5367 wl_0_108 wl_1_108 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5356 wl_0_107 wl_1_107 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5345 wl_0_103 wl_1_103 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4600 wl_0_84 wl_1_84 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4611 wl_0_89 wl_1_89 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4622 wl_0_92 wl_1_92 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5378 wl_0_106 wl_1_106 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5389 wl_0_105 wl_1_105 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3910 wl_0_67 wl_1_67 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3921 wl_0_75 wl_1_75 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4655 wl_0_81 wl_1_81 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4633 wl_0_85 wl_1_85 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4644 wl_0_92 wl_1_92 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3932 wl_0_68 wl_1_68 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3954 wl_0_69 wl_1_69 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3943 wl_0_75 wl_1_75 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4699 wl_0_79 wl_1_79 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4666 wl_0_86 wl_1_86 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4677 wl_0_87 wl_1_87 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4688 wl_0_92 wl_1_92 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3965 wl_0_67 wl_1_67 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3976 wl_0_67 wl_1_67 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3987 wl_0_74 wl_1_74 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3998 wl_0_70 wl_1_70 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7281 wl_0_107 wl_1_107 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7270 wl_0_100 wl_1_100 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7292 wl_0_98 wl_1_98 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6591 wl_0_87 wl_1_87 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6580 wl_0_92 wl_1_92 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5890 wl_0_66 wl_1_66 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3206 wl_0_56 wl_1_56 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2505 wl_0_6 wl_1_6 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3239 wl_0_42 wl_1_42 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3217 wl_0_47 wl_1_47 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3228 wl_0_53 wl_1_53 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2516 wl_0_12 wl_1_12 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2538 wl_0_9 wl_1_9 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2527 wl_0_9 wl_1_9 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1815 wl_0_20 wl_1_20 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1826 wl_0_9 wl_1_9 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2549 wl_0_4 wl_1_4 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1804 wl_0_32 wl_1_32 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1837 wl_0_31 wl_1_31 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1859 wl_0_43 wl_1_43 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1848 wl_0_54 wl_1_54 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5131 wl_0_122 wl_1_122 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5120 wl_0_116 wl_1_116 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5142 wl_0_115 wl_1_115 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5175 wl_0_112 wl_1_112 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5153 wl_0_112 wl_1_112 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5164 wl_0_111 wl_1_111 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4430 wl_0_68 wl_1_68 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5186 wl_0_118 wl_1_118 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5197 wl_0_107 wl_1_107 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4441 wl_0_71 wl_1_71 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4463 wl_0_73 wl_1_73 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4452 wl_0_74 wl_1_74 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4474 wl_0_78 wl_1_78 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3762 wl_0_28 wl_1_28 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3751 wl_0_39 wl_1_39 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3740 wl_0_50 wl_1_50 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4496 wl_0_72 wl_1_72 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4485 wl_0_71 wl_1_71 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3773 wl_0_17 wl_1_17 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3784 wl_0_6 wl_1_6 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3795 wl_0_60 wl_1_60 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_519 wl_0_14 wl_1_14 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_508 wl_0_13 wl_1_13 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3014 wl_0_34 wl_1_34 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3003 wl_0_45 wl_1_45 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2302 wl_0_15 wl_1_15 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2313 wl_0_27 wl_1_27 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3025 wl_0_46 wl_1_46 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3047 wl_0_49 wl_1_49 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3058 wl_0_51 wl_1_51 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3036 wl_0_60 wl_1_60 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2324 wl_0_15 wl_1_15 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2346 wl_0_15 wl_1_15 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2335 wl_0_7 wl_1_7 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1601 wl_0_52 wl_1_52 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3069 wl_0_62 wl_1_62 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2357 wl_0_20 wl_1_20 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2368 wl_0_11 wl_1_11 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2379 wl_0_0 wl_1_0 bl_0_24 bl_1_24 br_0_24 br_1_24
+ sky130_fd_bd_sram__openram_dp_cell_2379/a_38_n79# vdd_uq2558 gnd sky130_fd_bd_sram__openram_dp_cell_2379/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1634 wl_0_53 wl_1_53 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1612 wl_0_57 wl_1_57 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1623 wl_0_60 wl_1_60 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1645 wl_0_60 wl_1_60 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1656 wl_0_49 wl_1_49 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1667 wl_0_54 wl_1_54 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1678 wl_0_59 wl_1_59 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1689 wl_0_48 wl_1_48 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4271 wl_0_67 wl_1_67 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4260 wl_0_78 wl_1_78 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4282 wl_0_80 wl_1_80 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3570 wl_0_50 wl_1_50 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4293 wl_0_93 wl_1_93 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3581 wl_0_55 wl_1_55 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3592 wl_0_62 wl_1_62 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2880 wl_0_38 wl_1_38 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2891 wl_0_43 wl_1_43 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7803 wl_0_95 wl_1_95 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7825 wl_0_63 wl_1_63 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7814 wl_0_64 wl_1_64 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7869 wl_0_63 wl_1_63 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7858 wl_0_64 wl_1_64 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7847 wl_0_63 wl_1_63 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7836 wl_0_64 wl_1_64 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_305 wl_0_21 wl_1_21 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_327 wl_0_21 wl_1_21 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_316 wl_0_20 wl_1_20 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_338 wl_0_24 wl_1_24 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_349 wl_0_22 wl_1_22 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2110 wl_0_7 wl_1_7 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2121 wl_0_6 wl_1_6 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2154 wl_0_20 wl_1_20 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2143 wl_0_18 wl_1_18 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2132 wl_0_13 wl_1_13 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1420 wl_0_40 wl_1_40 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2198 wl_0_24 wl_1_24 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2187 wl_0_24 wl_1_24 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2176 wl_0_18 wl_1_18 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2165 wl_0_29 wl_1_29 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1431 wl_0_36 wl_1_36 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1453 wl_0_36 wl_1_36 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1442 wl_0_40 wl_1_40 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1486 wl_0_36 wl_1_36 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1475 wl_0_36 wl_1_36 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1464 wl_0_38 wl_1_38 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1497 wl_0_46 wl_1_46 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_850 wl_0_24 wl_1_24 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_861 wl_0_16 wl_1_16 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_894 wl_0_16 wl_1_16 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_883 wl_0_8 wl_1_8 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_872 wl_0_5 wl_1_5 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4090 wl_0_92 wl_1_92 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6409 wl_0_69 wl_1_69 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5708 wl_0_95 wl_1_95 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5719 wl_0_121 wl_1_121 bl_0_16 bl_1_16 br_0_16
+ br_1_16 bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7600 wl_0_114 wl_1_114 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7622 wl_0_112 wl_1_112 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7611 wl_0_103 wl_1_103 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7633 wl_0_95 wl_1_95 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6932 wl_0_126 wl_1_126 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7666 wl_0_121 wl_1_121 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6921 wl_0_117 wl_1_117 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6910 wl_0_117 wl_1_117 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7677 wl_0_110 wl_1_110 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7644 wl_0_96 wl_1_96 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7655 wl_0_95 wl_1_95 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6965 wl_0_125 wl_1_125 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6954 wl_0_122 wl_1_122 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6943 wl_0_117 wl_1_117 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7688 wl_0_99 wl_1_99 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7699 wl_0_88 wl_1_88 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6987 wl_0_126 wl_1_126 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6998 wl_0_115 wl_1_115 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6976 wl_0_114 wl_1_114 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_102 wl_0_7 wl_1_7 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_113 wl_0_4 wl_1_4 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_146 wl_0_8 wl_1_8 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_135 wl_0_6 wl_1_6 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_124 wl_0_5 wl_1_5 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_157 wl_0_9 wl_1_9 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_168 wl_0_2 wl_1_2 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_179 wl_0_5 wl_1_5 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1261 wl_0_33 wl_1_33 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1250 wl_0_42 wl_1_42 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1294 wl_0_34 wl_1_34 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1283 wl_0_45 wl_1_45 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1272 wl_0_56 wl_1_56 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_680 wl_0_20 wl_1_20 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_691 wl_0_29 wl_1_29 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6217 wl_0_86 wl_1_86 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6206 wl_0_87 wl_1_87 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6228 wl_0_93 wl_1_93 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5516 wl_0_127 wl_1_127 bl_0_29 bl_1_29 br_0_29
+ br_1_29 sky130_fd_bd_sram__openram_dp_cell_5516/a_38_n79# vdd_uq2238 gnd sky130_fd_bd_sram__openram_dp_cell_5516/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5505 wl_0_121 wl_1_121 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6239 wl_0_82 wl_1_82 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5538 wl_0_122 wl_1_122 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5549 wl_0_117 wl_1_117 bl_0_25 bl_1_25 br_0_25
+ br_1_25 bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5527 wl_0_116 wl_1_116 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4804 wl_0_99 wl_1_99 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4826 wl_0_106 wl_1_106 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4837 wl_0_106 wl_1_106 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4848 wl_0_105 wl_1_105 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4815 wl_0_99 wl_1_99 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4859 wl_0_110 wl_1_110 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8120 wl_0_9 wl_1_9 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8153 wl_0_63 wl_1_63 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8142 wl_0_64 wl_1_64 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8131 wl_0_63 wl_1_63 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7430 wl_0_126 wl_1_126 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7452 wl_0_115 wl_1_115 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7441 wl_0_113 wl_1_113 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8186 wl_0_64 wl_1_64 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8175 wl_0_63 wl_1_63 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8164 wl_0_64 wl_1_64 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7474 wl_0_124 wl_1_124 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7485 wl_0_121 wl_1_121 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7463 wl_0_118 wl_1_118 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6740 wl_0_104 wl_1_104 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7496 wl_0_121 wl_1_121 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6773 wl_0_106 wl_1_106 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6762 wl_0_104 wl_1_104 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6751 wl_0_102 wl_1_102 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6784 wl_0_108 wl_1_108 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6795 wl_0_101 wl_1_101 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1080 wl_0_52 wl_1_52 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1091 wl_0_62 wl_1_62 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2709 wl_0_29 wl_1_29 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6003 wl_0_69 wl_1_69 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6014 wl_0_76 wl_1_76 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6036 wl_0_75 wl_1_75 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6025 wl_0_76 wl_1_76 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5302 wl_0_109 wl_1_109 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5313 wl_0_98 wl_1_98 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5324 wl_0_97 wl_1_97 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6058 wl_0_81 wl_1_81 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6069 wl_0_84 wl_1_84 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6047 wl_0_91 wl_1_91 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5357 wl_0_108 wl_1_108 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5335 wl_0_105 wl_1_105 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5346 wl_0_101 wl_1_101 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4601 wl_0_83 wl_1_83 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4612 wl_0_88 wl_1_88 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4623 wl_0_91 wl_1_91 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5368 wl_0_107 wl_1_107 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5379 wl_0_105 wl_1_105 bl_0_22 bl_1_22 br_0_22
+ br_1_22 bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3900 wl_0_32 wl_1_32 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3911 wl_0_66 wl_1_66 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4634 wl_0_84 wl_1_84 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4656 wl_0_86 wl_1_86 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4645 wl_0_91 wl_1_91 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3933 wl_0_67 wl_1_67 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3944 wl_0_74 wl_1_74 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3922 wl_0_74 wl_1_74 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4667 wl_0_85 wl_1_85 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4678 wl_0_86 wl_1_86 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4689 wl_0_91 wl_1_91 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3966 wl_0_66 wl_1_66 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3977 wl_0_66 wl_1_66 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3955 wl_0_68 wl_1_68 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3988 wl_0_73 wl_1_73 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3999 wl_0_69 wl_1_69 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7260 wl_0_106 wl_1_106 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7282 wl_0_106 wl_1_106 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7271 wl_0_99 wl_1_99 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7293 wl_0_97 wl_1_97 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6592 wl_0_86 wl_1_86 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6570 wl_0_90 wl_1_90 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6581 wl_0_91 wl_1_91 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5880 wl_0_76 wl_1_76 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5891 wl_0_65 wl_1_65 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3207 wl_0_55 wl_1_55 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3218 wl_0_47 wl_1_47 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3229 wl_0_52 wl_1_52 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2528 wl_0_13 wl_1_13 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2517 wl_0_11 wl_1_11 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2506 wl_0_2 wl_1_2 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1816 wl_0_19 wl_1_19 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2539 wl_0_13 wl_1_13 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1827 wl_0_8 wl_1_8 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1805 wl_0_31 wl_1_31 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1838 wl_0_32 wl_1_32 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1849 wl_0_53 wl_1_53 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5110 wl_0_126 wl_1_126 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5132 wl_0_121 wl_1_121 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5121 wl_0_115 wl_1_115 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5143 wl_0_127 wl_1_127 bl_0_10 bl_1_10 br_0_10
+ br_1_10 sky130_fd_bd_sram__openram_dp_cell_5143/a_38_n79# vdd_uq3454 gnd sky130_fd_bd_sram__openram_dp_cell_5143/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5165 wl_0_112 wl_1_112 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5176 wl_0_111 wl_1_111 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5154 wl_0_111 wl_1_111 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4420 wl_0_66 wl_1_66 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4431 wl_0_67 wl_1_67 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5187 wl_0_117 wl_1_117 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5198 wl_0_112 wl_1_112 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4464 wl_0_66 wl_1_66 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4442 wl_0_70 wl_1_70 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4453 wl_0_73 wl_1_73 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3763 wl_0_27 wl_1_27 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3752 wl_0_38 wl_1_38 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3741 wl_0_49 wl_1_49 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3730 wl_0_60 wl_1_60 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4486 wl_0_70 wl_1_70 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4497 wl_0_71 wl_1_71 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4475 wl_0_77 wl_1_77 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3774 wl_0_16 wl_1_16 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3785 wl_0_5 wl_1_5 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3796 wl_0_59 wl_1_59 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7090 wl_0_114 wl_1_114 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_509 wl_0_4 wl_1_4 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3015 wl_0_33 wl_1_33 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3004 wl_0_44 wl_1_44 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2303 wl_0_15 wl_1_15 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3026 wl_0_45 wl_1_45 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3048 wl_0_52 wl_1_52 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3037 wl_0_59 wl_1_59 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2325 wl_0_17 wl_1_17 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2336 wl_0_6 wl_1_6 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2314 wl_0_26 wl_1_26 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2347 wl_0_30 wl_1_30 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3059 wl_0_50 wl_1_50 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1602 wl_0_51 wl_1_51 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2358 wl_0_19 wl_1_19 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2369 wl_0_10 wl_1_10 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1635 wl_0_52 wl_1_52 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1613 wl_0_56 wl_1_56 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1624 wl_0_59 wl_1_59 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1668 wl_0_53 wl_1_53 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1657 wl_0_54 wl_1_54 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1646 wl_0_59 wl_1_59 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1679 wl_0_58 wl_1_58 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4272 wl_0_66 wl_1_66 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4261 wl_0_77 wl_1_77 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4250 wl_0_88 wl_1_88 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3571 wl_0_49 wl_1_49 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3560 wl_0_58 wl_1_58 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4283 wl_0_79 wl_1_79 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4294 wl_0_92 wl_1_92 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3582 wl_0_54 wl_1_54 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3593 wl_0_61 wl_1_61 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2870 wl_0_35 wl_1_35 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2881 wl_0_37 wl_1_37 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2892 wl_0_42 wl_1_42 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7804 wl_0_96 wl_1_96 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7826 wl_0_64 wl_1_64 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7815 wl_0_63 wl_1_63 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7859 wl_0_63 wl_1_63 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7848 wl_0_64 wl_1_64 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7837 wl_0_63 wl_1_63 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_306 wl_0_20 wl_1_20 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_317 wl_0_19 wl_1_19 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_328 wl_0_20 wl_1_20 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_339 wl_0_23 wl_1_23 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2111 wl_0_6 wl_1_6 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2100 wl_0_1 wl_1_1 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2122 wl_0_5 wl_1_5 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2155 wl_0_19 wl_1_19 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2144 wl_0_17 wl_1_17 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2133 wl_0_28 wl_1_28 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1410 wl_0_43 wl_1_43 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2188 wl_0_23 wl_1_23 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2177 wl_0_17 wl_1_17 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2166 wl_0_28 wl_1_28 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1432 wl_0_35 wl_1_35 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1421 wl_0_39 wl_1_39 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1443 wl_0_43 wl_1_43 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2199 wl_0_30 wl_1_30 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1487 wl_0_35 wl_1_35 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1454 wl_0_35 wl_1_35 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1476 wl_0_35 wl_1_35 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1465 wl_0_37 wl_1_37 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1498 wl_0_45 wl_1_45 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_840 wl_0_15 wl_1_15 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_851 wl_0_23 wl_1_23 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_862 wl_0_16 wl_1_16 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_884 wl_0_7 wl_1_7 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_873 wl_0_4 wl_1_4 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4091 wl_0_91 wl_1_91 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4080 wl_0_93 wl_1_93 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_895 wl_0_15 wl_1_15 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3390 wl_0_35 wl_1_35 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5709 wl_0_96 wl_1_96 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7601 wl_0_113 wl_1_113 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7623 wl_0_111 wl_1_111 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7612 wl_0_102 wl_1_102 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7634 wl_0_96 wl_1_96 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6911 wl_0_127 wl_1_127 bl_0_36 bl_1_36 br_0_36
+ br_1_36 sky130_fd_bd_sram__openram_dp_cell_6911/a_38_n79# vdd_uq1790 gnd sky130_fd_bd_sram__openram_dp_cell_6911/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7667 wl_0_120 wl_1_120 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6900 wl_0_119 wl_1_119 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6922 wl_0_116 wl_1_116 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7645 wl_0_95 wl_1_95 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7656 wl_0_96 wl_1_96 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6933 wl_0_127 wl_1_127 bl_0_35 bl_1_35 br_0_35
+ br_1_35 sky130_fd_bd_sram__openram_dp_cell_6933/a_38_n79# vdd_uq1854 gnd sky130_fd_bd_sram__openram_dp_cell_6933/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6966 wl_0_124 wl_1_124 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6955 wl_0_121 wl_1_121 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6944 wl_0_116 wl_1_116 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7678 wl_0_109 wl_1_109 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7689 wl_0_98 wl_1_98 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6988 wl_0_125 wl_1_125 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6999 wl_0_114 wl_1_114 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6977 wl_0_113 wl_1_113 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_103 wl_0_8 wl_1_8 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_125 wl_0_4 wl_1_4 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_114 wl_0_3 wl_1_3 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_136 wl_0_5 wl_1_5 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_147 wl_0_7 wl_1_7 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_158 wl_0_8 wl_1_8 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_169 wl_0_1 wl_1_1 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1251 wl_0_41 wl_1_41 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1262 wl_0_48 wl_1_48 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1240 wl_0_52 wl_1_52 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1295 wl_0_33 wl_1_33 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1284 wl_0_44 wl_1_44 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1273 wl_0_55 wl_1_55 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_670 wl_0_20 wl_1_20 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_692 wl_0_28 wl_1_28 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_681 wl_0_30 wl_1_30 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6218 wl_0_85 wl_1_85 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6207 wl_0_86 wl_1_86 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5506 wl_0_120 wl_1_120 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6229 wl_0_92 wl_1_92 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5517 wl_0_126 wl_1_126 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5539 wl_0_121 wl_1_121 bl_0_28 bl_1_28 br_0_28
+ br_1_28 bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5528 wl_0_115 wl_1_115 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4805 wl_0_98 wl_1_98 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4816 wl_0_110 wl_1_110 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4827 wl_0_105 wl_1_105 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4838 wl_0_98 wl_1_98 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4849 wl_0_97 wl_1_97 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8110 wl_0_19 wl_1_19 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8121 wl_0_8 wl_1_8 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8154 wl_0_64 wl_1_64 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8143 wl_0_63 wl_1_63 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8132 wl_0_64 wl_1_64 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7431 wl_0_127 wl_1_127 bl_0_51 bl_1_51 br_0_51
+ br_1_51 sky130_fd_bd_sram__openram_dp_cell_7431/a_38_n79# vdd_uq830 gnd sky130_fd_bd_sram__openram_dp_cell_7431/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7442 wl_0_118 wl_1_118 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7420 wl_0_117 wl_1_117 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8187 wl_0_63 wl_1_63 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8176 wl_0_64 wl_1_64 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8165 wl_0_63 wl_1_63 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7475 wl_0_123 wl_1_123 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7453 wl_0_118 wl_1_118 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7464 wl_0_117 wl_1_117 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6741 wl_0_103 wl_1_103 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6730 wl_0_98 wl_1_98 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7497 wl_0_127 wl_1_127 bl_0_61 bl_1_61 br_0_61
+ br_1_61 sky130_fd_bd_sram__openram_dp_cell_7497/a_38_n79# vdd_uq190 gnd sky130_fd_bd_sram__openram_dp_cell_7497/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7486 wl_0_124 wl_1_124 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6774 wl_0_105 wl_1_105 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6763 wl_0_103 wl_1_103 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6752 wl_0_101 wl_1_101 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6785 wl_0_107 wl_1_107 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6796 wl_0_100 wl_1_100 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1070 wl_0_58 wl_1_58 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1081 wl_0_51 wl_1_51 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1092 wl_0_61 wl_1_61 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6004 wl_0_68 wl_1_68 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6015 wl_0_75 wl_1_75 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6026 wl_0_75 wl_1_75 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5303 wl_0_108 wl_1_108 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5325 wl_0_99 wl_1_99 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5314 wl_0_97 wl_1_97 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6037 wl_0_72 wl_1_72 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6059 wl_0_90 wl_1_90 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6048 wl_0_90 wl_1_90 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5358 wl_0_107 wl_1_107 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5336 wl_0_104 wl_1_104 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5347 wl_0_100 wl_1_100 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4602 wl_0_82 wl_1_82 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4613 wl_0_87 wl_1_87 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5369 wl_0_106 wl_1_106 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3901 wl_0_31 wl_1_31 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3912 wl_0_65 wl_1_65 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4635 wl_0_83 wl_1_83 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4646 wl_0_90 wl_1_90 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4624 wl_0_94 wl_1_94 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3934 wl_0_66 wl_1_66 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3923 wl_0_73 wl_1_73 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3945 wl_0_78 wl_1_78 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4668 wl_0_84 wl_1_84 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4679 wl_0_85 wl_1_85 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4657 wl_0_85 wl_1_85 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3967 wl_0_65 wl_1_65 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3956 wl_0_67 wl_1_67 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3978 wl_0_78 wl_1_78 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3989 wl_0_72 wl_1_72 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7250 wl_0_106 wl_1_106 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7261 wl_0_109 wl_1_109 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7283 wl_0_105 wl_1_105 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7294 wl_0_100 wl_1_100 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7272 wl_0_98 wl_1_98 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6560 wl_0_84 wl_1_84 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6571 wl_0_89 wl_1_89 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6582 wl_0_90 wl_1_90 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5870 wl_0_70 wl_1_70 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5881 wl_0_75 wl_1_75 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6593 wl_0_85 wl_1_85 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5892 wl_0_74 wl_1_74 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3208 wl_0_54 wl_1_54 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3219 wl_0_62 wl_1_62 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2529 wl_0_12 wl_1_12 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2518 wl_0_10 wl_1_10 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2507 wl_0_4 wl_1_4 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1817 wl_0_18 wl_1_18 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1806 wl_0_29 wl_1_29 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1828 wl_0_7 wl_1_7 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1839 wl_0_31 wl_1_31 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5100 wl_0_119 wl_1_119 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5111 wl_0_125 wl_1_125 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5133 wl_0_120 wl_1_120 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5122 wl_0_114 wl_1_114 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5144 wl_0_126 wl_1_126 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5166 wl_0_111 wl_1_111 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5155 wl_0_112 wl_1_112 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4421 wl_0_65 wl_1_65 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4410 wl_0_75 wl_1_75 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5177 wl_0_127 wl_1_127 bl_0_8 bl_1_8 br_0_8 br_1_8
+ sky130_fd_bd_sram__openram_dp_cell_5177/a_38_n79# vdd_uq3582 gnd sky130_fd_bd_sram__openram_dp_cell_5177/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5188 wl_0_116 wl_1_116 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5199 wl_0_111 wl_1_111 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3720 wl_0_44 wl_1_44 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4465 wl_0_65 wl_1_65 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4443 wl_0_69 wl_1_69 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4454 wl_0_72 wl_1_72 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4432 wl_0_78 wl_1_78 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3753 wl_0_37 wl_1_37 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3742 wl_0_48 wl_1_48 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3731 wl_0_59 wl_1_59 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4498 wl_0_65 wl_1_65 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4487 wl_0_69 wl_1_69 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4476 wl_0_76 wl_1_76 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3775 wl_0_15 wl_1_15 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3786 wl_0_4 wl_1_4 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3764 wl_0_26 wl_1_26 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3797 wl_0_58 wl_1_58 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7080 wl_0_124 wl_1_124 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7091 wl_0_113 wl_1_113 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6390 wl_0_78 wl_1_78 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3005 wl_0_43 wl_1_43 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2304 wl_0_16 wl_1_16 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3027 wl_0_44 wl_1_44 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3016 wl_0_46 wl_1_46 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3049 wl_0_51 wl_1_51 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3038 wl_0_58 wl_1_58 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2326 wl_0_16 wl_1_16 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2337 wl_0_5 wl_1_5 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2315 wl_0_25 wl_1_25 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2359 wl_0_18 wl_1_18 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2348 wl_0_29 wl_1_29 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1603 wl_0_50 wl_1_50 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1636 wl_0_51 wl_1_51 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1614 wl_0_55 wl_1_55 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1625 wl_0_62 wl_1_62 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1669 wl_0_52 wl_1_52 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1658 wl_0_53 wl_1_53 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1647 wl_0_58 wl_1_58 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4240 wl_0_92 wl_1_92 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4273 wl_0_65 wl_1_65 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4262 wl_0_76 wl_1_76 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4251 wl_0_87 wl_1_87 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3561 wl_0_57 wl_1_57 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3550 wl_0_58 wl_1_58 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4284 wl_0_80 wl_1_80 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4295 wl_0_91 wl_1_91 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2860 wl_0_45 wl_1_45 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3583 wl_0_53 wl_1_53 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3594 wl_0_60 wl_1_60 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3572 wl_0_62 wl_1_62 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2871 wl_0_34 wl_1_34 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2882 wl_0_36 wl_1_36 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2893 wl_0_41 wl_1_41 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7805 wl_0_95 wl_1_95 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7816 wl_0_64 wl_1_64 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7849 wl_0_63 wl_1_63 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7838 wl_0_64 wl_1_64 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7827 wl_0_63 wl_1_63 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_307 wl_0_19 wl_1_19 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_329 wl_0_19 wl_1_19 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_318 wl_0_30 wl_1_30 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2101 wl_0_0 wl_1_0 bl_0_20 bl_1_20 br_0_20 br_1_20
+ sky130_fd_bd_sram__openram_dp_cell_2101/a_38_n79# vdd_uq2814 gnd sky130_fd_bd_sram__openram_dp_cell_2101/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2112 wl_0_5 wl_1_5 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2145 wl_0_19 wl_1_19 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2123 wl_0_4 wl_1_4 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2134 wl_0_27 wl_1_27 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1400 wl_0_33 wl_1_33 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1411 wl_0_42 wl_1_42 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2189 wl_0_22 wl_1_22 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2156 wl_0_18 wl_1_18 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2167 wl_0_27 wl_1_27 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2178 wl_0_30 wl_1_30 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1433 wl_0_34 wl_1_34 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1422 wl_0_38 wl_1_38 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1444 wl_0_42 wl_1_42 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1455 wl_0_34 wl_1_34 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1477 wl_0_34 wl_1_34 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1466 wl_0_36 wl_1_36 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1488 wl_0_38 wl_1_38 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1499 wl_0_44 wl_1_44 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_841 wl_0_14 wl_1_14 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_830 wl_0_25 wl_1_25 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_852 wl_0_22 wl_1_22 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_863 wl_0_15 wl_1_15 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_885 wl_0_6 wl_1_6 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_874 wl_0_3 wl_1_3 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4070 wl_0_72 wl_1_72 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4081 wl_0_89 wl_1_89 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_896 wl_0_16 wl_1_16 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4092 wl_0_84 wl_1_84 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3391 wl_0_34 wl_1_34 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3380 wl_0_34 wl_1_34 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2690 wl_0_27 wl_1_27 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7602 wl_0_112 wl_1_112 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7624 wl_0_112 wl_1_112 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7613 wl_0_101 wl_1_101 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6912 wl_0_126 wl_1_126 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6923 wl_0_124 wl_1_124 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7668 wl_0_119 wl_1_119 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6901 wl_0_118 wl_1_118 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7635 wl_0_95 wl_1_95 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7646 wl_0_96 wl_1_96 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7657 wl_0_95 wl_1_95 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6956 wl_0_127 wl_1_127 bl_0_34 bl_1_34 br_0_34
+ br_1_34 sky130_fd_bd_sram__openram_dp_cell_6956/a_38_n79# vdd_uq1918 gnd sky130_fd_bd_sram__openram_dp_cell_6956/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6934 wl_0_126 wl_1_126 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6945 wl_0_115 wl_1_115 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7679 wl_0_108 wl_1_108 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6989 wl_0_124 wl_1_124 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6967 wl_0_123 wl_1_123 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6978 wl_0_120 wl_1_120 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_104 wl_0_7 wl_1_7 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_126 wl_0_12 wl_1_12 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_115 wl_0_2 wl_1_2 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_137 wl_0_4 wl_1_4 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_159 wl_0_7 wl_1_7 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_148 wl_0_6 wl_1_6 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1252 wl_0_40 wl_1_40 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1241 wl_0_51 wl_1_51 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1230 wl_0_56 wl_1_56 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1285 wl_0_43 wl_1_43 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1263 wl_0_48 wl_1_48 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1274 wl_0_54 wl_1_54 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1296 wl_0_48 wl_1_48 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_671 wl_0_19 wl_1_19 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_693 wl_0_27 wl_1_27 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_682 wl_0_29 wl_1_29 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_660 wl_0_29 wl_1_29 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6208 wl_0_85 wl_1_85 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6219 wl_0_94 wl_1_94 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5507 wl_0_119 wl_1_119 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5518 wl_0_125 wl_1_125 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5529 wl_0_114 wl_1_114 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4817 wl_0_109 wl_1_109 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4828 wl_0_104 wl_1_104 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4839 wl_0_97 wl_1_97 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4806 wl_0_97 wl_1_97 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8111 wl_0_18 wl_1_18 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8100 wl_0_29 wl_1_29 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8122 wl_0_7 wl_1_7 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8144 wl_0_64 wl_1_64 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8133 wl_0_63 wl_1_63 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7432 wl_0_126 wl_1_126 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7421 wl_0_120 wl_1_120 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7443 wl_0_118 wl_1_118 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7410 wl_0_115 wl_1_115 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8177 wl_0_63 wl_1_63 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8166 wl_0_64 wl_1_64 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8155 wl_0_63 wl_1_63 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7476 wl_0_127 wl_1_127 bl_0_58 bl_1_58 br_0_58
+ br_1_58 sky130_fd_bd_sram__openram_dp_cell_7476/a_38_n79# vdd_uq382 gnd sky130_fd_bd_sram__openram_dp_cell_7476/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7465 wl_0_124 wl_1_124 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7454 wl_0_117 wl_1_117 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6731 wl_0_97 wl_1_97 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8188 wl_0_64 wl_1_64 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6720 wl_0_74 wl_1_74 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7498 wl_0_126 wl_1_126 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7487 wl_0_123 wl_1_123 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6742 wl_0_102 wl_1_102 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6764 wl_0_102 wl_1_102 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6753 wl_0_100 wl_1_100 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6786 wl_0_110 wl_1_110 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6775 wl_0_104 wl_1_104 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6797 wl_0_99 wl_1_99 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1060 wl_0_40 wl_1_40 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1082 wl_0_50 wl_1_50 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1071 wl_0_57 wl_1_57 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1093 wl_0_60 wl_1_60 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_490 wl_0_14 wl_1_14 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6005 wl_0_67 wl_1_67 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6016 wl_0_74 wl_1_74 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6027 wl_0_74 wl_1_74 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5304 wl_0_107 wl_1_107 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5315 wl_0_106 wl_1_106 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6038 wl_0_71 wl_1_71 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6049 wl_0_89 wl_1_89 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5348 wl_0_110 wl_1_110 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5337 wl_0_103 wl_1_103 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5326 wl_0_98 wl_1_98 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4603 wl_0_81 wl_1_81 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4614 wl_0_86 wl_1_86 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5359 wl_0_106 wl_1_106 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3902 wl_0_32 wl_1_32 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4636 wl_0_82 wl_1_82 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4647 wl_0_89 wl_1_89 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4625 wl_0_93 wl_1_93 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3935 wl_0_65 wl_1_65 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3924 wl_0_72 wl_1_72 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3913 wl_0_73 wl_1_73 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4658 wl_0_84 wl_1_84 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4669 wl_0_83 wl_1_83 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3957 wl_0_66 wl_1_66 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3968 wl_0_75 wl_1_75 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3946 wl_0_77 wl_1_77 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3979 wl_0_77 wl_1_77 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7251 wl_0_105 wl_1_105 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7240 wl_0_103 wl_1_103 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7262 wl_0_108 wl_1_108 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7284 wl_0_104 wl_1_104 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7273 wl_0_97 wl_1_97 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7295 wl_0_110 wl_1_110 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6572 wl_0_88 wl_1_88 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6583 wl_0_89 wl_1_89 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6561 wl_0_92 wl_1_92 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6550 wl_0_94 wl_1_94 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5860 wl_0_66 wl_1_66 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5871 wl_0_69 wl_1_69 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6594 wl_0_84 wl_1_84 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5893 wl_0_73 wl_1_73 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5882 wl_0_74 wl_1_74 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3209 wl_0_53 wl_1_53 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2519 wl_0_9 wl_1_9 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2508 wl_0_3 wl_1_3 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1818 wl_0_17 wl_1_17 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1807 wl_0_28 wl_1_28 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1829 wl_0_6 wl_1_6 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5112 wl_0_124 wl_1_124 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5101 wl_0_118 wl_1_118 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5123 wl_0_113 wl_1_113 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5145 wl_0_125 wl_1_125 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5134 wl_0_119 wl_1_119 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5167 wl_0_112 wl_1_112 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5156 wl_0_111 wl_1_111 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4400 wl_0_66 wl_1_66 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4422 wl_0_72 wl_1_72 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4411 wl_0_74 wl_1_74 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5178 wl_0_126 wl_1_126 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5189 wl_0_115 wl_1_115 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3710 wl_0_54 wl_1_54 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4444 wl_0_68 wl_1_68 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4455 wl_0_71 wl_1_71 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4433 wl_0_77 wl_1_77 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3754 wl_0_36 wl_1_36 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3721 wl_0_43 wl_1_43 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3743 wl_0_47 wl_1_47 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3732 wl_0_58 wl_1_58 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4488 wl_0_68 wl_1_68 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4466 wl_0_69 wl_1_69 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4477 wl_0_75 wl_1_75 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3776 wl_0_14 wl_1_14 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3787 wl_0_3 wl_1_3 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3765 wl_0_25 wl_1_25 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4499 wl_0_76 wl_1_76 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3798 wl_0_57 wl_1_57 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7081 wl_0_123 wl_1_123 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7070 wl_0_114 wl_1_114 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7092 wl_0_112 wl_1_112 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6380 wl_0_66 wl_1_66 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6391 wl_0_77 wl_1_77 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5690 wl_0_95 wl_1_95 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3006 wl_0_42 wl_1_42 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3028 wl_0_43 wl_1_43 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3017 wl_0_45 wl_1_45 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3039 wl_0_57 wl_1_57 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2316 wl_0_24 wl_1_24 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2305 wl_0_15 wl_1_15 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2327 wl_0_15 wl_1_15 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2338 wl_0_4 wl_1_4 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2349 wl_0_28 wl_1_28 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1604 wl_0_49 wl_1_49 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1615 wl_0_54 wl_1_54 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1626 wl_0_61 wl_1_61 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1637 wl_0_50 wl_1_50 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1648 wl_0_57 wl_1_57 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1659 wl_0_62 wl_1_62 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4230 wl_0_82 wl_1_82 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4263 wl_0_75 wl_1_75 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4252 wl_0_86 wl_1_86 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4241 wl_0_91 wl_1_91 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3562 wl_0_56 wl_1_56 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3551 wl_0_57 wl_1_57 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3540 wl_0_58 wl_1_58 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4274 wl_0_79 wl_1_79 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4285 wl_0_79 wl_1_79 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4296 wl_0_90 wl_1_90 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2850 wl_0_16 wl_1_16 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3584 wl_0_52 wl_1_52 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3595 wl_0_59 wl_1_59 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3573 wl_0_61 wl_1_61 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2883 wl_0_35 wl_1_35 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2894 wl_0_40 wl_1_40 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2861 wl_0_44 wl_1_44 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2872 wl_0_46 wl_1_46 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7806 wl_0_96 wl_1_96 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7817 wl_0_63 wl_1_63 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7839 wl_0_63 wl_1_63 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7828 wl_0_64 wl_1_64 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_308 wl_0_18 wl_1_18 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_319 wl_0_29 wl_1_29 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2113 wl_0_14 wl_1_14 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2102 wl_0_11 wl_1_11 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2124 wl_0_3 wl_1_3 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2135 wl_0_26 wl_1_26 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2146 wl_0_28 wl_1_28 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1401 wl_0_36 wl_1_36 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2157 wl_0_17 wl_1_17 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2168 wl_0_26 wl_1_26 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2179 wl_0_29 wl_1_29 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1423 wl_0_37 wl_1_37 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1412 wl_0_41 wl_1_41 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1434 wl_0_44 wl_1_44 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1456 wl_0_33 wl_1_33 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1478 wl_0_33 wl_1_33 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1467 wl_0_35 wl_1_35 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1445 wl_0_41 wl_1_41 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1489 wl_0_37 wl_1_37 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_820 wl_0_15 wl_1_15 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_842 wl_0_13 wl_1_13 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_831 wl_0_24 wl_1_24 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_853 wl_0_21 wl_1_21 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_864 wl_0_16 wl_1_16 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_875 wl_0_2 wl_1_2 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4060 wl_0_67 wl_1_67 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4071 wl_0_71 wl_1_71 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4082 wl_0_88 wl_1_88 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_897 wl_0_15 wl_1_15 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_886 wl_0_5 wl_1_5 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3370 wl_0_44 wl_1_44 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4093 wl_0_83 wl_1_83 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3392 wl_0_33 wl_1_33 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3381 wl_0_33 wl_1_33 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2680 wl_0_17 wl_1_17 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2691 wl_0_26 wl_1_26 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1990 wl_0_3 wl_1_3 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7603 wl_0_111 wl_1_111 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7625 wl_0_111 wl_1_111 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7614 wl_0_100 wl_1_100 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6913 wl_0_125 wl_1_125 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6902 wl_0_117 wl_1_117 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7636 wl_0_96 wl_1_96 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7647 wl_0_95 wl_1_95 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7658 wl_0_96 wl_1_96 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6957 wl_0_126 wl_1_126 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6935 wl_0_125 wl_1_125 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6924 wl_0_123 wl_1_123 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7669 wl_0_118 wl_1_118 bl_0_48 bl_1_48 br_0_48
+ br_1_48 bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6946 wl_0_114 wl_1_114 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6968 wl_0_122 wl_1_122 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6979 wl_0_119 wl_1_119 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_127 wl_0_14 wl_1_14 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_105 wl_0_13 wl_1_13 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_116 wl_0_1 wl_1_1 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_138 wl_0_10 wl_1_10 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_149 wl_0_5 wl_1_5 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1253 wl_0_39 wl_1_39 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1242 wl_0_50 wl_1_50 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1220 wl_0_54 wl_1_54 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1231 wl_0_55 wl_1_55 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1286 wl_0_42 wl_1_42 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1264 wl_0_47 wl_1_47 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1275 wl_0_53 wl_1_53 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1297 wl_0_47 wl_1_47 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_650 wl_0_24 wl_1_24 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_672 wl_0_18 wl_1_18 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_683 wl_0_28 wl_1_28 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_661 wl_0_28 wl_1_28 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_694 wl_0_19 wl_1_19 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6209 wl_0_84 wl_1_84 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5519 wl_0_124 wl_1_124 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5508 wl_0_118 wl_1_118 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4818 wl_0_108 wl_1_108 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4807 wl_0_105 wl_1_105 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4829 wl_0_103 wl_1_103 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8101 wl_0_28 wl_1_28 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7400 wl_0_120 wl_1_120 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8112 wl_0_17 wl_1_17 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8123 wl_0_6 wl_1_6 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8145 wl_0_63 wl_1_63 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8134 wl_0_64 wl_1_64 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7433 wl_0_125 wl_1_125 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7422 wl_0_119 wl_1_119 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7411 wl_0_114 wl_1_114 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8178 wl_0_64 wl_1_64 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8167 wl_0_63 wl_1_63 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8156 wl_0_64 wl_1_64 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7466 wl_0_123 wl_1_123 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7444 wl_0_118 wl_1_118 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7455 wl_0_116 wl_1_116 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6732 wl_0_101 wl_1_101 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8189 wl_0_63 wl_1_63 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6721 wl_0_73 wl_1_73 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6710 wl_0_84 wl_1_84 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7488 wl_0_127 wl_1_127 bl_0_62 bl_1_62 br_0_62
+ br_1_62 sky130_fd_bd_sram__openram_dp_cell_7488/a_38_n79# vdd_uq99 gnd sky130_fd_bd_sram__openram_dp_cell_7488/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7477 wl_0_126 wl_1_126 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7499 wl_0_125 wl_1_125 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6743 wl_0_101 wl_1_101 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6765 wl_0_101 wl_1_101 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6754 wl_0_99 wl_1_99 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6787 wl_0_109 wl_1_109 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6776 wl_0_103 wl_1_103 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6798 wl_0_98 wl_1_98 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1061 wl_0_39 wl_1_39 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1050 wl_0_41 wl_1_41 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1083 wl_0_49 wl_1_49 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1072 wl_0_56 wl_1_56 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1094 wl_0_59 wl_1_59 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_491 wl_0_13 wl_1_13 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_480 wl_0_3 wl_1_3 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6006 wl_0_66 wl_1_66 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6017 wl_0_73 wl_1_73 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5305 wl_0_106 wl_1_106 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5316 wl_0_105 wl_1_105 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6039 wl_0_70 wl_1_70 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6028 wl_0_73 wl_1_73 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5349 wl_0_109 wl_1_109 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5338 wl_0_102 wl_1_102 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5327 wl_0_97 wl_1_97 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4604 wl_0_84 wl_1_84 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3903 wl_0_31 wl_1_31 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4637 wl_0_81 wl_1_81 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4615 wl_0_85 wl_1_85 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4626 wl_0_92 wl_1_92 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3936 wl_0_65 wl_1_65 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3914 wl_0_72 wl_1_72 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3925 wl_0_71 wl_1_71 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4659 wl_0_83 wl_1_83 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4648 wl_0_88 wl_1_88 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3958 wl_0_65 wl_1_65 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3969 wl_0_74 wl_1_74 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3947 wl_0_76 wl_1_76 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7230 wl_0_104 wl_1_104 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7241 wl_0_102 wl_1_102 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7263 wl_0_107 wl_1_107 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7252 wl_0_104 wl_1_104 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7285 wl_0_103 wl_1_103 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7274 wl_0_104 wl_1_104 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6540 wl_0_88 wl_1_88 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7296 wl_0_109 wl_1_109 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6573 wl_0_87 wl_1_87 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6562 wl_0_91 wl_1_91 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6551 wl_0_93 wl_1_93 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5861 wl_0_65 wl_1_65 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6595 wl_0_83 wl_1_83 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6584 wl_0_94 wl_1_94 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5850 wl_0_95 wl_1_95 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5872 wl_0_68 wl_1_68 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5894 wl_0_72 wl_1_72 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5883 wl_0_73 wl_1_73 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2509 wl_0_5 wl_1_5 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1808 wl_0_27 wl_1_27 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1819 wl_0_16 wl_1_16 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5113 wl_0_123 wl_1_123 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5124 wl_0_118 wl_1_118 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5102 wl_0_117 wl_1_117 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5146 wl_0_124 wl_1_124 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5135 wl_0_118 wl_1_118 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5157 wl_0_112 wl_1_112 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4401 wl_0_65 wl_1_65 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4412 wl_0_73 wl_1_73 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5179 wl_0_125 wl_1_125 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5168 wl_0_111 wl_1_111 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3700 wl_0_34 wl_1_34 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3711 wl_0_53 wl_1_53 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4445 wl_0_67 wl_1_67 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4456 wl_0_70 wl_1_70 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4423 wl_0_71 wl_1_71 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4434 wl_0_78 wl_1_78 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3722 wl_0_32 wl_1_32 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3744 wl_0_46 wl_1_46 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3733 wl_0_57 wl_1_57 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4489 wl_0_67 wl_1_67 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4467 wl_0_68 wl_1_68 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4478 wl_0_78 wl_1_78 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3766 wl_0_24 wl_1_24 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3777 wl_0_13 wl_1_13 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3755 wl_0_35 wl_1_35 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3788 wl_0_2 wl_1_2 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3799 wl_0_56 wl_1_56 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7060 wl_0_124 wl_1_124 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7071 wl_0_126 wl_1_126 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7082 wl_0_122 wl_1_122 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7093 wl_0_111 wl_1_111 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6381 wl_0_65 wl_1_65 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6370 wl_0_76 wl_1_76 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6392 wl_0_76 wl_1_76 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5680 wl_0_95 wl_1_95 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5691 wl_0_96 wl_1_96 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4990 wl_0_127 wl_1_127 bl_0_0 bl_1_0 br_0_0 br_1_0
+ sky130_fd_bd_sram__openram_dp_cell_4990/a_38_n79# vdd_uq4094 gnd sky130_fd_bd_sram__openram_dp_cell_4990/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3007 wl_0_41 wl_1_41 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3029 wl_0_42 wl_1_42 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3018 wl_0_45 wl_1_45 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2317 wl_0_23 wl_1_23 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2306 wl_0_16 wl_1_16 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2328 wl_0_14 wl_1_14 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2339 wl_0_3 wl_1_3 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1605 wl_0_50 wl_1_50 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1616 wl_0_53 wl_1_53 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1627 wl_0_60 wl_1_60 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1638 wl_0_49 wl_1_49 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1649 wl_0_56 wl_1_56 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4231 wl_0_81 wl_1_81 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4220 wl_0_92 wl_1_92 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4264 wl_0_74 wl_1_74 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4242 wl_0_80 wl_1_80 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4253 wl_0_85 wl_1_85 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3530 wl_0_52 wl_1_52 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3552 wl_0_56 wl_1_56 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3541 wl_0_57 wl_1_57 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4286 wl_0_80 wl_1_80 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4275 wl_0_80 wl_1_80 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4297 wl_0_89 wl_1_89 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2840 wl_0_16 wl_1_16 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2851 wl_0_15 wl_1_15 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3585 wl_0_51 wl_1_51 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3563 wl_0_55 wl_1_55 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3596 wl_0_58 wl_1_58 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3574 wl_0_62 wl_1_62 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2884 wl_0_34 wl_1_34 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2862 wl_0_43 wl_1_43 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2873 wl_0_45 wl_1_45 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2895 wl_0_39 wl_1_39 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7807 wl_0_95 wl_1_95 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7829 wl_0_63 wl_1_63 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7818 wl_0_64 wl_1_64 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_309 wl_0_17 wl_1_17 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2103 wl_0_10 wl_1_10 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2114 wl_0_13 wl_1_13 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2125 wl_0_2 wl_1_2 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2136 wl_0_25 wl_1_25 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1402 wl_0_35 wl_1_35 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2158 wl_0_18 wl_1_18 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2169 wl_0_25 wl_1_25 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2147 wl_0_27 wl_1_27 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1424 wl_0_36 wl_1_36 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1413 wl_0_40 wl_1_40 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1435 wl_0_43 wl_1_43 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1446 wl_0_40 wl_1_40 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1468 wl_0_43 wl_1_43 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1457 wl_0_46 wl_1_46 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1479 wl_0_34 wl_1_34 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_821 wl_0_16 wl_1_16 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_832 wl_0_23 wl_1_23 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_810 wl_0_25 wl_1_25 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_854 wl_0_20 wl_1_20 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_865 wl_0_15 wl_1_15 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_843 wl_0_12 wl_1_12 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4061 wl_0_66 wl_1_66 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4072 wl_0_70 wl_1_70 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4050 wl_0_77 wl_1_77 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_898 wl_0_15 wl_1_15 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_876 wl_0_1 wl_1_1 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_887 wl_0_4 wl_1_4 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3360 wl_0_44 wl_1_44 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4094 wl_0_82 wl_1_82 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4083 wl_0_87 wl_1_87 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3382 wl_0_36 wl_1_36 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3371 wl_0_43 wl_1_43 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3393 wl_0_46 wl_1_46 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2681 wl_0_17 wl_1_17 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2670 wl_0_17 wl_1_17 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2692 wl_0_25 wl_1_25 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1980 wl_0_12 wl_1_12 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1991 wl_0_2 wl_1_2 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7604 wl_0_110 wl_1_110 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7615 wl_0_99 wl_1_99 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6914 wl_0_124 wl_1_124 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6903 wl_0_116 wl_1_116 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7626 wl_0_112 wl_1_112 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7637 wl_0_95 wl_1_95 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7648 wl_0_96 wl_1_96 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7659 wl_0_95 wl_1_95 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6936 wl_0_124 wl_1_124 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6925 wl_0_115 wl_1_115 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6947 wl_0_113 wl_1_113 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6958 wl_0_125 wl_1_125 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6969 wl_0_121 wl_1_121 bl_0_38 bl_1_38 br_0_38
+ br_1_38 bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_128 wl_0_13 wl_1_13 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_106 wl_0_12 wl_1_12 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_117 wl_0_0 wl_1_0 bl_0_53 bl_1_53 br_0_53 br_1_53
+ sky130_fd_bd_sram__openram_dp_cell_117/a_38_n79# vdd_uq702 gnd sky130_fd_bd_sram__openram_dp_cell_117/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_139 wl_0_9 wl_1_9 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1210 wl_0_55 wl_1_55 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1243 wl_0_49 wl_1_49 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1221 wl_0_53 wl_1_53 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1232 wl_0_54 wl_1_54 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1254 wl_0_38 wl_1_38 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1265 wl_0_47 wl_1_47 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1276 wl_0_52 wl_1_52 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1287 wl_0_41 wl_1_41 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1298 wl_0_48 wl_1_48 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_640 wl_0_0 wl_1_0 bl_0_33 bl_1_33 br_0_33 br_1_33
+ sky130_fd_bd_sram__openram_dp_cell_640/a_38_n79# vdd_uq1982 gnd sky130_fd_bd_sram__openram_dp_cell_640/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_673 wl_0_17 wl_1_17 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_651 wl_0_23 wl_1_23 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_684 wl_0_27 wl_1_27 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_662 wl_0_27 wl_1_27 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_695 wl_0_18 wl_1_18 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3190 wl_0_50 wl_1_50 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5509 wl_0_117 wl_1_117 bl_0_30 bl_1_30 br_0_30
+ br_1_30 bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4819 wl_0_107 wl_1_107 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4808 wl_0_104 wl_1_104 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8102 wl_0_27 wl_1_27 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8113 wl_0_16 wl_1_16 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8124 wl_0_5 wl_1_5 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8135 wl_0_63 wl_1_63 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7412 wl_0_127 wl_1_127 bl_0_52 bl_1_52 br_0_52
+ br_1_52 sky130_fd_bd_sram__openram_dp_cell_7412/a_38_n79# vdd_uq766 gnd sky130_fd_bd_sram__openram_dp_cell_7412/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7434 wl_0_124 wl_1_124 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7401 wl_0_119 wl_1_119 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7423 wl_0_118 wl_1_118 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8168 wl_0_64 wl_1_64 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8157 wl_0_63 wl_1_63 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8146 wl_0_64 wl_1_64 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7467 wl_0_122 wl_1_122 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7445 wl_0_117 wl_1_117 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7456 wl_0_115 wl_1_115 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8179 wl_0_63 wl_1_63 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6722 wl_0_72 wl_1_72 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6711 wl_0_83 wl_1_83 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6700 wl_0_94 wl_1_94 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7489 wl_0_126 wl_1_126 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7478 wl_0_125 wl_1_125 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6744 wl_0_100 wl_1_100 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6733 wl_0_100 wl_1_100 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6755 wl_0_98 wl_1_98 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6788 wl_0_108 wl_1_108 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6777 wl_0_102 wl_1_102 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6766 wl_0_100 wl_1_100 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6799 wl_0_97 wl_1_97 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1051 wl_0_40 wl_1_40 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1040 wl_0_44 wl_1_44 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1062 wl_0_38 wl_1_38 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1084 wl_0_53 wl_1_53 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1073 wl_0_55 wl_1_55 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1095 wl_0_58 wl_1_58 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7990 wl_0_11 wl_1_11 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_492 wl_0_12 wl_1_12 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_470 wl_0_1 wl_1_1 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_481 wl_0_2 wl_1_2 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6007 wl_0_65 wl_1_65 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6018 wl_0_72 wl_1_72 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5306 wl_0_105 wl_1_105 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6029 wl_0_78 wl_1_78 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5317 wl_0_104 wl_1_104 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5339 wl_0_101 wl_1_101 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5328 wl_0_98 wl_1_98 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4605 wl_0_94 wl_1_94 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4616 wl_0_84 wl_1_84 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4638 wl_0_90 wl_1_90 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4627 wl_0_91 wl_1_91 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3904 wl_0_32 wl_1_32 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3926 wl_0_70 wl_1_70 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3915 wl_0_71 wl_1_71 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4649 wl_0_87 wl_1_87 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3959 wl_0_73 wl_1_73 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3948 wl_0_75 wl_1_75 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3937 wl_0_78 wl_1_78 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7242 wl_0_110 wl_1_110 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7220 wl_0_103 wl_1_103 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7231 wl_0_103 wl_1_103 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7264 wl_0_106 wl_1_106 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7253 wl_0_103 wl_1_103 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7275 wl_0_103 wl_1_103 bl_0_49 bl_1_49 br_0_49
+ br_1_49 bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6530 wl_0_94 wl_1_94 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7297 wl_0_108 wl_1_108 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7286 wl_0_102 wl_1_102 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6574 wl_0_86 wl_1_86 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6541 wl_0_87 wl_1_87 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6563 wl_0_90 wl_1_90 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6552 wl_0_92 wl_1_92 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5840 wl_0_65 wl_1_65 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5862 wl_0_78 wl_1_78 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6596 wl_0_82 wl_1_82 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6585 wl_0_93 wl_1_93 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5851 wl_0_96 wl_1_96 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5873 wl_0_67 wl_1_67 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5895 wl_0_71 wl_1_71 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5884 wl_0_72 wl_1_72 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1809 wl_0_26 wl_1_26 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5114 wl_0_122 wl_1_122 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5103 wl_0_116 wl_1_116 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5147 wl_0_123 wl_1_123 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5136 wl_0_117 wl_1_117 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5125 wl_0_117 wl_1_117 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5158 wl_0_111 wl_1_111 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4413 wl_0_72 wl_1_72 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4402 wl_0_75 wl_1_75 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5169 wl_0_112 wl_1_112 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3701 wl_0_33 wl_1_33 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4446 wl_0_66 wl_1_66 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4424 wl_0_70 wl_1_70 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4435 wl_0_77 wl_1_77 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3723 wl_0_31 wl_1_31 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3745 wl_0_45 wl_1_45 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3712 wl_0_52 wl_1_52 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3734 wl_0_56 wl_1_56 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4468 wl_0_67 wl_1_67 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4457 wl_0_69 wl_1_69 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4479 wl_0_77 wl_1_77 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3767 wl_0_23 wl_1_23 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3778 wl_0_12 wl_1_12 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3756 wl_0_34 wl_1_34 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3789 wl_0_1 wl_1_1 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7050 wl_0_116 wl_1_116 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7072 wl_0_125 wl_1_125 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7061 wl_0_123 wl_1_123 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7083 wl_0_121 wl_1_121 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7094 wl_0_110 wl_1_110 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6382 wl_0_67 wl_1_67 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6360 wl_0_75 wl_1_75 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6371 wl_0_75 wl_1_75 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5670 wl_0_111 wl_1_111 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6393 wl_0_68 wl_1_68 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5681 wl_0_96 wl_1_96 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5692 wl_0_95 wl_1_95 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4991 wl_0_126 wl_1_126 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4980 wl_0_113 wl_1_113 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3008 wl_0_40 wl_1_40 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3019 wl_0_44 wl_1_44 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2318 wl_0_22 wl_1_22 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2307 wl_0_15 wl_1_15 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2329 wl_0_13 wl_1_13 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1606 wl_0_49 wl_1_49 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1617 wl_0_52 wl_1_52 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1639 wl_0_58 wl_1_58 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1628 wl_0_59 wl_1_59 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4210 wl_0_85 wl_1_85 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4221 wl_0_91 wl_1_91 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4243 wl_0_79 wl_1_79 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4254 wl_0_84 wl_1_84 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4232 wl_0_84 wl_1_84 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3531 wl_0_51 wl_1_51 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3553 wl_0_55 wl_1_55 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3542 wl_0_56 wl_1_56 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3520 wl_0_62 wl_1_62 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4265 wl_0_73 wl_1_73 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4287 wl_0_79 wl_1_79 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4276 wl_0_79 wl_1_79 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4298 wl_0_88 wl_1_88 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2841 wl_0_15 wl_1_15 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2830 wl_0_5 wl_1_5 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3586 wl_0_50 wl_1_50 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3564 wl_0_54 wl_1_54 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3575 wl_0_61 wl_1_61 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2885 wl_0_33 wl_1_33 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2863 wl_0_42 wl_1_42 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2874 wl_0_44 wl_1_44 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2852 wl_0_44 wl_1_44 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3597 wl_0_57 wl_1_57 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2896 wl_0_38 wl_1_38 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6190 wl_0_89 wl_1_89 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7808 wl_0_96 wl_1_96 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7819 wl_0_63 wl_1_63 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2104 wl_0_9 wl_1_9 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2137 wl_0_24 wl_1_24 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2115 wl_0_12 wl_1_12 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2126 wl_0_4 wl_1_4 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2159 wl_0_17 wl_1_17 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2148 wl_0_26 wl_1_26 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1403 wl_0_34 wl_1_34 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1425 wl_0_35 wl_1_35 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1414 wl_0_39 wl_1_39 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1447 wl_0_39 wl_1_39 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1436 wl_0_42 wl_1_42 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1469 wl_0_42 wl_1_42 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1458 wl_0_45 wl_1_45 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_833 wl_0_22 wl_1_22 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_822 wl_0_15 wl_1_15 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_811 wl_0_24 wl_1_24 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_800 wl_0_29 wl_1_29 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_855 wl_0_19 wl_1_19 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_866 wl_0_11 wl_1_11 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_844 wl_0_30 wl_1_30 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4062 wl_0_65 wl_1_65 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4040 wl_0_73 wl_1_73 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4051 wl_0_76 wl_1_76 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4073 wl_0_75 wl_1_75 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_877 wl_0_0 wl_1_0 bl_0_39 bl_1_39 br_0_39 br_1_39
+ sky130_fd_bd_sram__openram_dp_cell_877/a_38_n79# vdd_uq1598 gnd sky130_fd_bd_sram__openram_dp_cell_877/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_888 wl_0_3 wl_1_3 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_899 wl_0_33 wl_1_33 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3350 wl_0_42 wl_1_42 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3361 wl_0_43 wl_1_43 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4095 wl_0_81 wl_1_81 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4084 wl_0_86 wl_1_86 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3383 wl_0_35 wl_1_35 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3372 wl_0_42 wl_1_42 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3394 wl_0_45 wl_1_45 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2693 wl_0_24 wl_1_24 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2671 wl_0_18 wl_1_18 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2660 wl_0_17 wl_1_17 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2682 wl_0_27 wl_1_27 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1981 wl_0_11 wl_1_11 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1970 wl_0_2 wl_1_2 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1992 wl_0_1 wl_1_1 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7605 wl_0_109 wl_1_109 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7616 wl_0_98 wl_1_98 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6904 wl_0_115 wl_1_115 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7627 wl_0_111 wl_1_111 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7638 wl_0_96 wl_1_96 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7649 wl_0_95 wl_1_95 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6915 wl_0_123 wl_1_123 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6937 wl_0_123 wl_1_123 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6948 wl_0_115 wl_1_115 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6926 wl_0_114 wl_1_114 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6959 wl_0_124 wl_1_124 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_107 wl_0_11 wl_1_11 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_118 wl_0_3 wl_1_3 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_129 wl_0_12 wl_1_12 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1200 wl_0_53 wl_1_53 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1244 wl_0_48 wl_1_48 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1222 wl_0_52 wl_1_52 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1233 wl_0_53 wl_1_53 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1211 wl_0_54 wl_1_54 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1255 wl_0_48 wl_1_48 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1277 wl_0_51 wl_1_51 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1266 wl_0_62 wl_1_62 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1288 wl_0_40 wl_1_40 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1299 wl_0_47 wl_1_47 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_630 wl_0_7 wl_1_7 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_641 wl_0_4 wl_1_4 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_652 wl_0_22 wl_1_22 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_674 wl_0_22 wl_1_22 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_663 wl_0_26 wl_1_26 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_696 wl_0_17 wl_1_17 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_685 wl_0_26 wl_1_26 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3191 wl_0_49 wl_1_49 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3180 wl_0_52 wl_1_52 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2490 wl_0_4 wl_1_4 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4809 wl_0_98 wl_1_98 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8114 wl_0_15 wl_1_15 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8125 wl_0_4 wl_1_4 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8103 wl_0_26 wl_1_26 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8136 wl_0_64 wl_1_64 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7413 wl_0_126 wl_1_126 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7402 wl_0_120 wl_1_120 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7424 wl_0_117 wl_1_117 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8169 wl_0_63 wl_1_63 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8158 wl_0_64 wl_1_64 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8147 wl_0_63 wl_1_63 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7446 wl_0_116 wl_1_116 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7435 wl_0_114 wl_1_114 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7457 wl_0_114 wl_1_114 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6723 wl_0_71 wl_1_71 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6712 wl_0_82 wl_1_82 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6701 wl_0_93 wl_1_93 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7479 wl_0_127 wl_1_127 bl_0_63 bl_1_63 br_0_63
+ br_1_63 sky130_fd_bd_sram__openram_dp_cell_7479/a_38_n79# vdd gnd sky130_fd_bd_sram__openram_dp_cell_7479/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7468 wl_0_121 wl_1_121 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6734 wl_0_110 wl_1_110 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6745 wl_0_99 wl_1_99 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6756 wl_0_97 wl_1_97 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6767 wl_0_110 wl_1_110 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6789 wl_0_107 wl_1_107 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6778 wl_0_101 wl_1_101 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1030 wl_0_33 wl_1_33 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1041 wl_0_36 wl_1_36 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1052 wl_0_39 wl_1_39 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1063 wl_0_37 wl_1_37 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1085 wl_0_52 wl_1_52 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1074 wl_0_54 wl_1_54 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1096 wl_0_57 wl_1_57 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7980 wl_0_21 wl_1_21 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7991 wl_0_10 wl_1_10 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_460 wl_0_16 wl_1_16 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_482 wl_0_1 wl_1_1 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_471 wl_0_2 wl_1_2 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_493 wl_0_4 wl_1_4 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6008 wl_0_67 wl_1_67 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5307 wl_0_104 wl_1_104 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6019 wl_0_71 wl_1_71 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5318 wl_0_103 wl_1_103 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5329 wl_0_97 wl_1_97 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4617 wl_0_83 wl_1_83 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4628 wl_0_90 wl_1_90 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4606 wl_0_94 wl_1_94 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3905 wl_0_31 wl_1_31 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3927 wl_0_69 wl_1_69 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3916 wl_0_70 wl_1_70 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4639 wl_0_89 wl_1_89 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3949 wl_0_74 wl_1_74 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3938 wl_0_77 wl_1_77 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7210 wl_0_110 wl_1_110 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7221 wl_0_102 wl_1_102 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7232 wl_0_102 wl_1_102 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7243 wl_0_109 wl_1_109 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7265 wl_0_105 wl_1_105 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7254 wl_0_102 wl_1_102 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7276 wl_0_97 wl_1_97 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6520 wl_0_90 wl_1_90 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6531 wl_0_93 wl_1_93 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7298 wl_0_107 wl_1_107 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7287 wl_0_101 wl_1_101 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6542 wl_0_86 wl_1_86 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6553 wl_0_91 wl_1_91 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6564 wl_0_94 wl_1_94 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5830 wl_0_75 wl_1_75 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6597 wl_0_81 wl_1_81 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6575 wl_0_85 wl_1_85 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6586 wl_0_92 wl_1_92 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5852 wl_0_95 wl_1_95 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5841 wl_0_96 wl_1_96 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5874 wl_0_66 wl_1_66 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5896 wl_0_70 wl_1_70 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5885 wl_0_71 wl_1_71 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5863 wl_0_77 wl_1_77 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_290 wl_0_30 wl_1_30 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5115 wl_0_121 wl_1_121 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5104 wl_0_115 wl_1_115 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5126 wl_0_127 wl_1_127 bl_0_11 bl_1_11 br_0_11
+ br_1_11 sky130_fd_bd_sram__openram_dp_cell_5126/a_38_n79# vdd_uq3390 gnd sky130_fd_bd_sram__openram_dp_cell_5126/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5148 wl_0_122 wl_1_122 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5137 wl_0_116 wl_1_116 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4403 wl_0_74 wl_1_74 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5159 wl_0_112 wl_1_112 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3702 wl_0_62 wl_1_62 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4447 wl_0_65 wl_1_65 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4425 wl_0_69 wl_1_69 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4414 wl_0_71 wl_1_71 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4436 wl_0_76 wl_1_76 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3724 wl_0_32 wl_1_32 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3713 wl_0_51 wl_1_51 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3735 wl_0_55 wl_1_55 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4469 wl_0_66 wl_1_66 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4458 wl_0_68 wl_1_68 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3768 wl_0_22 wl_1_22 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3757 wl_0_33 wl_1_33 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3746 wl_0_44 wl_1_44 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3779 wl_0_11 wl_1_11 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7040 wl_0_126 wl_1_126 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7051 wl_0_115 wl_1_115 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7062 wl_0_122 wl_1_122 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7084 wl_0_120 wl_1_120 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7073 wl_0_113 wl_1_113 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7095 wl_0_109 wl_1_109 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6350 wl_0_67 wl_1_67 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6361 wl_0_74 wl_1_74 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6372 wl_0_74 wl_1_74 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5671 wl_0_112 wl_1_112 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5660 wl_0_101 wl_1_101 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6383 wl_0_66 wl_1_66 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6394 wl_0_67 wl_1_67 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5682 wl_0_95 wl_1_95 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5693 wl_0_96 wl_1_96 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4992 wl_0_125 wl_1_125 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4981 wl_0_114 wl_1_114 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4970 wl_0_113 wl_1_113 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3009 wl_0_39 wl_1_39 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2319 wl_0_21 wl_1_21 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2308 wl_0_30 wl_1_30 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1618 wl_0_51 wl_1_51 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1607 wl_0_62 wl_1_62 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1629 wl_0_58 wl_1_58 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4211 wl_0_84 wl_1_84 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4200 wl_0_88 wl_1_88 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4222 wl_0_90 wl_1_90 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3510 wl_0_54 wl_1_54 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4255 wl_0_83 wl_1_83 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4233 wl_0_83 wl_1_83 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4244 wl_0_94 wl_1_94 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3532 wl_0_50 wl_1_50 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3543 wl_0_55 wl_1_55 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3521 wl_0_61 wl_1_61 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4266 wl_0_72 wl_1_72 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4277 wl_0_79 wl_1_79 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4288 wl_0_80 wl_1_80 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2842 wl_0_16 wl_1_16 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2820 wl_0_15 wl_1_15 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2831 wl_0_4 wl_1_4 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3587 wl_0_49 wl_1_49 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3554 wl_0_52 wl_1_52 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3565 wl_0_53 wl_1_53 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3576 wl_0_60 wl_1_60 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4299 wl_0_87 wl_1_87 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2864 wl_0_41 wl_1_41 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2875 wl_0_43 wl_1_43 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2853 wl_0_43 wl_1_43 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3598 wl_0_56 wl_1_56 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2886 wl_0_33 wl_1_33 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2897 wl_0_37 wl_1_37 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6180 wl_0_87 wl_1_87 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6191 wl_0_94 wl_1_94 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5490 wl_0_126 wl_1_126 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7809 wl_0_95 wl_1_95 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2116 wl_0_11 wl_1_11 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2105 wl_0_8 wl_1_8 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2127 wl_0_3 wl_1_3 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2138 wl_0_23 wl_1_23 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2149 wl_0_25 wl_1_25 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1404 wl_0_33 wl_1_33 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1426 wl_0_34 wl_1_34 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1415 wl_0_38 wl_1_38 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1448 wl_0_38 wl_1_38 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1459 wl_0_44 wl_1_44 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1437 wl_0_46 wl_1_46 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_823 wl_0_16 wl_1_16 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_812 wl_0_23 wl_1_23 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_801 wl_0_28 wl_1_28 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4030 wl_0_77 wl_1_77 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_834 wl_0_21 wl_1_21 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_856 wl_0_18 wl_1_18 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_845 wl_0_29 wl_1_29 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4041 wl_0_72 wl_1_72 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4052 wl_0_75 wl_1_75 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4063 wl_0_76 wl_1_76 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_878 wl_0_13 wl_1_13 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_867 wl_0_10 wl_1_10 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_889 wl_0_2 wl_1_2 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3351 wl_0_41 wl_1_41 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3340 wl_0_44 wl_1_44 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4085 wl_0_85 wl_1_85 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4074 wl_0_86 wl_1_86 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4096 wl_0_90 wl_1_90 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2650 wl_0_20 wl_1_20 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3384 wl_0_34 wl_1_34 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3373 wl_0_41 wl_1_41 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3362 wl_0_42 wl_1_42 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3395 wl_0_44 wl_1_44 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2661 wl_0_22 wl_1_22 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2672 wl_0_17 wl_1_17 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2683 wl_0_29 wl_1_29 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2694 wl_0_23 wl_1_23 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1982 wl_0_11 wl_1_11 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1960 wl_0_6 wl_1_6 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1971 wl_0_1 wl_1_1 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1993 wl_0_0 wl_1_0 bl_0_30 bl_1_30 br_0_30 br_1_30
+ sky130_fd_bd_sram__openram_dp_cell_1993/a_38_n79# vdd_uq2174 gnd sky130_fd_bd_sram__openram_dp_cell_1993/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7606 wl_0_108 wl_1_108 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6905 wl_0_114 wl_1_114 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7617 wl_0_97 wl_1_97 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7628 wl_0_96 wl_1_96 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7639 wl_0_95 wl_1_95 bl_0_58 bl_1_58 br_0_58 br_1_58
+ bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6916 wl_0_122 wl_1_122 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6938 wl_0_122 wl_1_122 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6927 wl_0_113 wl_1_113 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6949 wl_0_117 wl_1_117 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_108 wl_0_10 wl_1_10 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_119 wl_0_2 wl_1_2 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1201 wl_0_49 wl_1_49 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1234 wl_0_52 wl_1_52 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1223 wl_0_51 wl_1_51 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1212 wl_0_53 wl_1_53 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1245 wl_0_47 wl_1_47 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1256 wl_0_47 wl_1_47 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1267 wl_0_61 wl_1_61 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1289 wl_0_39 wl_1_39 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1278 wl_0_50 wl_1_50 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_620 wl_0_9 wl_1_9 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_631 wl_0_6 wl_1_6 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_653 wl_0_21 wl_1_21 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_675 wl_0_21 wl_1_21 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_642 wl_0_3 wl_1_3 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_664 wl_0_25 wl_1_25 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_686 wl_0_25 wl_1_25 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_697 wl_0_26 wl_1_26 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3170 wl_0_62 wl_1_62 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3181 wl_0_51 wl_1_51 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3192 wl_0_53 wl_1_53 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2480 wl_0_0 wl_1_0 bl_0_6 bl_1_6 br_0_6 br_1_6
+ sky130_fd_bd_sram__openram_dp_cell_2480/a_38_n79# vdd_uq3710 gnd sky130_fd_bd_sram__openram_dp_cell_2480/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2491 wl_0_1 wl_1_1 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1790 wl_0_43 wl_1_43 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8115 wl_0_14 wl_1_14 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8126 wl_0_3 wl_1_3 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8104 wl_0_25 wl_1_25 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7414 wl_0_125 wl_1_125 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7403 wl_0_119 wl_1_119 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7425 wl_0_116 wl_1_116 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8159 wl_0_63 wl_1_63 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8148 wl_0_64 wl_1_64 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8137 wl_0_63 wl_1_63 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7447 wl_0_115 wl_1_115 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7436 wl_0_113 wl_1_113 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7458 wl_0_113 wl_1_113 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6713 wl_0_81 wl_1_81 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6702 wl_0_92 wl_1_92 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7469 wl_0_126 wl_1_126 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6735 wl_0_109 wl_1_109 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6746 wl_0_98 wl_1_98 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6724 wl_0_70 wl_1_70 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6768 wl_0_110 wl_1_110 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6757 wl_0_109 wl_1_109 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6779 wl_0_100 wl_1_100 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1042 wl_0_35 wl_1_35 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1031 wl_0_40 wl_1_40 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1020 wl_0_40 wl_1_40 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1064 wl_0_36 wl_1_36 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1053 wl_0_38 wl_1_38 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1086 wl_0_51 wl_1_51 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1075 wl_0_53 wl_1_53 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1097 wl_0_62 wl_1_62 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7970 wl_0_31 wl_1_31 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7981 wl_0_20 wl_1_20 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7992 wl_0_9 wl_1_9 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_450 wl_0_4 wl_1_4 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_461 wl_0_15 wl_1_15 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_472 wl_0_1 wl_1_1 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_483 wl_0_0 wl_1_0 bl_0_43 bl_1_43 br_0_43 br_1_43
+ sky130_fd_bd_sram__openram_dp_cell_483/a_38_n79# vdd_uq1342 gnd sky130_fd_bd_sram__openram_dp_cell_483/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_494 wl_0_3 wl_1_3 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6009 wl_0_66 wl_1_66 bl_0_52 bl_1_52 br_0_52 br_1_52
+ bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5308 wl_0_103 wl_1_103 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5319 wl_0_102 wl_1_102 bl_0_27 bl_1_27 br_0_27
+ br_1_27 bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4618 wl_0_82 wl_1_82 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4629 wl_0_89 wl_1_89 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4607 wl_0_93 wl_1_93 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3917 wl_0_69 wl_1_69 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3906 wl_0_71 wl_1_71 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3928 wl_0_68 wl_1_68 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3939 wl_0_76 wl_1_76 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7233 wl_0_110 wl_1_110 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7211 wl_0_109 wl_1_109 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7200 wl_0_105 wl_1_105 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7222 wl_0_101 wl_1_101 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7244 wl_0_108 wl_1_108 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7266 wl_0_104 wl_1_104 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7255 wl_0_101 wl_1_101 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6510 wl_0_82 wl_1_82 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6521 wl_0_89 wl_1_89 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7299 wl_0_106 wl_1_106 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7288 wl_0_100 wl_1_100 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7277 wl_0_98 wl_1_98 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5820 wl_0_85 wl_1_85 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6543 wl_0_85 wl_1_85 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6554 wl_0_90 wl_1_90 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6532 wl_0_92 wl_1_92 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6565 wl_0_93 wl_1_93 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5831 wl_0_74 wl_1_74 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6576 wl_0_84 wl_1_84 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6598 wl_0_88 wl_1_88 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6587 wl_0_91 wl_1_91 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5853 wl_0_96 wl_1_96 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5842 wl_0_95 wl_1_95 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5875 wl_0_65 wl_1_65 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5886 wl_0_70 wl_1_70 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5864 wl_0_76 wl_1_76 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5897 wl_0_69 wl_1_69 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_280 wl_0_28 wl_1_28 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_291 wl_0_29 wl_1_29 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5105 wl_0_114 wl_1_114 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5127 wl_0_126 wl_1_126 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5149 wl_0_121 wl_1_121 bl_0_10 bl_1_10 br_0_10
+ br_1_10 bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5116 wl_0_120 wl_1_120 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5138 wl_0_115 wl_1_115 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4404 wl_0_73 wl_1_73 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4426 wl_0_68 wl_1_68 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4415 wl_0_70 wl_1_70 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4437 wl_0_75 wl_1_75 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3725 wl_0_31 wl_1_31 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3714 wl_0_50 wl_1_50 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3736 wl_0_54 wl_1_54 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3703 wl_0_61 wl_1_61 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4459 wl_0_67 wl_1_67 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4448 wl_0_78 wl_1_78 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3769 wl_0_21 wl_1_21 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3758 wl_0_32 wl_1_32 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3747 wl_0_43 wl_1_43 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7041 wl_0_125 wl_1_125 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7030 wl_0_118 wl_1_118 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7074 wl_0_124 wl_1_124 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7063 wl_0_121 wl_1_121 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7052 wl_0_114 wl_1_114 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7085 wl_0_119 wl_1_119 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7096 wl_0_108 wl_1_108 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6351 wl_0_66 wl_1_66 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6362 wl_0_73 wl_1_73 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6373 wl_0_73 wl_1_73 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6340 wl_0_77 wl_1_77 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5650 wl_0_111 wl_1_111 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5661 wl_0_100 wl_1_100 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6395 wl_0_65 wl_1_65 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6384 wl_0_65 wl_1_65 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4960 wl_0_115 wl_1_115 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5672 wl_0_111 wl_1_111 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5683 wl_0_96 wl_1_96 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5694 wl_0_95 wl_1_95 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4993 wl_0_127 wl_1_127 bl_0_1 bl_1_1 br_0_1 br_1_1
+ sky130_fd_bd_sram__openram_dp_cell_4993/a_38_n79# vdd_uq4030 gnd sky130_fd_bd_sram__openram_dp_cell_4993/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4982 wl_0_118 wl_1_118 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4971 wl_0_116 wl_1_116 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2309 wl_0_16 wl_1_16 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1608 wl_0_61 wl_1_61 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1619 wl_0_50 wl_1_50 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4212 wl_0_83 wl_1_83 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4201 wl_0_94 wl_1_94 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3500 wl_0_50 wl_1_50 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4234 wl_0_82 wl_1_82 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4223 wl_0_89 wl_1_89 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4245 wl_0_93 wl_1_93 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3533 wl_0_49 wl_1_49 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3511 wl_0_53 wl_1_53 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3544 wl_0_54 wl_1_54 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3522 wl_0_60 wl_1_60 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4267 wl_0_71 wl_1_71 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4289 wl_0_79 wl_1_79 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4278 wl_0_80 wl_1_80 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4256 wl_0_82 wl_1_82 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2821 wl_0_14 wl_1_14 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2810 wl_0_9 wl_1_9 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2832 wl_0_3 wl_1_3 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3555 wl_0_51 wl_1_51 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3566 wl_0_52 wl_1_52 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3577 wl_0_59 wl_1_59 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2843 wl_0_15 wl_1_15 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2865 wl_0_40 wl_1_40 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2876 wl_0_42 wl_1_42 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2854 wl_0_42 wl_1_42 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3599 wl_0_55 wl_1_55 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3588 wl_0_60 wl_1_60 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2898 wl_0_36 wl_1_36 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2887 wl_0_40 wl_1_40 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6181 wl_0_86 wl_1_86 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6170 wl_0_91 wl_1_91 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6192 wl_0_93 wl_1_93 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5491 wl_0_125 wl_1_125 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5480 wl_0_117 wl_1_117 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4790 wl_0_105 wl_1_105 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2117 wl_0_10 wl_1_10 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2106 wl_0_7 wl_1_7 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2128 wl_0_2 wl_1_2 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2139 wl_0_22 wl_1_22 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1416 wl_0_37 wl_1_37 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1405 wl_0_40 wl_1_40 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1427 wl_0_33 wl_1_33 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1438 wl_0_45 wl_1_45 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1449 wl_0_46 wl_1_46 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_813 wl_0_16 wl_1_16 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_824 wl_0_15 wl_1_15 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_802 wl_0_27 wl_1_27 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4020 wl_0_68 wl_1_68 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_835 wl_0_20 wl_1_20 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_857 wl_0_17 wl_1_17 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_846 wl_0_28 wl_1_28 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4042 wl_0_71 wl_1_71 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4053 wl_0_74 wl_1_74 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4064 wl_0_78 wl_1_78 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4031 wl_0_78 wl_1_78 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_879 wl_0_12 wl_1_12 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_868 wl_0_9 wl_1_9 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3352 wl_0_40 wl_1_40 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3330 wl_0_44 wl_1_44 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3341 wl_0_43 wl_1_43 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4086 wl_0_84 wl_1_84 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4075 wl_0_85 wl_1_85 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4097 wl_0_89 wl_1_89 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2640 wl_0_30 wl_1_30 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3385 wl_0_33 wl_1_33 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3374 wl_0_40 wl_1_40 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3363 wl_0_41 wl_1_41 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2673 wl_0_24 wl_1_24 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2662 wl_0_21 wl_1_21 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2651 wl_0_19 wl_1_19 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2684 wl_0_28 wl_1_28 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3396 wl_0_43 wl_1_43 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2695 wl_0_22 wl_1_22 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1972 wl_0_0 wl_1_0 bl_0_26 bl_1_26 br_0_26 br_1_26
+ sky130_fd_bd_sram__openram_dp_cell_1972/a_38_n79# vdd_uq2430 gnd sky130_fd_bd_sram__openram_dp_cell_1972/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1961 wl_0_5 wl_1_5 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1950 wl_0_31 wl_1_31 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1983 wl_0_10 wl_1_10 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1994 wl_0_10 wl_1_10 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7607 wl_0_107 wl_1_107 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7618 wl_0_112 wl_1_112 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7629 wl_0_95 wl_1_95 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6917 wl_0_121 wl_1_121 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6939 wl_0_121 wl_1_121 bl_0_35 bl_1_35 br_0_35
+ br_1_35 bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6928 wl_0_114 wl_1_114 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6906 wl_0_113 wl_1_113 bl_0_37 bl_1_37 br_0_37
+ br_1_37 bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_109 wl_0_9 wl_1_9 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1235 wl_0_48 wl_1_48 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1202 wl_0_52 wl_1_52 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1213 wl_0_52 wl_1_52 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1224 wl_0_62 wl_1_62 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1257 wl_0_37 wl_1_37 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1246 wl_0_46 wl_1_46 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1268 wl_0_60 wl_1_60 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1279 wl_0_49 wl_1_49 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_621 wl_0_8 wl_1_8 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_610 wl_0_1 wl_1_1 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_632 wl_0_5 wl_1_5 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_654 wl_0_20 wl_1_20 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_643 wl_0_13 wl_1_13 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_665 wl_0_24 wl_1_24 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_676 wl_0_18 wl_1_18 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_687 wl_0_24 wl_1_24 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_698 wl_0_25 wl_1_25 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3160 wl_0_55 wl_1_55 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3182 wl_0_50 wl_1_50 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3193 wl_0_52 wl_1_52 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3171 wl_0_61 wl_1_61 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2470 wl_0_0 wl_1_0 bl_0_13 bl_1_13 br_0_13 br_1_13
+ sky130_fd_bd_sram__openram_dp_cell_2470/a_38_n79# vdd_uq3262 gnd sky130_fd_bd_sram__openram_dp_cell_2470/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2492 wl_0_0 wl_1_0 bl_0_2 bl_1_2 br_0_2 br_1_2
+ sky130_fd_bd_sram__openram_dp_cell_2492/a_38_n79# vdd_uq3966 gnd sky130_fd_bd_sram__openram_dp_cell_2492/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2481 wl_0_3 wl_1_3 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1780 wl_0_53 wl_1_53 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1791 wl_0_42 wl_1_42 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8105 wl_0_24 wl_1_24 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8116 wl_0_13 wl_1_13 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8127 wl_0_2 wl_1_2 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7415 wl_0_124 wl_1_124 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7404 wl_0_118 wl_1_118 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8149 wl_0_63 wl_1_63 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8138 wl_0_64 wl_1_64 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7437 wl_0_117 wl_1_117 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7426 wl_0_115 wl_1_115 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7448 wl_0_114 wl_1_114 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6714 wl_0_80 wl_1_80 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6703 wl_0_91 wl_1_91 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7459 wl_0_114 wl_1_114 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6736 wl_0_108 wl_1_108 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6747 wl_0_97 wl_1_97 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6725 wl_0_69 wl_1_69 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6769 wl_0_110 wl_1_110 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6758 wl_0_108 wl_1_108 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1010 wl_0_34 wl_1_34 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1043 wl_0_34 wl_1_34 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1032 wl_0_39 wl_1_39 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1021 wl_0_39 wl_1_39 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1054 wl_0_33 wl_1_33 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1065 wl_0_46 wl_1_46 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1076 wl_0_52 wl_1_52 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1087 wl_0_50 wl_1_50 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1098 wl_0_56 wl_1_56 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7971 wl_0_30 wl_1_30 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7960 wl_0_41 wl_1_41 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7982 wl_0_19 wl_1_19 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7993 wl_0_8 wl_1_8 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_440 wl_0_14 wl_1_14 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_462 wl_0_15 wl_1_15 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_473 wl_0_9 wl_1_9 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_451 wl_0_3 wl_1_3 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_484 wl_0_0 wl_1_0 bl_0_44 bl_1_44 br_0_44 br_1_44
+ sky130_fd_bd_sram__openram_dp_cell_484/a_38_n79# vdd_uq1278 gnd sky130_fd_bd_sram__openram_dp_cell_484/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_495 wl_0_2 wl_1_2 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5309 wl_0_102 wl_1_102 bl_0_29 bl_1_29 br_0_29
+ br_1_29 bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4619 wl_0_81 wl_1_81 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4608 wl_0_92 wl_1_92 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3907 wl_0_70 wl_1_70 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3918 wl_0_78 wl_1_78 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3929 wl_0_67 wl_1_67 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7212 wl_0_108 wl_1_108 bl_0_57 bl_1_57 br_0_57
+ br_1_57 bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7201 wl_0_104 wl_1_104 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7223 wl_0_100 wl_1_100 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7234 wl_0_109 wl_1_109 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7245 wl_0_107 wl_1_107 bl_0_59 bl_1_59 br_0_59
+ br_1_59 bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7267 wl_0_103 wl_1_103 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7256 wl_0_100 wl_1_100 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6511 wl_0_81 wl_1_81 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6522 wl_0_88 wl_1_88 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6500 wl_0_92 wl_1_92 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7278 wl_0_110 wl_1_110 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7289 wl_0_99 wl_1_99 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6544 wl_0_84 wl_1_84 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6555 wl_0_89 wl_1_89 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6533 wl_0_91 wl_1_91 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5810 wl_0_95 wl_1_95 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5832 wl_0_73 wl_1_73 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5821 wl_0_84 wl_1_84 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6577 wl_0_83 wl_1_83 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6588 wl_0_90 wl_1_90 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6566 wl_0_94 wl_1_94 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5843 wl_0_96 wl_1_96 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5887 wl_0_69 wl_1_69 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5876 wl_0_76 wl_1_76 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5865 wl_0_75 wl_1_75 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6599 wl_0_87 wl_1_87 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5854 wl_0_95 wl_1_95 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5898 wl_0_68 wl_1_68 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7790 wl_0_96 wl_1_96 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_292 wl_0_28 wl_1_28 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_281 wl_0_27 wl_1_27 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_270 wl_0_29 wl_1_29 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5106 wl_0_113 wl_1_113 bl_0_13 bl_1_13 br_0_13
+ br_1_13 bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5128 wl_0_125 wl_1_125 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5117 wl_0_119 wl_1_119 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5139 wl_0_114 wl_1_114 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4427 wl_0_67 wl_1_67 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4416 wl_0_70 wl_1_70 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4405 wl_0_72 wl_1_72 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4438 wl_0_74 wl_1_74 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3726 wl_0_32 wl_1_32 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3715 wl_0_49 wl_1_49 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3704 wl_0_60 wl_1_60 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4449 wl_0_77 wl_1_77 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3759 wl_0_31 wl_1_31 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3748 wl_0_42 wl_1_42 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3737 wl_0_53 wl_1_53 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7020 wl_0_118 wl_1_118 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7031 wl_0_117 wl_1_117 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7042 wl_0_124 wl_1_124 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7075 wl_0_123 wl_1_123 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7064 wl_0_120 wl_1_120 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7053 wl_0_113 wl_1_113 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6330 wl_0_78 wl_1_78 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7086 wl_0_118 wl_1_118 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7097 wl_0_107 wl_1_107 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6352 wl_0_65 wl_1_65 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6363 wl_0_72 wl_1_72 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6341 wl_0_76 wl_1_76 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5640 wl_0_121 wl_1_121 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5651 wl_0_110 wl_1_110 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5662 wl_0_99 wl_1_99 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6385 wl_0_65 wl_1_65 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6396 wl_0_66 wl_1_66 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6374 wl_0_72 wl_1_72 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5673 wl_0_112 wl_1_112 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4950 wl_0_107 wl_1_107 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5684 wl_0_95 wl_1_95 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5695 wl_0_96 wl_1_96 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4983 wl_0_118 wl_1_118 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4972 wl_0_115 wl_1_115 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4961 wl_0_114 wl_1_114 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4994 wl_0_126 wl_1_126 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1609 wl_0_60 wl_1_60 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4213 wl_0_82 wl_1_82 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4202 wl_0_93 wl_1_93 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3501 wl_0_49 wl_1_49 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4235 wl_0_81 wl_1_81 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4224 wl_0_88 wl_1_88 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4246 wl_0_92 wl_1_92 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3512 wl_0_52 wl_1_52 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3534 wl_0_60 wl_1_60 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3523 wl_0_59 wl_1_59 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4268 wl_0_70 wl_1_70 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4279 wl_0_79 wl_1_79 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4257 wl_0_81 wl_1_81 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2800 wl_0_20 wl_1_20 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2822 wl_0_13 wl_1_13 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2811 wl_0_8 wl_1_8 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2833 wl_0_2 wl_1_2 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3567 wl_0_51 wl_1_51 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3545 wl_0_53 wl_1_53 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3578 wl_0_58 wl_1_58 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3556 wl_0_62 wl_1_62 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2844 wl_0_16 wl_1_16 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2866 wl_0_39 wl_1_39 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2855 wl_0_41 wl_1_41 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3589 wl_0_59 wl_1_59 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2899 wl_0_35 wl_1_35 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2877 wl_0_41 wl_1_41 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2888 wl_0_46 wl_1_46 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6160 wl_0_88 wl_1_88 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6171 wl_0_94 wl_1_94 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5470 wl_0_117 wl_1_117 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6182 wl_0_85 wl_1_85 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6193 wl_0_92 wl_1_92 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5492 wl_0_124 wl_1_124 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5481 wl_0_116 wl_1_116 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4780 wl_0_105 wl_1_105 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4791 wl_0_104 wl_1_104 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2118 wl_0_9 wl_1_9 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2107 wl_0_6 wl_1_6 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2129 wl_0_1 wl_1_1 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1406 wl_0_39 wl_1_39 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1417 wl_0_43 wl_1_43 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1428 wl_0_33 wl_1_33 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1439 wl_0_41 wl_1_41 bl_0_50 bl_1_50 br_0_50 br_1_50
+ bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_814 wl_0_15 wl_1_15 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_803 wl_0_26 wl_1_26 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4021 wl_0_67 wl_1_67 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4010 wl_0_74 wl_1_74 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_836 wl_0_19 wl_1_19 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_847 wl_0_27 wl_1_27 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_825 wl_0_30 wl_1_30 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4043 wl_0_70 wl_1_70 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4054 wl_0_73 wl_1_73 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4032 wl_0_77 wl_1_77 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_858 wl_0_16 wl_1_16 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_869 wl_0_8 wl_1_8 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3320 wl_0_38 wl_1_38 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3342 wl_0_42 wl_1_42 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3331 wl_0_43 wl_1_43 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4065 wl_0_77 wl_1_77 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4076 wl_0_84 wl_1_84 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4087 wl_0_83 wl_1_83 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2630 wl_0_26 wl_1_26 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2641 wl_0_29 wl_1_29 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3386 wl_0_35 wl_1_35 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3364 wl_0_40 wl_1_40 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3353 wl_0_39 wl_1_39 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3375 wl_0_39 wl_1_39 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4098 wl_0_88 wl_1_88 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2674 wl_0_23 wl_1_23 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2663 wl_0_18 wl_1_18 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2652 wl_0_25 wl_1_25 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3397 wl_0_46 wl_1_46 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2685 wl_0_19 wl_1_19 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1973 wl_0_1 wl_1_1 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1962 wl_0_4 wl_1_4 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2696 wl_0_30 wl_1_30 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1940 wl_0_31 wl_1_31 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1951 wl_0_32 wl_1_32 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1995 wl_0_14 wl_1_14 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1984 wl_0_9 wl_1_9 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7619 wl_0_111 wl_1_111 bl_0_54 bl_1_54 br_0_54
+ br_1_54 bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7608 wl_0_106 wl_1_106 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6918 wl_0_120 wl_1_120 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6907 wl_0_118 wl_1_118 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6929 wl_0_113 wl_1_113 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1214 wl_0_51 wl_1_51 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1225 wl_0_61 wl_1_61 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1203 wl_0_62 wl_1_62 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1258 wl_0_36 wl_1_36 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1247 wl_0_45 wl_1_45 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1236 wl_0_47 wl_1_47 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1269 wl_0_59 wl_1_59 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_611 wl_0_14 wl_1_14 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_622 wl_0_7 wl_1_7 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_600 wl_0_8 wl_1_8 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_655 wl_0_19 wl_1_19 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_644 wl_0_12 wl_1_12 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_633 wl_0_4 wl_1_4 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_666 wl_0_23 wl_1_23 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_677 wl_0_17 wl_1_17 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_688 wl_0_23 wl_1_23 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_699 wl_0_26 wl_1_26 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3161 wl_0_54 wl_1_54 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3150 wl_0_60 wl_1_60 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3183 wl_0_49 wl_1_49 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3194 wl_0_51 wl_1_51 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3172 wl_0_60 wl_1_60 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2460 wl_0_7 wl_1_7 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2482 wl_0_2 wl_1_2 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2471 wl_0_4 wl_1_4 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2493 wl_0_1 wl_1_1 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1770 wl_0_31 wl_1_31 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1781 wl_0_52 wl_1_52 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1792 wl_0_41 wl_1_41 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8106 wl_0_23 wl_1_23 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8117 wl_0_12 wl_1_12 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7416 wl_0_123 wl_1_123 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7405 wl_0_117 wl_1_117 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8128 wl_0_1 wl_1_1 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8139 wl_0_63 wl_1_63 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7438 wl_0_116 wl_1_116 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7427 wl_0_114 wl_1_114 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7449 wl_0_113 wl_1_113 bl_0_63 bl_1_63 br_0_63
+ br_1_63 bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6704 wl_0_90 wl_1_90 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6737 wl_0_107 wl_1_107 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6726 wl_0_68 wl_1_68 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6715 wl_0_79 wl_1_79 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6759 wl_0_107 wl_1_107 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6748 wl_0_99 wl_1_99 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1000 wl_0_44 wl_1_44 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1011 wl_0_33 wl_1_33 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1033 wl_0_38 wl_1_38 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1022 wl_0_38 wl_1_38 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1044 wl_0_33 wl_1_33 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1055 wl_0_37 wl_1_37 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1066 wl_0_45 wl_1_45 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1077 wl_0_51 wl_1_51 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1088 wl_0_49 wl_1_49 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1099 wl_0_55 wl_1_55 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7961 wl_0_40 wl_1_40 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7950 wl_0_51 wl_1_51 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7983 wl_0_18 wl_1_18 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7994 wl_0_7 wl_1_7 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7972 wl_0_29 wl_1_29 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_441 wl_0_13 wl_1_13 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_430 wl_0_24 wl_1_24 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_463 wl_0_16 wl_1_16 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_474 wl_0_8 wl_1_8 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_452 wl_0_2 wl_1_2 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_485 wl_0_9 wl_1_9 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_496 wl_0_1 wl_1_1 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2290 wl_0_29 wl_1_29 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4609 wl_0_91 wl_1_91 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3908 wl_0_69 wl_1_69 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3919 wl_0_77 wl_1_77 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7213 wl_0_110 wl_1_110 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7202 wl_0_103 wl_1_103 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7224 wl_0_99 wl_1_99 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7246 wl_0_110 wl_1_110 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7235 wl_0_108 wl_1_108 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7257 wl_0_99 wl_1_99 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6512 wl_0_88 wl_1_88 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6501 wl_0_91 wl_1_91 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7279 wl_0_109 wl_1_109 bl_0_51 bl_1_51 br_0_51
+ br_1_51 bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5800 wl_0_105 wl_1_105 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7268 wl_0_102 wl_1_102 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6545 wl_0_83 wl_1_83 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6556 wl_0_88 wl_1_88 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6523 wl_0_87 wl_1_87 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5811 wl_0_94 wl_1_94 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6534 wl_0_94 wl_1_94 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5833 wl_0_72 wl_1_72 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6578 wl_0_82 wl_1_82 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5822 wl_0_83 wl_1_83 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6589 wl_0_89 wl_1_89 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6567 wl_0_93 wl_1_93 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5844 wl_0_95 wl_1_95 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5866 wl_0_74 wl_1_74 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5877 wl_0_75 wl_1_75 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5855 wl_0_96 wl_1_96 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5899 wl_0_67 wl_1_67 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5888 wl_0_68 wl_1_68 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7780 wl_0_70 wl_1_70 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7791 wl_0_95 wl_1_95 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_271 wl_0_28 wl_1_28 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_260 wl_0_29 wl_1_29 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_282 wl_0_30 wl_1_30 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_293 wl_0_27 wl_1_27 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5129 wl_0_124 wl_1_124 bl_0_11 bl_1_11 br_0_11
+ br_1_11 bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5107 wl_0_120 wl_1_120 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5118 wl_0_118 wl_1_118 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4428 wl_0_66 wl_1_66 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4417 wl_0_69 wl_1_69 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4406 wl_0_71 wl_1_71 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3727 wl_0_31 wl_1_31 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3716 wl_0_48 wl_1_48 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3705 wl_0_59 wl_1_59 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4439 wl_0_73 wl_1_73 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3749 wl_0_41 wl_1_41 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3738 wl_0_52 wl_1_52 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7021 wl_0_127 wl_1_127 bl_0_43 bl_1_43 br_0_43
+ br_1_43 sky130_fd_bd_sram__openram_dp_cell_7021/a_38_n79# vdd_uq1342 gnd sky130_fd_bd_sram__openram_dp_cell_7021/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7010 wl_0_120 wl_1_120 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7032 wl_0_116 wl_1_116 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7043 wl_0_123 wl_1_123 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7065 wl_0_119 wl_1_119 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7054 wl_0_114 wl_1_114 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6320 wl_0_72 wl_1_72 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7076 wl_0_127 wl_1_127 bl_0_45 bl_1_45 br_0_45
+ br_1_45 sky130_fd_bd_sram__openram_dp_cell_7076/a_38_n79# vdd_uq1214 gnd sky130_fd_bd_sram__openram_dp_cell_7076/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7087 wl_0_117 wl_1_117 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7098 wl_0_106 wl_1_106 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6353 wl_0_69 wl_1_69 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6364 wl_0_71 wl_1_71 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6342 wl_0_75 wl_1_75 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6331 wl_0_77 wl_1_77 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5641 wl_0_120 wl_1_120 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5652 wl_0_109 wl_1_109 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5630 wl_0_100 wl_1_100 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6375 wl_0_71 wl_1_71 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6386 wl_0_75 wl_1_75 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6397 wl_0_78 wl_1_78 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5674 wl_0_111 wl_1_111 bl_0_18 bl_1_18 br_0_18
+ br_1_18 bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4951 wl_0_106 wl_1_106 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4940 wl_0_103 wl_1_103 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5663 wl_0_98 wl_1_98 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5685 wl_0_96 wl_1_96 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4984 wl_0_117 wl_1_117 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4973 wl_0_117 wl_1_117 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4962 wl_0_113 wl_1_113 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5696 wl_0_95 wl_1_95 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4995 wl_0_125 wl_1_125 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4203 wl_0_92 wl_1_92 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4214 wl_0_81 wl_1_81 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4225 wl_0_87 wl_1_87 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4236 wl_0_94 wl_1_94 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3513 wl_0_51 wl_1_51 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3524 wl_0_58 wl_1_58 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3535 wl_0_59 wl_1_59 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3502 wl_0_62 wl_1_62 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4269 wl_0_69 wl_1_69 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4258 wl_0_80 wl_1_80 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4247 wl_0_91 wl_1_91 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2801 wl_0_19 wl_1_19 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2823 wl_0_12 wl_1_12 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2812 wl_0_7 wl_1_7 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3568 wl_0_50 wl_1_50 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3546 wl_0_52 wl_1_52 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3557 wl_0_61 wl_1_61 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2845 wl_0_15 wl_1_15 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2834 wl_0_1 wl_1_1 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2856 wl_0_46 wl_1_46 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3579 wl_0_57 wl_1_57 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2867 wl_0_38 wl_1_38 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2878 wl_0_40 wl_1_40 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2889 wl_0_45 wl_1_45 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6150 wl_0_83 wl_1_83 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6161 wl_0_87 wl_1_87 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6172 wl_0_93 wl_1_93 bl_0_59 bl_1_59 br_0_59 br_1_59
+ bl_1_59 vdd_uq318 gnd br_1_59 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5460 wl_0_118 wl_1_118 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6183 wl_0_84 wl_1_84 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6194 wl_0_91 wl_1_91 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5471 wl_0_126 wl_1_126 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5493 wl_0_123 wl_1_123 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5482 wl_0_115 wl_1_115 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4792 wl_0_103 wl_1_103 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4781 wl_0_104 wl_1_104 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4770 wl_0_80 wl_1_80 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2119 wl_0_8 wl_1_8 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2108 wl_0_0 wl_1_0 bl_0_21 bl_1_21 br_0_21 br_1_21
+ sky130_fd_bd_sram__openram_dp_cell_2108/a_38_n79# vdd_uq2750 gnd sky130_fd_bd_sram__openram_dp_cell_2108/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1407 wl_0_46 wl_1_46 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1418 wl_0_42 wl_1_42 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1429 wl_0_44 wl_1_44 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_815 wl_0_16 wl_1_16 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_804 wl_0_30 wl_1_30 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4000 wl_0_68 wl_1_68 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4011 wl_0_73 wl_1_73 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_837 wl_0_18 wl_1_18 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_848 wl_0_26 wl_1_26 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_826 wl_0_29 wl_1_29 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3310 wl_0_36 wl_1_36 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4022 wl_0_66 wl_1_66 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4044 wl_0_69 wl_1_69 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4055 wl_0_72 wl_1_72 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4033 wl_0_78 wl_1_78 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_859 wl_0_15 wl_1_15 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3321 wl_0_37 wl_1_37 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3343 wl_0_41 wl_1_41 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3332 wl_0_42 wl_1_42 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4066 wl_0_76 wl_1_76 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4088 wl_0_82 wl_1_82 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4077 wl_0_83 wl_1_83 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2620 wl_0_23 wl_1_23 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2631 wl_0_25 wl_1_25 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3354 wl_0_38 wl_1_38 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3376 wl_0_38 wl_1_38 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3365 wl_0_39 wl_1_39 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4099 wl_0_87 wl_1_87 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2653 wl_0_24 wl_1_24 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2675 wl_0_22 wl_1_22 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2664 wl_0_17 wl_1_17 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2642 wl_0_28 wl_1_28 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1930 wl_0_32 wl_1_32 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3387 wl_0_34 wl_1_34 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3398 wl_0_45 wl_1_45 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2686 wl_0_18 wl_1_18 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1963 wl_0_3 wl_1_3 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2697 wl_0_29 wl_1_29 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1941 wl_0_32 wl_1_32 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1952 wl_0_31 wl_1_31 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1996 wl_0_13 wl_1_13 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1985 wl_0_8 wl_1_8 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1974 wl_0_0 wl_1_0 bl_0_28 bl_1_28 br_0_28 br_1_28
+ sky130_fd_bd_sram__openram_dp_cell_1974/a_38_n79# vdd_uq2302 gnd sky130_fd_bd_sram__openram_dp_cell_1974/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5290 wl_0_108 wl_1_108 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7609 wl_0_105 wl_1_105 bl_0_55 bl_1_55 br_0_55
+ br_1_55 bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6919 wl_0_119 wl_1_119 bl_0_36 bl_1_36 br_0_36
+ br_1_36 bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6908 wl_0_116 wl_1_116 bl_0_34 bl_1_34 br_0_34
+ br_1_34 bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1215 wl_0_50 wl_1_50 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1226 wl_0_60 wl_1_60 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1204 wl_0_61 wl_1_61 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1259 wl_0_35 wl_1_35 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1248 wl_0_44 wl_1_44 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1237 wl_0_55 wl_1_55 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_612 wl_0_13 wl_1_13 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_601 wl_0_7 wl_1_7 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_623 wl_0_6 wl_1_6 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_634 wl_0_3 wl_1_3 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_645 wl_0_30 wl_1_30 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_656 wl_0_30 wl_1_30 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_667 wl_0_22 wl_1_22 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_689 wl_0_22 wl_1_22 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_678 wl_0_20 wl_1_20 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3140 wl_0_55 wl_1_55 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3151 wl_0_59 wl_1_59 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2450 wl_0_2 wl_1_2 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3162 wl_0_53 wl_1_53 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3184 wl_0_56 wl_1_56 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3173 wl_0_59 wl_1_59 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2461 wl_0_6 wl_1_6 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2483 wl_0_6 wl_1_6 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2472 wl_0_3 wl_1_3 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3195 wl_0_50 wl_1_50 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2494 wl_0_0 wl_1_0 bl_0_1 bl_1_1 br_0_1 br_1_1
+ sky130_fd_bd_sram__openram_dp_cell_2494/a_38_n79# vdd_uq4030 gnd sky130_fd_bd_sram__openram_dp_cell_2494/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1760 wl_0_39 wl_1_39 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1771 wl_0_62 wl_1_62 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1793 wl_0_40 wl_1_40 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1782 wl_0_51 wl_1_51 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8107 wl_0_22 wl_1_22 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8118 wl_0_11 wl_1_11 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7406 wl_0_116 wl_1_116 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8129 wl_0_0 wl_1_0 bl_0_31 bl_1_31 br_0_31 br_1_31
+ sky130_fd_bd_sram__openram_dp_cell_8129/a_38_n79# vdd_uq2110 gnd sky130_fd_bd_sram__openram_dp_cell_8129/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7417 wl_0_122 wl_1_122 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7439 wl_0_115 wl_1_115 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7428 wl_0_113 wl_1_113 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6705 wl_0_89 wl_1_89 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6738 wl_0_106 wl_1_106 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6716 wl_0_78 wl_1_78 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6727 wl_0_80 wl_1_80 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6749 wl_0_98 wl_1_98 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1012 wl_0_36 wl_1_36 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1034 wl_0_37 wl_1_37 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1023 wl_0_37 wl_1_37 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1001 wl_0_43 wl_1_43 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1056 wl_0_36 wl_1_36 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1045 wl_0_45 wl_1_45 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1067 wl_0_61 wl_1_61 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1089 wl_0_49 wl_1_49 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1078 wl_0_50 wl_1_50 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7962 wl_0_39 wl_1_39 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7951 wl_0_50 wl_1_50 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7940 wl_0_61 wl_1_61 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7984 wl_0_17 wl_1_17 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7995 wl_0_6 wl_1_6 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7973 wl_0_28 wl_1_28 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_420 wl_0_16 wl_1_16 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_431 wl_0_23 wl_1_23 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_464 wl_0_15 wl_1_15 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_442 wl_0_12 wl_1_12 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_453 wl_0_1 wl_1_1 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_486 wl_0_8 wl_1_8 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_475 wl_0_7 wl_1_7 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_497 wl_0_0 wl_1_0 bl_0_45 bl_1_45 br_0_45 br_1_45
+ sky130_fd_bd_sram__openram_dp_cell_497/a_38_n79# vdd_uq1214 gnd sky130_fd_bd_sram__openram_dp_cell_497/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2280 wl_0_18 wl_1_18 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2291 wl_0_28 wl_1_28 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1590 wl_0_59 wl_1_59 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3909 wl_0_68 wl_1_68 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7214 wl_0_109 wl_1_109 bl_0_62 bl_1_62 br_0_62
+ br_1_62 bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7203 wl_0_102 wl_1_102 bl_0_60 bl_1_60 br_0_60
+ br_1_60 bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7247 wl_0_109 wl_1_109 bl_0_61 bl_1_61 br_0_61
+ br_1_61 bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7236 wl_0_107 wl_1_107 bl_0_58 bl_1_58 br_0_58
+ br_1_58 bl_1_58 vdd_uq382 gnd br_1_58 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7225 wl_0_98 wl_1_98 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7258 wl_0_98 wl_1_98 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6513 wl_0_87 wl_1_87 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6502 wl_0_88 wl_1_88 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5801 wl_0_104 wl_1_104 bl_0_15 bl_1_15 br_0_15
+ br_1_15 bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7269 wl_0_101 wl_1_101 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6546 wl_0_82 wl_1_82 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6524 wl_0_86 wl_1_86 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6535 wl_0_93 wl_1_93 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5834 wl_0_71 wl_1_71 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6579 wl_0_81 wl_1_81 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5823 wl_0_82 wl_1_82 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6557 wl_0_87 wl_1_87 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6568 wl_0_92 wl_1_92 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5812 wl_0_93 wl_1_93 bl_0_15 bl_1_15 br_0_15 br_1_15
+ bl_1_15 vdd_uq3134 gnd br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5867 wl_0_73 wl_1_73 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5878 wl_0_78 wl_1_78 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5856 wl_0_95 wl_1_95 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5845 wl_0_96 wl_1_96 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5889 wl_0_67 wl_1_67 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7770 wl_0_80 wl_1_80 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7792 wl_0_96 wl_1_96 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7781 wl_0_69 wl_1_69 bl_0_47 bl_1_47 br_0_47 br_1_47
+ bl_1_47 vdd_uq1086 gnd br_1_47 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_250 wl_0_17 wl_1_17 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_261 wl_0_28 wl_1_28 bl_0_49 bl_1_49 br_0_49 br_1_49
+ bl_1_49 vdd_uq958 gnd br_1_49 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_272 wl_0_27 wl_1_27 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_283 wl_0_29 wl_1_29 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_294 wl_0_26 wl_1_26 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5108 wl_0_119 wl_1_119 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5119 wl_0_117 wl_1_117 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4429 wl_0_65 wl_1_65 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4418 wl_0_68 wl_1_68 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4407 wl_0_78 wl_1_78 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3717 wl_0_47 wl_1_47 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3706 wl_0_58 wl_1_58 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3739 wl_0_51 wl_1_51 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3728 wl_0_62 wl_1_62 bl_0_16 bl_1_16 br_0_16 br_1_16
+ bl_1_16 vdd_uq3070 gnd br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7022 wl_0_126 wl_1_126 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7011 wl_0_119 wl_1_119 bl_0_44 bl_1_44 br_0_44
+ br_1_44 bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7000 wl_0_113 wl_1_113 bl_0_45 bl_1_45 br_0_45
+ br_1_45 bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7044 wl_0_122 wl_1_122 bl_0_42 bl_1_42 br_0_42
+ br_1_42 bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7066 wl_0_118 wl_1_118 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7033 wl_0_115 wl_1_115 bl_0_43 bl_1_43 br_0_43
+ br_1_43 bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7055 wl_0_113 wl_1_113 bl_0_41 bl_1_41 br_0_41
+ br_1_41 bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6321 wl_0_71 wl_1_71 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6310 wl_0_71 wl_1_71 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7077 wl_0_127 wl_1_127 bl_0_40 bl_1_40 br_0_40
+ br_1_40 sky130_fd_bd_sram__openram_dp_cell_7077/a_38_n79# vdd_uq1534 gnd sky130_fd_bd_sram__openram_dp_cell_7077/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7088 wl_0_116 wl_1_116 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7099 wl_0_105 wl_1_105 bl_0_40 bl_1_40 br_0_40
+ br_1_40 bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6354 wl_0_68 wl_1_68 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6343 wl_0_74 wl_1_74 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6332 wl_0_76 wl_1_76 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5642 wl_0_119 wl_1_119 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5620 wl_0_110 wl_1_110 bl_0_24 bl_1_24 br_0_24
+ br_1_24 bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5653 wl_0_108 wl_1_108 bl_0_23 bl_1_23 br_0_23
+ br_1_23 bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5631 wl_0_99 wl_1_99 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6365 wl_0_70 wl_1_70 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6376 wl_0_70 wl_1_70 bl_0_43 bl_1_43 br_0_43 br_1_43
+ bl_1_43 vdd_uq1342 gnd br_1_43 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6387 wl_0_74 wl_1_74 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6398 wl_0_76 wl_1_76 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4941 wl_0_102 wl_1_102 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4930 wl_0_101 wl_1_101 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5664 wl_0_97 wl_1_97 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5675 wl_0_96 wl_1_96 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5686 wl_0_95 wl_1_95 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4974 wl_0_118 wl_1_118 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4963 wl_0_117 wl_1_117 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4952 wl_0_105 wl_1_105 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5697 wl_0_96 wl_1_96 bl_0_24 bl_1_24 br_0_24 br_1_24
+ bl_1_24 vdd_uq2558 gnd br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4996 wl_0_124 wl_1_124 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4985 wl_0_116 wl_1_116 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4226 wl_0_86 wl_1_86 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4215 wl_0_87 wl_1_87 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4204 wl_0_91 wl_1_91 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4237 wl_0_93 wl_1_93 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3514 wl_0_50 wl_1_50 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3525 wl_0_57 wl_1_57 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3503 wl_0_61 wl_1_61 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4259 wl_0_79 wl_1_79 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4248 wl_0_90 wl_1_90 bl_0_23 bl_1_23 br_0_23 br_1_23
+ bl_1_23 vdd_uq2622 gnd br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2802 wl_0_18 wl_1_18 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2824 wl_0_11 wl_1_11 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2813 wl_0_6 wl_1_6 bl_0_7 bl_1_7 br_0_7 br_1_7
+ bl_1_7 vdd_uq3646 gnd br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3569 wl_0_49 wl_1_49 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3547 wl_0_51 wl_1_51 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3558 wl_0_60 wl_1_60 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3536 wl_0_62 wl_1_62 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2846 wl_0_16 wl_1_16 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2835 wl_0_0 wl_1_0 bl_0_8 bl_1_8 br_0_8 br_1_8
+ sky130_fd_bd_sram__openram_dp_cell_2835/a_38_n79# vdd_uq3582 gnd sky130_fd_bd_sram__openram_dp_cell_2835/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2857 wl_0_45 wl_1_45 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2868 wl_0_37 wl_1_37 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2879 wl_0_39 wl_1_39 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6140 wl_0_81 wl_1_81 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6151 wl_0_82 wl_1_82 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6162 wl_0_86 wl_1_86 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5450 wl_0_120 wl_1_120 bl_0_17 bl_1_17 br_0_17
+ br_1_17 bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5461 wl_0_117 wl_1_117 bl_0_21 bl_1_21 br_0_21
+ br_1_21 bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6184 wl_0_83 wl_1_83 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6195 wl_0_90 wl_1_90 bl_0_61 bl_1_61 br_0_61 br_1_61
+ bl_1_61 vdd_uq190 gnd br_1_61 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6173 wl_0_94 wl_1_94 bl_0_62 bl_1_62 br_0_62 br_1_62
+ bl_1_62 vdd_uq99 gnd br_1_62 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5472 wl_0_125 wl_1_125 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5494 wl_0_122 wl_1_122 bl_0_19 bl_1_19 br_0_19
+ br_1_19 bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5483 wl_0_114 wl_1_114 bl_0_20 bl_1_20 br_0_20
+ br_1_20 bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4782 wl_0_103 wl_1_103 bl_0_12 bl_1_12 br_0_12
+ br_1_12 bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4793 wl_0_102 wl_1_102 bl_0_14 bl_1_14 br_0_14
+ br_1_14 bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4760 wl_0_72 wl_1_72 bl_0_8 bl_1_8 br_0_8 br_1_8
+ bl_1_8 vdd_uq3582 gnd br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4771 wl_0_79 wl_1_79 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2109 wl_0_8 wl_1_8 bl_0_19 bl_1_19 br_0_19 br_1_19
+ bl_1_19 vdd_uq2878 gnd br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1408 wl_0_45 wl_1_45 bl_0_60 bl_1_60 br_0_60 br_1_60
+ bl_1_60 vdd_uq254 gnd br_1_60 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1419 wl_0_41 wl_1_41 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_805 wl_0_29 wl_1_29 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4001 wl_0_67 wl_1_67 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4012 wl_0_72 wl_1_72 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_838 wl_0_17 wl_1_17 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_816 wl_0_15 wl_1_15 bl_0_46 bl_1_46 br_0_46 br_1_46
+ bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_827 wl_0_28 wl_1_28 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3300 wl_0_48 wl_1_48 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4023 wl_0_65 wl_1_65 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4045 wl_0_68 wl_1_68 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4034 wl_0_77 wl_1_77 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_849 wl_0_25 wl_1_25 bl_0_40 bl_1_40 br_0_40 br_1_40
+ bl_1_40 vdd_uq1534 gnd br_1_40 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3311 wl_0_35 wl_1_35 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3322 wl_0_36 wl_1_36 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3333 wl_0_41 wl_1_41 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4056 wl_0_71 wl_1_71 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4067 wl_0_75 wl_1_75 bl_0_17 bl_1_17 br_0_17 br_1_17
+ bl_1_17 vdd_uq3006 gnd br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4078 wl_0_82 wl_1_82 bl_0_20 bl_1_20 br_0_20 br_1_20
+ bl_1_20 vdd_uq2814 gnd br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2632 wl_0_24 wl_1_24 bl_0_2 bl_1_2 br_0_2 br_1_2
+ bl_1_2 vdd_uq3966 gnd br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2621 wl_0_22 wl_1_22 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2610 wl_0_28 wl_1_28 bl_0_1 bl_1_1 br_0_1 br_1_1
+ bl_1_1 vdd_uq4030 gnd br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3355 wl_0_37 wl_1_37 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3377 wl_0_37 wl_1_37 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3366 wl_0_38 wl_1_38 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3344 wl_0_46 wl_1_46 bl_0_27 bl_1_27 br_0_27 br_1_27
+ bl_1_27 vdd_uq2366 gnd br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4089 wl_0_81 wl_1_81 bl_0_22 bl_1_22 br_0_22 br_1_22
+ bl_1_22 vdd_uq2686 gnd br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2654 wl_0_23 wl_1_23 bl_0_4 bl_1_4 br_0_4 br_1_4
+ bl_1_4 vdd_uq3838 gnd br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2665 wl_0_20 wl_1_20 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2643 wl_0_27 wl_1_27 bl_0_6 bl_1_6 br_0_6 br_1_6
+ bl_1_6 vdd_uq3710 gnd br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1920 wl_0_31 wl_1_31 bl_0_57 bl_1_57 br_0_57 br_1_57
+ bl_1_57 vdd_uq446 gnd br_1_57 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3388 wl_0_33 wl_1_33 bl_0_18 bl_1_18 br_0_18 br_1_18
+ bl_1_18 vdd_uq2942 gnd br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3399 wl_0_44 wl_1_44 bl_0_21 bl_1_21 br_0_21 br_1_21
+ bl_1_21 vdd_uq2750 gnd br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2676 wl_0_21 wl_1_21 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1953 wl_0_13 wl_1_13 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1964 wl_0_2 wl_1_2 bl_0_29 bl_1_29 br_0_29 br_1_29
+ bl_1_29 vdd_uq2238 gnd br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2698 wl_0_28 wl_1_28 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2687 wl_0_30 wl_1_30 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1942 wl_0_31 wl_1_31 bl_0_42 bl_1_42 br_0_42 br_1_42
+ bl_1_42 vdd_uq1406 gnd br_1_42 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1931 wl_0_31 wl_1_31 bl_0_54 bl_1_54 br_0_54 br_1_54
+ bl_1_54 vdd_uq638 gnd br_1_54 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1975 wl_0_12 wl_1_12 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1997 wl_0_12 wl_1_12 bl_0_25 bl_1_25 br_0_25 br_1_25
+ bl_1_25 vdd_uq2494 gnd br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1986 wl_0_7 wl_1_7 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5291 wl_0_107 wl_1_107 bl_0_26 bl_1_26 br_0_26
+ br_1_26 bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5280 wl_0_98 wl_1_98 bl_0_30 bl_1_30 br_0_30 br_1_30
+ bl_1_30 vdd_uq2174 gnd br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4590 wl_0_94 wl_1_94 bl_0_3 bl_1_3 br_0_3 br_1_3
+ bl_1_3 vdd_uq3902 gnd br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6909 wl_0_118 wl_1_118 bl_0_33 bl_1_33 br_0_33
+ br_1_33 bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1216 wl_0_49 wl_1_49 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1205 wl_0_60 wl_1_60 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1249 wl_0_43 wl_1_43 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1238 wl_0_54 wl_1_54 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1227 wl_0_59 wl_1_59 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_613 wl_0_12 wl_1_12 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_602 wl_0_6 wl_1_6 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_635 wl_0_2 wl_1_2 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_624 wl_0_5 wl_1_5 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_646 wl_0_29 wl_1_29 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_657 wl_0_29 wl_1_29 bl_0_38 bl_1_38 br_0_38 br_1_38
+ bl_1_38 vdd_uq1662 gnd br_1_38 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_679 wl_0_21 wl_1_21 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_668 wl_0_30 wl_1_30 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3130 wl_0_54 wl_1_54 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3141 wl_0_54 wl_1_54 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3152 wl_0_58 wl_1_58 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2440 wl_0_2 wl_1_2 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3163 wl_0_52 wl_1_52 bl_0_12 bl_1_12 br_0_12 br_1_12
+ bl_1_12 vdd_uq3326 gnd br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3185 wl_0_55 wl_1_55 bl_0_13 bl_1_13 br_0_13 br_1_13
+ bl_1_13 vdd_uq3262 gnd br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3174 wl_0_58 wl_1_58 bl_0_14 bl_1_14 br_0_14 br_1_14
+ bl_1_14 vdd_uq3198 gnd br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2451 wl_0_1 wl_1_1 bl_0_11 bl_1_11 br_0_11 br_1_11
+ bl_1_11 vdd_uq3390 gnd br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2473 wl_0_2 wl_1_2 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2462 wl_0_5 wl_1_5 bl_0_10 bl_1_10 br_0_10 br_1_10
+ bl_1_10 vdd_uq3454 gnd br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3196 wl_0_62 wl_1_62 bl_0_9 bl_1_9 br_0_9 br_1_9
+ bl_1_9 vdd_uq3518 gnd br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2495 wl_0_1 wl_1_1 bl_0_0 bl_1_0 br_0_0 br_1_0
+ bl_1_0 vdd_uq4094 gnd br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2484 wl_0_5 wl_1_5 bl_0_5 bl_1_5 br_0_5 br_1_5
+ bl_1_5 vdd_uq3774 gnd br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1761 wl_0_38 wl_1_38 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1750 wl_0_49 wl_1_49 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1772 wl_0_61 wl_1_61 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1794 wl_0_39 wl_1_39 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1783 wl_0_50 wl_1_50 bl_0_48 bl_1_48 br_0_48 br_1_48
+ bl_1_48 vdd_uq999 gnd br_1_48 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8108 wl_0_21 wl_1_21 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7407 wl_0_115 wl_1_115 bl_0_53 bl_1_53 br_0_53
+ br_1_53 bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8119 wl_0_10 wl_1_10 bl_0_31 bl_1_31 br_0_31 br_1_31
+ bl_1_31 vdd_uq2110 gnd br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7418 wl_0_121 wl_1_121 bl_0_52 bl_1_52 br_0_52
+ br_1_52 bl_1_52 vdd_uq766 gnd br_1_52 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7429 wl_0_113 wl_1_113 bl_0_50 bl_1_50 br_0_50
+ br_1_50 bl_1_50 vdd_uq894 gnd br_1_50 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6717 wl_0_77 wl_1_77 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6728 wl_0_79 wl_1_79 bl_0_44 bl_1_44 br_0_44 br_1_44
+ bl_1_44 vdd_uq1278 gnd br_1_44 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6706 wl_0_88 wl_1_88 bl_0_39 bl_1_39 br_0_39 br_1_39
+ bl_1_39 vdd_uq1598 gnd br_1_39 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6739 wl_0_105 wl_1_105 bl_0_46 bl_1_46 br_0_46
+ br_1_46 bl_1_46 vdd_uq1150 gnd br_1_46 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1013 wl_0_35 wl_1_35 bl_0_36 bl_1_36 br_0_36 br_1_36
+ bl_1_36 vdd_uq1790 gnd br_1_36 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1002 wl_0_42 wl_1_42 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1024 wl_0_46 wl_1_46 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1035 wl_0_36 wl_1_36 bl_0_34 bl_1_34 br_0_34 br_1_34
+ bl_1_34 vdd_uq1918 gnd br_1_34 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1057 wl_0_43 wl_1_43 bl_0_35 bl_1_35 br_0_35 br_1_35
+ bl_1_35 vdd_uq1854 gnd br_1_35 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1046 wl_0_44 wl_1_44 bl_0_37 bl_1_37 br_0_37 br_1_37
+ bl_1_37 vdd_uq1726 gnd br_1_37 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1068 wl_0_60 wl_1_60 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1079 wl_0_49 wl_1_49 bl_0_33 bl_1_33 br_0_33 br_1_33
+ bl_1_33 vdd_uq1982 gnd br_1_33 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7952 wl_0_49 wl_1_49 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7941 wl_0_60 wl_1_60 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7930 wl_0_71 wl_1_71 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7985 wl_0_16 wl_1_16 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7996 wl_0_5 wl_1_5 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7974 wl_0_27 wl_1_27 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7963 wl_0_38 wl_1_38 bl_0_32 bl_1_32 br_0_32 br_1_32
+ bl_1_32 vdd_uq2046 gnd br_1_32 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_432 wl_0_22 wl_1_22 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_421 wl_0_15 wl_1_15 bl_0_53 bl_1_53 br_0_53 br_1_53
+ bl_1_53 vdd_uq702 gnd br_1_53 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_410 wl_0_1 wl_1_1 bl_0_55 bl_1_55 br_0_55 br_1_55
+ bl_1_55 vdd_uq574 gnd br_1_55 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_443 wl_0_11 wl_1_11 bl_0_56 bl_1_56 br_0_56 br_1_56
+ bl_1_56 vdd_uq510 gnd br_1_56 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_465 wl_0_6 wl_1_6 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_454 wl_0_0 wl_1_0 bl_0_56 bl_1_56 br_0_56 br_1_56
+ sky130_fd_bd_sram__openram_dp_cell_454/a_38_n79# vdd_uq510 gnd sky130_fd_bd_sram__openram_dp_cell_454/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_498 wl_0_10 wl_1_10 bl_0_41 bl_1_41 br_0_41 br_1_41
+ bl_1_41 vdd_uq1470 gnd br_1_41 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_487 wl_0_7 wl_1_7 bl_0_45 bl_1_45 br_0_45 br_1_45
+ bl_1_45 vdd_uq1214 gnd br_1_45 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_476 wl_0_0 wl_1_0 bl_0_41 bl_1_41 br_0_41 br_1_41
+ sky130_fd_bd_sram__openram_dp_cell_476/a_38_n79# vdd_uq1470 gnd sky130_fd_bd_sram__openram_dp_cell_476/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2281 wl_0_17 wl_1_17 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2292 wl_0_27 wl_1_27 bl_0_26 bl_1_26 br_0_26 br_1_26
+ bl_1_26 vdd_uq2430 gnd br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2270 wl_0_28 wl_1_28 bl_0_28 bl_1_28 br_0_28 br_1_28
+ bl_1_28 vdd_uq2302 gnd br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1580 wl_0_54 wl_1_54 bl_0_51 bl_1_51 br_0_51 br_1_51
+ bl_1_51 vdd_uq830 gnd br_1_51 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1591 wl_0_58 wl_1_58 bl_0_63 bl_1_63 br_0_63 br_1_63
+ bl_1_63 vdd gnd br_1_63 sky130_fd_bd_sram__openram_dp_cell
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_replica_bitcell_array wl_1_113 wl_0_114
+ wl_1_114 wl_0_115 wl_0_116 wl_1_116 wl_0_117 wl_0_118 wl_0_119 wl_1_122 wl_1_123
+ wl_0_125 wl_1_125 wl_0_126 wl_0_127 rbl_wl_1_1 wl_1_96 wl_1_98 wl_1_101 wl_0_103
+ wl_0_104 wl_0_105 wl_0_106 wl_0_107 wl_1_107 wl_0_108 wl_0_109 wl_1_110 wl_1_83
+ wl_1_84 wl_1_85 wl_1_86 wl_1_72 wl_1_87 wl_1_89 wl_1_64 wl_1_91 wl_1_92 wl_1_73
+ wl_1_74 wl_1_65 wl_1_93 wl_1_94 wl_1_95 wl_1_75 wl_1_69 wl_1_77 wl_1_66 wl_1_78
+ wl_1_80 wl_1_70 wl_1_81 wl_1_67 wl_1_71 wl_1_82 wl_1_31 wl_1_32 wl_1_34 wl_1_36
+ wl_0_37 wl_1_37 wl_0_38 wl_1_38 wl_0_39 wl_1_40 wl_1_41 wl_1_42 wl_1_43 wl_1_44
+ wl_1_45 wl_1_46 wl_1_47 wl_0_48 wl_0_49 wl_1_49 wl_1_50 wl_1_51 wl_1_52 wl_1_53
+ wl_1_55 wl_1_56 wl_1_58 wl_0_59 wl_1_59 wl_1_60 wl_1_61 wl_1_62 wl_1_63 wl_0_1 wl_1_30
+ wl_1_1 wl_0_2 wl_1_13 wl_0_26 wl_1_2 wl_1_14 wl_0_3 wl_1_3 wl_0_15 wl_1_26 wl_0_4
+ wl_0_16 wl_1_16 wl_0_17 wl_1_17 wl_0_28 wl_0_18 wl_1_28 wl_0_29 wl_0_19 wl_1_19
+ rbl_wl_0_0 wl_0_27 wl_1_8 wl_1_20 wl_0_9 wl_1_0 wl_1_10 wl_1_22 wl_1_11 wl_1_23
+ wl_1_25 br_0_15 bl_1_16 br_0_16 br_1_16 bl_1_17 br_0_17 br_1_17 bl_1_18 br_0_18
+ br_1_18 bl_1_19 br_0_19 br_1_19 br_0_20 br_1_20 br_0_21 br_1_21 br_0_22 br_1_22
+ bl_1_23 br_0_23 br_1_23 bl_1_24 br_0_24 br_1_24 bl_1_25 br_0_25 br_1_25 bl_1_26
+ br_0_26 br_1_26 bl_1_27 br_0_27 br_1_27 bl_1_28 br_0_28 br_1_28 bl_1_29 br_0_29
+ br_1_29 br_0_30 br_1_30 br_0_31 br_1_31 br_0_12 br_1_12 bl_1_13 br_0_13 br_1_13
+ bl_1_14 br_0_14 br_1_14 rbl_br_0_0 bl_1_15 rbl_br_1_0 br_1_15 bl_0_0 br_0_0 br_1_0
+ bl_0_1 br_0_1 br_1_1 bl_0_2 br_0_2 br_1_2 bl_0_3 br_0_3 br_1_3 bl_0_4 bl_1_4 br_0_4
+ bl_0_5 br_0_10 br_1_10 br_0_11 br_1_11 bl_1_12 rbl_bl_0_0 rbl_bl_1_0 bl_1_48 br_1_48
+ bl_1_49 br_0_49 br_1_49 br_0_50 br_0_51 br_1_51 br_0_52 br_1_52 br_0_53 br_1_53
+ br_0_54 br_1_54 br_0_55 br_1_55 bl_1_56 br_0_56 br_1_56 bl_1_57 br_0_57 br_1_57
+ bl_1_58 br_0_58 br_1_58 bl_1_59 br_0_59 br_1_59 br_0_60 br_0_61 br_0_62 br_1_62
+ br_0_63 br_1_63 rbl_bl_0_1 rbl_br_0_1 bl_1_34 br_0_34 br_1_34 bl_1_35 br_0_35 br_1_35
+ br_0_46 br_0_48 bl_1_36 br_0_36 br_1_36 bl_1_37 bl_1_46 br_0_37 br_1_37 bl_1_38
+ br_0_38 br_0_32 br_1_38 br_1_32 br_1_46 bl_1_39 br_0_39 br_1_39 bl_1_47 br_0_47
+ br_0_40 br_1_40 br_0_41 br_1_41 br_0_33 br_1_47 br_0_42 br_1_42 br_0_43 br_1_33
+ br_1_43 br_0_44 br_1_44 bl_1_45 br_0_45 br_1_45 gnd_uq775 gnd_uq776 bl_1_3 bl_1_2
+ bl_1_1 wl_0_0 bl_1_0 bl_0_19 bl_0_29 bl_0_18 bl_0_39 bl_0_17 bl_0_28 wl_0_113 wl_0_102
+ wl_0_124 wl_0_36 wl_0_58 wl_0_47 wl_0_25 wl_0_14 bl_0_38 bl_0_49 bl_0_27 bl_0_16
+ wl_1_119 wl_0_123 wl_0_112 wl_0_101 wl_0_68 wl_0_57 wl_0_46 wl_0_35 wl_0_24 wl_0_13
+ bl_0_59 bl_0_48 bl_0_15 bl_0_26 bl_0_37 wl_0_122 wl_0_111 wl_0_100 wl_0_78 wl_0_67
+ wl_0_56 wl_0_45 wl_0_34 wl_0_23 wl_0_12 bl_0_47 bl_0_58 bl_0_36 bl_0_14 bl_0_25
+ wl_0_121 wl_0_110 wl_0_99 wl_0_88 wl_0_77 wl_0_66 wl_0_55 wl_0_44 wl_0_33 wl_0_22
+ wl_0_11 bl_0_57 bl_0_46 bl_0_24 bl_0_35 bl_0_13 wl_1_104 wl_0_120 wl_0_98 wl_0_87
+ wl_0_54 wl_0_76 wl_0_65 wl_0_43 wl_0_32 wl_0_21 wl_0_10 bl_0_56 bl_0_45 bl_0_23
+ bl_0_34 bl_0_12 wl_1_90 wl_0_97 wl_0_86 wl_0_75 wl_0_64 wl_0_20 wl_0_53 wl_0_42
+ wl_0_31 bl_0_44 bl_0_33 bl_0_55 bl_0_11 bl_0_22 wl_0_96 wl_0_74 wl_0_63 wl_0_85
+ wl_0_30 wl_0_52 wl_0_41 bl_0_32 bl_0_54 bl_0_43 bl_0_21 bl_0_10 wl_0_95 wl_0_84
+ wl_0_73 wl_0_62 wl_0_51 wl_0_40 bl_0_53 bl_0_42 bl_0_20 bl_0_31 wl_0_94 wl_0_83
+ wl_0_72 wl_0_50 wl_0_61 bl_0_41 bl_0_52 bl_0_63 bl_0_30 wl_1_115 wl_1_106 br_1_61
+ br_1_50 wl_0_93 wl_0_82 wl_0_71 wl_0_60 bl_0_51 bl_0_62 bl_0_40 bl_1_55 bl_1_33
+ bl_1_22 bl_1_44 bl_1_11 br_1_60 wl_0_92 wl_0_81 wl_0_70 bl_0_50 bl_0_61 bl_1_54
+ bl_1_21 bl_1_43 bl_1_32 bl_1_10 wl_1_5 wl_0_91 wl_0_69 wl_0_80 bl_0_60 bl_1_53 bl_1_31
+ bl_1_42 bl_1_20 wl_1_118 wl_1_109 wl_1_100 wl_0_90 wl_0_79 rbl_bl_1_1 bl_1_63 bl_1_52
+ bl_1_41 bl_1_30 wl_0_89 wl_1_127 wl_1_7 bl_1_62 bl_1_51 bl_1_40 wl_1_121 wl_1_112
+ bl_1_61 bl_1_50 wl_1_103 bl_1_60 wl_1_124 rbl_br_1_1 wl_1_18 wl_1_9 wl_1_57 wl_1_48
+ wl_1_39 wl_1_105 wl_1_21 wl_1_12 wl_1_33 wl_1_4 wl_1_117 wl_1_108 wl_1_99 br_1_9
+ br_0_9 br_1_8 bl_1_9 wl_1_24 wl_1_76 wl_1_15 br_0_8 wl_1_126 wl_1_6 wl_1_54 wl_0_8
+ bl_0_9 br_1_7 bl_1_8 wl_1_120 br_0_7 wl_1_111 wl_1_102 wl_0_7 bl_0_8 br_1_6 bl_1_7
+ br_0_6 wl_0_6 bl_0_7 br_1_5 wl_1_35 wl_1_68 bl_1_6 wl_1_88 wl_1_27 wl_1_79 wl_1_97
+ wl_1_29 br_0_5 wl_0_5 bl_0_6 br_1_4 bl_1_5 gnd vdd
Xsky130_sram_1kbyte_1rw1r_32x256_8_replica_column_0_0 wl_0_96 wl_0_97 wl_0_98 wl_0_99
+ wl_0_100 wl_0_101 wl_0_102 wl_0_103 wl_0_104 wl_0_105 wl_0_106 wl_0_107 wl_0_108
+ wl_0_109 wl_0_110 wl_0_111 wl_0_112 wl_0_113 wl_0_114 wl_0_115 wl_0_116 wl_0_117
+ wl_0_118 wl_0_119 wl_0_120 wl_0_121 wl_0_122 wl_0_123 wl_0_124 wl_0_125 wl_0_126
+ wl_0_127 gnd_uq776 wl_1_97 wl_1_98 wl_1_99 wl_1_100 wl_1_101 wl_1_102 wl_1_103 wl_1_105
+ wl_1_106 wl_1_107 wl_1_108 wl_1_109 wl_1_110 wl_1_111 wl_1_112 wl_1_113 wl_1_114
+ wl_1_115 wl_1_116 wl_1_117 wl_1_118 wl_1_119 wl_1_120 wl_1_121 wl_1_122 wl_1_123
+ wl_1_124 wl_1_125 wl_1_126 wl_1_127 rbl_wl_1_1 wl_1_64 wl_1_65 wl_1_66 wl_1_67 wl_1_68
+ wl_1_69 wl_1_70 wl_1_71 wl_1_72 wl_1_73 wl_1_74 wl_1_75 wl_1_76 wl_1_77 wl_1_78
+ wl_1_79 wl_1_80 wl_1_81 wl_1_82 wl_1_83 wl_1_84 wl_1_85 wl_1_86 wl_1_87 wl_1_88
+ wl_1_89 wl_1_90 wl_1_91 wl_1_92 wl_1_94 wl_1_95 wl_1_96 wl_0_65 wl_0_66 wl_0_67
+ wl_0_69 wl_0_70 wl_0_71 wl_0_72 wl_0_73 wl_0_74 wl_0_75 wl_0_76 wl_0_77 wl_0_78
+ wl_0_79 wl_0_80 wl_0_81 wl_0_82 wl_0_84 wl_0_85 wl_0_86 wl_0_87 wl_0_88 wl_0_89
+ wl_0_90 wl_0_91 wl_0_92 wl_0_93 wl_0_94 wl_0_95 wl_0_64 wl_0_32 wl_0_33 wl_0_34
+ wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43 wl_0_44
+ wl_0_45 wl_0_46 wl_0_47 wl_0_48 wl_0_49 wl_0_50 wl_0_52 wl_0_53 wl_0_54 wl_0_55
+ wl_0_56 wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_1_31 wl_1_32
+ wl_1_33 wl_1_34 wl_1_35 wl_1_36 wl_1_37 wl_1_38 wl_1_39 wl_1_40 wl_1_41 wl_1_42
+ wl_1_43 wl_1_44 wl_1_45 wl_1_46 wl_1_48 wl_1_49 wl_1_50 wl_1_51 wl_1_52 wl_1_53
+ wl_1_54 wl_1_55 wl_1_56 wl_1_57 wl_1_58 wl_1_59 wl_1_60 wl_1_61 wl_1_62 wl_1_63
+ gnd_uq775 wl_1_0 wl_1_1 wl_1_2 wl_1_3 wl_1_4 wl_1_5 wl_1_6 wl_1_7 wl_1_8 wl_1_9
+ wl_1_10 wl_1_11 wl_1_12 wl_1_13 wl_1_14 wl_1_15 wl_1_16 wl_1_17 wl_1_18 wl_1_19
+ wl_1_20 wl_1_21 wl_1_22 wl_1_23 wl_1_24 wl_1_25 wl_1_27 wl_1_28 wl_1_29 wl_1_30
+ wl_0_31 rbl_wl_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8
+ wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19
+ wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29
+ wl_0_30 vdd wl_1_104 wl_0_83 wl_0_68 wl_0_51 wl_1_26 wl_1_47 wl_1_93 rbl_bl_1_1
+ rbl_br_1_1 gnd rbl_bl_0_1 rbl_br_0_1 sky130_sram_1kbyte_1rw1r_32x256_8_replica_column_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_dummy_array_0 vdd bl_0_0 br_0_0 bl_1_0 br_1_0 bl_0_1
+ br_0_1 bl_1_1 br_1_1 bl_0_2 br_0_2 br_1_2 bl_0_3 br_0_3 bl_1_3 br_1_3 bl_0_4 br_0_4
+ bl_1_4 br_1_4 bl_0_5 br_0_5 bl_1_5 br_1_5 bl_0_6 br_0_6 bl_1_6 br_1_6 bl_0_7 br_0_7
+ bl_1_7 br_1_7 bl_0_8 br_0_8 bl_1_8 br_1_8 bl_0_9 br_0_9 bl_1_9 br_1_9 bl_0_10 br_0_10
+ bl_1_10 br_1_10 bl_0_11 br_0_11 bl_1_11 br_1_11 bl_0_12 br_0_12 bl_1_12 br_1_12
+ bl_0_13 br_0_13 bl_1_13 br_1_13 bl_0_14 br_0_14 bl_1_14 br_1_14 bl_0_15 br_0_15
+ bl_1_15 br_1_15 bl_0_16 br_0_16 bl_1_16 br_1_16 bl_0_17 br_0_17 bl_1_17 br_1_17
+ bl_0_18 br_0_18 bl_1_18 br_1_18 bl_0_19 br_0_19 bl_1_19 br_1_19 bl_0_20 br_0_20
+ br_1_20 bl_0_21 br_0_21 bl_1_21 br_1_21 bl_0_22 br_0_22 br_1_22 bl_0_23 br_0_23
+ bl_1_23 br_1_23 bl_0_24 br_0_24 bl_1_24 br_1_24 bl_0_25 br_0_25 bl_1_25 br_1_25
+ bl_0_26 br_0_26 bl_1_26 br_1_26 bl_0_27 br_0_27 bl_1_27 br_1_27 bl_0_28 br_0_28
+ bl_1_28 br_1_28 bl_0_29 br_0_29 bl_1_29 br_1_29 bl_0_30 br_0_30 bl_1_30 br_1_30
+ bl_0_31 br_0_31 bl_1_31 br_1_31 bl_0_32 br_0_32 bl_1_32 br_1_32 bl_0_33 br_0_33
+ br_1_33 bl_0_34 br_0_34 bl_1_34 br_1_34 br_0_35 bl_1_35 br_1_35 bl_0_36 br_0_36
+ bl_1_36 br_1_36 bl_0_37 br_0_37 bl_1_37 br_1_37 bl_0_38 br_0_38 bl_1_38 br_1_38
+ bl_0_39 br_0_39 bl_1_39 br_1_39 bl_0_40 br_0_40 br_1_40 bl_0_41 br_0_41 bl_1_41
+ br_1_41 bl_0_42 br_0_42 bl_1_42 br_1_42 bl_0_43 br_0_43 bl_1_43 br_1_43 bl_0_44
+ br_0_44 bl_1_44 br_1_44 bl_0_45 br_0_45 bl_1_45 br_1_45 bl_0_46 br_0_46 bl_1_46
+ br_1_46 bl_0_47 br_0_47 bl_1_47 br_1_47 bl_0_48 br_0_48 bl_1_48 br_1_48 bl_0_49
+ br_0_49 bl_1_49 br_1_49 bl_0_50 br_0_50 bl_1_50 br_1_50 bl_0_51 br_0_51 br_1_51
+ bl_0_52 br_0_52 bl_1_52 br_1_52 bl_0_53 br_0_53 br_1_53 bl_0_54 br_0_54 bl_1_54
+ br_1_54 bl_0_55 br_0_55 bl_1_55 br_1_55 bl_0_56 br_0_56 bl_1_56 br_1_56 bl_0_57
+ br_0_57 bl_1_57 br_1_57 bl_0_58 bl_1_58 br_1_58 bl_0_59 br_0_59 bl_1_59 br_1_59
+ bl_0_60 br_0_60 bl_1_60 br_1_60 bl_0_61 br_0_61 bl_1_61 br_1_61 bl_0_62 br_0_62
+ bl_1_62 br_1_62 bl_0_63 br_0_63 bl_1_63 br_1_63 vdd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd bl_1_63 br_1_19 bl_1_27
+ br_1_9 br_1_48 br_1_58 bl_1_31 br_1_38 bl_1_2 vdd bl_1_46 vdd br_1_28 vdd br_1_18
+ bl_1_50 bl_1_17 vdd br_1_8 br_1_47 br_1_57 bl_1_21 vdd br_1_37 vdd vdd bl_1_36 vdd
+ br_1_27 bl_1_54 vdd vdd bl_1_40 br_1_17 bl_1_7 vdd bl_1_58 br_1_7 br_1_46 br_1_56
+ bl_1_11 vdd br_1_36 bl_1_62 vdd vdd bl_1_26 vdd br_1_26 vdd vdd br_1_16 bl_1_30
+ vdd bl_1_51 br_1_6 bl_1_33 br_1_45 br_1_55 bl_1_1 bl_1_45 vdd br_1_35 vdd bl_1_49
+ vdd bl_1_16 vdd br_1_25 vdd vdd bl_1_53 bl_1_20 br_1_15 vdd br_1_44 br_1_5 br_1_54
+ bl_1_35 vdd br_1_34 bl_1_39 vdd vdd bl_1_6 vdd br_1_24 bl_1_57 vdd vdd bl_1_43 bl_1_10
+ br_1_14 vdd bl_0_35 bl_1_61 br_1_4 bl_1_25 vdd vdd bl_1_29 vdd vdd bl_1_20 bl_1_2
+ vdd bl_1_33 bl_1_0 bl_1_44 vdd br_1_53 br_1_63 bl_1_48 bl_1_15 vdd br_1_43 bl_1_52
+ vdd bl_1_19 vdd vdd br_1_33 vdd bl_1_23 br_1_23 bl_1_34 vdd br_1_13 br_1_52 br_1_62
+ bl_1_38 bl_1_5 vdd bl_1_53 br_1_3 br_1_42 bl_1_56 bl_1_42 bl_1_9 vdd vdd vdd br_1_32
+ bl_1_60 vdd bl_1_13 br_1_22 bl_1_24 vdd br_1_12 br_1_51 br_1_61 bl_1_28 vdd br_1_2
+ br_1_41 bl_1_32 vdd vdd vdd br_1_31 vdd bl_1_3 br_1_21 bl_1_47 bl_1_14 vdd br_1_11
+ br_0_58 br_1_50 br_1_60 bl_1_51 bl_1_18 vdd br_1_1 br_1_40 rbl_wl_1_1 bl_1_22 vdd
+ vdd vdd br_1_30 gnd_uq776 vdd bl_1_40 br_1_20 bl_1_37 bl_1_22 bl_1_4 vdd br_1_10
+ br_1_49 bl_1_55 br_1_59 bl_1_41 bl_1_8 vdd br_1_0 br_1_39 bl_1_59 gnd bl_1_12 vdd
+ br_1_29 sky130_sram_1kbyte_1rw1r_32x256_8_dummy_array
Xsky130_sram_1kbyte_1rw1r_32x256_8_dummy_array_1 vdd bl_0_0 br_0_0 bl_1_0 br_1_0 bl_0_1
+ br_0_1 bl_1_1 br_1_1 bl_0_2 br_0_2 br_1_2 bl_0_3 br_0_3 bl_1_3 br_1_3 bl_0_4 br_0_4
+ bl_1_4 br_1_4 bl_0_5 br_0_5 bl_1_5 br_1_5 bl_0_6 br_0_6 bl_1_6 br_1_6 bl_0_7 br_0_7
+ bl_1_7 br_1_7 bl_0_8 br_0_8 bl_1_8 br_1_8 bl_0_9 br_0_9 bl_1_9 br_1_9 bl_0_10 br_0_10
+ bl_1_10 br_1_10 bl_0_11 br_0_11 bl_1_11 br_1_11 bl_0_12 br_0_12 bl_1_12 br_1_12
+ bl_0_13 br_0_13 bl_1_13 br_1_13 bl_0_14 br_0_14 bl_1_14 br_1_14 bl_0_15 br_0_15
+ bl_1_15 br_1_15 bl_0_16 br_0_16 bl_1_16 br_1_16 bl_0_17 br_0_17 bl_1_17 br_1_17
+ bl_0_18 br_0_18 bl_1_18 br_1_18 bl_0_19 br_0_19 bl_1_19 br_1_19 bl_0_20 br_0_20
+ br_1_20 bl_0_21 br_0_21 bl_1_21 br_1_21 bl_0_22 br_0_22 br_1_22 bl_0_23 br_0_23
+ bl_1_23 br_1_23 bl_0_24 br_0_24 bl_1_24 br_1_24 bl_0_25 br_0_25 bl_1_25 br_1_25
+ bl_0_26 br_0_26 bl_1_26 br_1_26 bl_0_27 br_0_27 bl_1_27 br_1_27 bl_0_28 br_0_28
+ bl_1_28 br_1_28 bl_0_29 br_0_29 bl_1_29 br_1_29 bl_0_30 br_0_30 bl_1_30 br_1_30
+ bl_0_31 br_0_31 bl_1_31 br_1_31 bl_0_32 br_0_32 bl_1_32 br_1_32 bl_0_33 br_0_33
+ br_1_33 bl_0_34 br_0_34 bl_1_34 br_1_34 br_0_35 bl_1_35 br_1_35 bl_0_36 br_0_36
+ bl_1_36 br_1_36 bl_0_37 br_0_37 bl_1_37 br_1_37 bl_0_38 br_0_38 bl_1_38 br_1_38
+ bl_0_39 br_0_39 bl_1_39 br_1_39 bl_0_40 br_0_40 br_1_40 bl_0_41 br_0_41 bl_1_41
+ br_1_41 bl_0_42 br_0_42 bl_1_42 br_1_42 bl_0_43 br_0_43 bl_1_43 br_1_43 bl_0_44
+ br_0_44 bl_1_44 br_1_44 bl_0_45 br_0_45 bl_1_45 br_1_45 bl_0_46 br_0_46 bl_1_46
+ br_1_46 bl_0_47 br_0_47 bl_1_47 br_1_47 bl_0_48 br_0_48 bl_1_48 br_1_48 bl_0_49
+ br_0_49 bl_1_49 br_1_49 bl_0_50 br_0_50 bl_1_50 br_1_50 bl_0_51 br_0_51 br_1_51
+ bl_0_52 br_0_52 bl_1_52 br_1_52 bl_0_53 br_0_53 br_1_53 bl_0_54 br_0_54 bl_1_54
+ br_1_54 bl_0_55 br_0_55 bl_1_55 br_1_55 bl_0_56 br_0_56 bl_1_56 br_1_56 bl_0_57
+ br_0_57 bl_1_57 br_1_57 bl_0_58 bl_1_58 br_1_58 bl_0_59 br_0_59 bl_1_59 br_1_59
+ bl_0_60 br_0_60 bl_1_60 br_1_60 bl_0_61 br_0_61 bl_1_61 br_1_61 bl_0_62 br_0_62
+ bl_1_62 br_1_62 bl_0_63 br_0_63 bl_1_63 br_1_63 vdd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd bl_1_63 br_1_19 bl_1_27
+ br_1_9 br_1_48 br_1_58 bl_1_31 br_1_38 bl_1_2 vdd bl_1_46 vdd br_1_28 vdd br_1_18
+ bl_1_50 bl_1_17 vdd br_1_8 br_1_47 br_1_57 bl_1_21 vdd br_1_37 vdd vdd bl_1_36 vdd
+ br_1_27 bl_1_54 vdd vdd bl_1_40 br_1_17 bl_1_7 vdd bl_1_58 br_1_7 br_1_46 br_1_56
+ bl_1_11 vdd br_1_36 bl_1_62 vdd vdd bl_1_26 vdd br_1_26 vdd vdd br_1_16 bl_1_30
+ vdd bl_1_51 br_1_6 bl_1_33 br_1_45 br_1_55 bl_1_1 bl_1_45 vdd br_1_35 vdd bl_1_49
+ vdd bl_1_16 vdd br_1_25 vdd vdd bl_1_53 bl_1_20 br_1_15 vdd br_1_44 br_1_5 br_1_54
+ bl_1_35 vdd br_1_34 bl_1_39 vdd vdd bl_1_6 vdd br_1_24 bl_1_57 vdd vdd bl_1_43 bl_1_10
+ br_1_14 vdd bl_0_35 bl_1_61 br_1_4 bl_1_25 vdd vdd bl_1_29 vdd vdd bl_1_20 bl_1_2
+ vdd bl_1_33 bl_1_0 bl_1_44 vdd br_1_53 br_1_63 bl_1_48 bl_1_15 vdd br_1_43 bl_1_52
+ vdd bl_1_19 vdd vdd br_1_33 vdd bl_1_23 br_1_23 bl_1_34 vdd br_1_13 br_1_52 br_1_62
+ bl_1_38 bl_1_5 vdd bl_1_53 br_1_3 br_1_42 bl_1_56 bl_1_42 bl_1_9 vdd vdd vdd br_1_32
+ bl_1_60 vdd bl_1_13 br_1_22 bl_1_24 vdd br_1_12 br_1_51 br_1_61 bl_1_28 vdd br_1_2
+ br_1_41 bl_1_32 vdd vdd vdd br_1_31 vdd bl_1_3 br_1_21 bl_1_47 bl_1_14 vdd br_1_11
+ br_0_58 br_1_50 br_1_60 bl_1_51 bl_1_18 vdd br_1_1 br_1_40 gnd_uq775 bl_1_22 vdd
+ vdd vdd br_1_30 rbl_wl_0_0 vdd bl_1_40 br_1_20 bl_1_37 bl_1_22 bl_1_4 vdd br_1_10
+ br_1_49 bl_1_55 br_1_59 bl_1_41 bl_1_8 vdd br_1_0 br_1_39 bl_1_59 gnd bl_1_12 vdd
+ br_1_29 sky130_sram_1kbyte_1rw1r_32x256_8_dummy_array
Xsky130_sram_1kbyte_1rw1r_32x256_8_replica_column_0 wl_1_97 wl_1_98 wl_1_99 wl_1_105
+ wl_1_108 wl_1_111 wl_1_114 wl_1_117 wl_1_120 wl_1_122 wl_1_123 wl_1_126 wl_0_96
+ wl_0_102 wl_0_103 wl_0_104 wl_0_105 wl_0_106 wl_0_107 wl_0_108 wl_0_113 wl_0_114
+ wl_0_115 wl_0_116 wl_0_117 wl_0_118 wl_0_124 wl_0_125 wl_0_126 wl_0_127 gnd_uq776
+ wl_1_96 wl_0_66 wl_0_69 wl_0_75 wl_0_81 wl_0_84 wl_0_90 wl_1_64 wl_1_65 wl_1_66
+ wl_1_67 wl_1_68 wl_1_69 wl_1_70 wl_1_71 wl_1_73 wl_1_74 wl_1_75 wl_1_76 wl_1_77
+ wl_1_78 wl_1_79 wl_1_80 wl_1_81 wl_1_82 wl_1_83 wl_1_84 wl_1_85 wl_1_86 wl_1_87
+ wl_1_90 wl_1_91 wl_1_92 wl_1_94 wl_1_95 wl_0_36 wl_0_37 wl_0_38 wl_0_47 wl_0_48
+ wl_0_54 wl_0_58 wl_0_59 wl_0_62 wl_1_31 wl_1_32 wl_1_34 wl_1_35 wl_1_37 wl_1_38
+ wl_1_39 wl_1_40 wl_1_41 wl_1_43 wl_1_44 wl_1_46 wl_1_47 wl_1_49 wl_1_50 wl_1_52
+ wl_1_53 wl_1_54 wl_1_55 wl_1_57 wl_1_58 wl_1_59 wl_1_60 wl_1_61 wl_1_62 wl_1_0 wl_1_1
+ wl_1_2 wl_1_5 wl_1_8 wl_1_9 wl_1_10 wl_1_11 wl_1_13 wl_1_14 wl_1_16 wl_1_17 wl_1_19
+ wl_1_20 wl_1_22 wl_1_23 wl_1_25 wl_1_26 wl_1_28 wl_1_29 wl_0_0 wl_0_1 wl_0_2 wl_0_3
+ wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_25
+ wl_0_26 wl_0_27 wl_0_28 vdd wl_0_123 wl_0_87 wl_0_78 wl_0_35 wl_0_99 wl_0_29 wl_0_20
+ wl_0_11 wl_0_120 wl_0_111 wl_0_55 wl_0_50 wl_0_41 wl_0_92 wl_0_32 wl_0_23 wl_1_113
+ wl_1_104 wl_0_83 wl_0_74 wl_0_65 wl_0_122 wl_0_53 wl_0_44 wl_0_95 wl_1_7 wl_1_125
+ wl_1_116 wl_1_107 wl_0_86 wl_0_68 wl_0_77 wl_0_61 wl_0_98 wl_1_89 wl_1_119 wl_1_110
+ wl_1_101 wl_0_89 wl_0_80 wl_0_71 wl_0_46 wl_0_19 wl_0_10 wl_0_119 wl_0_110 wl_0_101
+ rbl_wl_1_1 wl_1_4 wl_0_49 wl_0_40 wl_0_31 wl_0_13 wl_0_22 wl_1_112 wl_1_103 wl_0_82
+ wl_0_73 wl_0_64 wl_0_57 wl_0_112 wl_0_52 wl_0_43 wl_0_34 wl_0_94 wl_1_15 wl_1_6
+ wl_1_124 wl_1_115 wl_1_106 wl_0_85 wl_0_76 wl_0_67 wl_0_60 wl_0_97 wl_1_88 wl_1_45
+ gnd_uq775 wl_1_36 wl_1_27 wl_1_18 wl_1_127 wl_1_118 wl_1_109 wl_1_100 wl_0_88 wl_0_79
+ wl_0_70 rbl_wl_0_0 wl_0_45 wl_0_9 wl_0_109 wl_0_100 wl_1_48 wl_1_30 wl_1_21 wl_1_12
+ wl_1_3 wl_1_121 wl_0_91 wl_0_39 wl_0_30 wl_0_21 wl_0_12 wl_0_121 wl_1_72 wl_1_63
+ wl_1_56 wl_1_51 wl_1_102 wl_1_42 wl_1_93 wl_1_33 wl_1_24 wl_0_72 wl_0_63 wl_0_56
+ wl_0_51 wl_0_42 wl_0_33 wl_0_93 wl_0_24 rbl_bl_1_0 rbl_br_1_0 rbl_br_0_0 rbl_bl_0_0
+ gnd sky130_sram_1kbyte_1rw1r_32x256_8_replica_column
Xsky130_sram_1kbyte_1rw1r_32x256_8_bitcell_array_0 wl_0_125 wl_1_80 wl_1_81 wl_0_59
+ wl_0_48 wl_0_49 wl_1_51 wl_0_37 wl_0_28 wl_0_26 wl_0_19 wl_0_15 wl_0_4 br_1_30 br_0_19
+ bl_1_12 bl_1_4 bl_1_5 bl_1_56 bl_1_57 br_1_51 bl_1_45 br_1_40 br_1_41 bl_1_37 bl_1_34
+ gnd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ br_1_54 br_1_5 br_1_37 br_1_63 bl_1_59 bl_1_22 bl_1_56 bl_1_62 bl_1_41 br_1_22 bl_1_28
+ bl_1_32 br_1_33 bl_1_9 bl_1_21 bl_1_11 bl_1_60 br_1_38 br_1_49 bl_1_47 bl_1_29 bl_1_11
+ bl_1_9 bl_1_40 bl_1_45 br_1_25 br_1_63 br_1_35 br_1_0 br_1_19 br_1_17 br_1_44 bl_1_2
+ br_1_37 bl_1_15 bl_1_58 br_1_26 bl_1_15 br_1_16 bl_1_46 br_1_59 br_1_20 br_1_59
+ br_1_61 br_1_24 bl_1_14 br_1_47 br_1_49 br_1_53 bl_1_58 bl_1_31 bl_1_34 br_1_51
+ br_1_51 br_1_55 br_1_21 br_1_27 bl_1_25 br_1_7 bl_1_5 bl_1_17 br_1_52 br_1_18 bl_1_14
+ bl_1_27 bl_1_24 br_1_9 br_1_10 br_1_58 br_1_30 bl_1_31 bl_1_20 bl_1_4 bl_1_52 bl_1_54
+ br_1_34 bl_1_19 br_1_34 br_1_32 bl_1_4 bl_1_34 br_1_30 br_1_23 br_1_28 bl_1_40 bl_1_33
+ br_1_60 bl_1_38 br_1_13 bl_1_1 bl_1_56 bl_1_39 br_1_43 br_1_38 br_1_17 br_1_22 br_1_24
+ br_1_6 br_1_50 br_1_39 bl_1_25 bl_1_0 bl_1_16 br_1_56 br_1_2 bl_1_43 br_1_40 br_1_1
+ bl_1_47 br_1_3 bl_1_3 bl_1_35 br_1_31 bl_1_2 br_1_5 bl_1_10 bl_1_43 bl_1_29 br_1_4
+ br_1_18 br_1_27 br_1_28 bl_1_6 bl_1_45 br_1_44 bl_1_57 br_1_42 bl_1_42 br_1_12 br_1_57
+ bl_1_7 br_1_57 br_1_29 br_1_11 br_1_56 br_1_15 br_1_13 bl_1_30 br_1_11 br_1_41 bl_1_28
+ bl_1_10 br_1_21 br_1_48 bl_1_5 bl_1_60 bl_1_55 bl_1_7 bl_1_26 br_1_9 br_1_45 bl_1_49
+ br_1_60 br_1_15 br_1_2 br_1_14 bl_1_33 bl_1_50 br_1_33 bl_1_63 br_1_46 bl_1_51 bl_1_61
+ bl_1_50 br_1_41 bl_1_53 bl_1_12 bl_1_37 br_1_62 bl_1_3 bl_1_0 bl_1_44 br_1_25 br_1_40
+ br_1_55 br_1_52 bl_1_53 bl_1_52 br_1_29 br_1_23 br_1_10 bl_1_54 bl_1_37 bl_1_38
+ bl_1_48 bl_1_17 bl_1_8 br_1_50 br_1_8 bl_1_49 bl_1_35 bl_1_13 br_1_53 bl_1_57 bl_1_59
+ br_1_14 bl_1_44 br_1_12 br_1_7 bl_1_36 br_1_4 br_1_42 bl_1_13 br_1_58 br_1_32 br_1_47
+ br_1_45 bl_1_55 br_1_1 bl_1_62 bl_1_26 br_1_54 bl_1_8 br_1_36 bl_1_22 br_1_48 bl_1_23
+ bl_1_32 bl_1_16 bl_1_46 bl_1_61 wl_0_83 br_1_50 wl_1_28 bl_1_6 wl_1_19 wl_1_113
+ wl_1_4 wl_1_0 br_0_50 wl_1_98 br_1_6 wl_1_46 br_1_36 bl_1_51 br_1_26 br_1_19 wl_0_67
+ wl_0_113 br_1_61 wl_1_86 wl_0_78 bl_0_34 br_1_31 wl_0_0 bl_1_48 br_1_39 wl_0_98
+ wl_1_40 wl_0_60 bl_0_10 wl_0_46 br_1_20 wl_1_58 wl_1_107 bl_1_18 bl_1_50 bl_1_1
+ wl_1_49 wl_1_10 wl_0_9 br_1_8 wl_1_76 wl_1_64 wl_0_65 bl_1_24 wl_0_86 bl_0_23 br_1_3
+ bl_1_41 bl_1_63 wl_1_43 bl_0_37 wl_1_123 wl_0_40 bl_0_56 bl_1_18 bl_1_16 wl_0_58
+ wl_1_125 wl_0_107 bl_1_19 bl_0_50 wl_0_10 wl_1_116 wl_1_97 br_1_21 wl_0_29 br_1_38
+ wl_1_13 bl_0_1 wl_0_8 wl_0_34 bl_0_7 wl_0_76 wl_0_63 wl_0_95 br_0_52 br_1_18 wl_0_64
+ bl_1_23 bl_1_6 bl_1_31 bl_0_45 wl_0_93 br_1_25 bl_0_2 wl_1_75 wl_1_20 wl_1_29 bl_1_42
+ wl_0_43 br_1_4 bl_0_53 wl_1_110 br_0_8 br_1_0 bl_0_40 wl_1_36 br_0_32 wl_0_22 wl_0_74
+ bl_1_63 wl_1_120 vdd wl_0_123 bl_0_58 wl_1_54 bl_1_51 bl_1_49 wl_0_69 bl_0_8 bl_1_61
+ wl_1_56 br_1_62 br_1_45 wl_0_106 br_0_56 bl_1_36 wl_1_79 bl_0_35 br_1_60 wl_1_101
+ bl_0_16 wl_1_35 bl_0_43 wl_0_104 wl_0_105 bl_1_0 br_1_2 wl_1_100 wl_0_116 wl_0_108
+ wl_1_42 bl_1_3 wl_0_97 br_1_9 wl_1_31 br_1_59 wl_0_7 wl_1_90 wl_0_52 br_1_31 wl_1_119
+ wl_1_114 br_1_0 wl_1_99 br_1_12 br_0_26 br_0_24 bl_0_44 br_0_21 br_1_39 bl_1_12
+ wl_1_111 br_0_38 wl_1_84 wl_0_13 br_0_36 wl_1_89 br_0_37 bl_1_39 br_1_58 bl_1_27
+ bl_1_20 wl_1_9 bl_0_14 bl_0_47 bl_0_25 wl_0_32 wl_1_68 bl_0_5 bl_0_17 wl_1_17 wl_0_25
+ br_0_18 br_1_16 wl_1_77 br_1_53 bl_0_9 bl_0_6 bl_1_46 bl_0_59 bl_0_31 bl_1_38 br_1_63
+ br_0_33 wl_1_27 wl_1_2 br_0_42 wl_1_12 bl_1_41 br_0_28 bl_1_19 wl_0_47 bl_1_18 wl_0_87
+ br_0_23 br_0_25 wl_0_66 bl_0_13 wl_0_6 wl_1_3 wl_0_45 wl_1_117 wl_1_1 wl_1_112 wl_0_75
+ wl_0_20 bl_1_39 bl_1_33 wl_0_38 br_1_3 wl_1_50 bl_0_42 wl_1_11 wl_0_36 wl_1_103
+ br_1_20 br_0_30 wl_0_61 wl_0_16 bl_0_4 wl_0_55 br_0_4 wl_1_32 wl_1_122 wl_1_14 wl_1_18
+ wl_0_110 wl_1_108 bl_1_30 bl_1_30 bl_0_60 wl_0_57 bl_1_17 bl_0_11 br_0_43 wl_1_126
+ br_1_43 wl_1_30 bl_0_54 wl_0_24 br_1_23 bl_0_32 br_0_6 bl_0_63 br_1_26 wl_1_87 wl_0_80
+ br_1_29 br_0_34 br_0_47 wl_0_120 br_1_49 br_1_46 bl_0_12 bl_1_7 wl_1_88 br_1_35
+ bl_1_27 wl_0_54 wl_1_109 bl_0_51 bl_0_49 br_1_44 bl_1_35 wl_0_71 wl_1_105 br_0_11
+ wl_1_121 br_0_41 wl_1_45 wl_0_94 bl_0_62 bl_1_48 wl_1_24 wl_1_63 wl_1_61 wl_1_62
+ wl_0_127 bl_1_32 bl_0_61 br_0_31 wl_1_106 br_0_29 wl_0_56 br_1_34 bl_0_48 br_0_45
+ br_1_27 wl_0_51 wl_0_85 br_1_22 wl_1_52 wl_0_102 br_0_14 wl_1_78 wl_0_118 br_1_19
+ wl_1_5 wl_0_5 br_0_51 wl_0_88 wl_0_44 br_0_46 bl_1_15 wl_0_79 br_0_48 br_0_60 wl_0_101
+ wl_1_92 wl_0_70 wl_0_109 br_1_46 wl_1_94 wl_1_47 wl_0_35 wl_1_60 wl_0_33 wl_0_62
+ wl_1_127 br_1_42 br_0_10 bl_1_14 wl_1_83 wl_1_33 bl_0_0 wl_0_100 br_0_2 wl_1_104
+ wl_1_85 br_1_17 wl_0_92 wl_0_42 vdd wl_0_39 br_0_61 bl_0_3 wl_1_7 wl_1_95 br_0_54
+ wl_0_53 bl_0_52 br_0_9 wl_0_31 br_0_13 br_0_59 br_1_7 bl_1_10 wl_0_90 bl_1_47 bl_1_52
+ bl_1_11 br_1_24 bl_1_36 wl_0_119 bl_0_24 bl_1_55 bl_0_28 br_0_49 wl_1_102 wl_0_114
+ wl_1_53 bl_1_21 br_1_28 br_0_0 wl_0_99 br_0_12 wl_0_72 wl_1_23 br_1_8 wl_0_81 bl_0_15
+ br_0_39 wl_0_111 br_1_33 bl_1_53 wl_1_8 br_1_57 bl_0_26 br_1_10 br_0_57 wl_0_84
+ br_1_55 wl_0_89 wl_0_122 bl_1_13 bl_0_29 bl_0_39 br_1_62 wl_0_73 br_0_7 wl_1_74
+ br_0_58 bl_0_27 br_0_55 bl_1_20 bl_1_1 wl_0_14 bl_0_20 wl_1_59 br_1_5 wl_1_70 bl_1_24
+ wl_1_26 wl_0_68 bl_0_30 wl_1_65 br_1_16 bl_1_9 br_1_32 wl_0_91 bl_1_8 br_1_61 br_1_37
+ br_0_5 bl_0_57 wl_0_17 wl_1_38 wl_1_91 br_1_47 bl_1_54 wl_1_66 bl_0_36 wl_1_71 br_0_16
+ bl_0_21 br_1_48 wl_1_41 wl_1_22 wl_0_77 wl_0_82 br_0_53 wl_0_23 bl_1_2 bl_1_26 br_1_56
+ wl_0_21 wl_1_82 wl_1_44 bl_0_46 br_1_11 br_1_13 bl_0_38 wl_1_118 br_0_63 wl_1_6
+ br_0_1 bl_1_62 bl_1_22 bl_1_42 wl_1_21 wl_1_39 wl_0_27 wl_1_93 wl_1_124 wl_0_2 br_0_27
+ bl_1_25 wl_0_12 wl_1_73 wl_0_126 br_1_43 bl_1_43 bl_0_41 wl_1_69 br_1_52 bl_0_19
+ wl_0_96 br_0_22 wl_0_41 br_0_62 bl_0_22 bl_0_18 bl_1_21 vdd br_1_14 br_1_6 wl_0_18
+ wl_1_34 wl_1_48 wl_1_115 bl_1_59 wl_0_3 br_0_15 wl_0_117 wl_0_121 wl_1_96 br_1_15
+ wl_0_1 wl_0_112 br_1_36 wl_0_124 bl_0_33 bl_1_40 br_0_3 bl_1_29 wl_1_25 wl_1_72
+ br_0_40 wl_1_15 wl_1_37 br_0_17 wl_0_30 br_0_35 br_1_54 wl_0_50 wl_1_57 vdd wl_0_11
+ bl_1_58 br_1_35 bl_1_28 br_0_44 bl_1_23 bl_1_44 wl_0_103 br_0_20 bl_1_60 bl_0_55
+ wl_1_55 wl_0_115 wl_1_16 vdd wl_1_67 br_1_1 sky130_sram_1kbyte_1rw1r_32x256_8_bitcell_array
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_port_address wl_en addr_0 addr_1 addr_2
+ addr_3 addr_4 addr_5 addr_6 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72
+ wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86
+ wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100
+ wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112
+ wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124
+ wl_125 wl_126 wl_127 rbl_wl wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11
+ wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25
+ wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39
+ wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53
+ wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_0 vdd_uq2 vdd_uq3
+ vdd_uq78 vdd_uq76 vdd_uq8 vdd vdd_uq406 vdd_uq407 gnd_uq8 gnd_uq9 gnd_uq3 gnd_uq20
+ gnd_uq25 gnd_uq26 vdd_uq35 vdd_uq27 vdd_uq51 vdd_uq4 gnd_uq37 vdd_uq34 gnd vdd_uq405
Xsky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0 addr_0 addr_1 addr_2 addr_3
+ addr_4 addr_5 addr_6 sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_1 sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_2
+ sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_3 sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_4
+ sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_5 sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_6
+ sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_7 sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_8
+ sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_9 sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_10
+ sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_11 sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_12
+ sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_13 sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_14
+ sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder_0/predecode_15 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_64
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_65 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_66
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_67 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_68
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_69 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_70
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_71 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_72
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_73 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_74
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_75 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_76
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_77 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_78
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_79 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_80
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_81 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_82
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_83 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_84
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_85 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_86
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_87 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_88
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_89 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_90
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_91 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_92
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_93 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_94
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_95 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_96
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_97 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_98
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_99 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_100
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_101 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_102
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_103 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_104
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_105 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_106
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_107 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_108
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_109 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_110
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_111 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_112
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_113 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_114
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_115 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_116
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_117 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_118
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_119 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_120
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_121 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_122
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_123 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_124
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_125 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_126
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_0 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_2 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_3
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_4 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_5
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_6 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_7
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_8 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_9
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_10 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_11
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_12 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_13
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_14 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_15
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_16 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_17
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_18 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_19
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_20 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_21
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_22 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_23
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_24 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_25
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_26 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_27
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_28 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_29
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_30 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_31
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_32 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_33
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_34 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_35
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_36 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_37
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_38 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_39
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_40 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_41
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_42 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_43
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_44 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_45
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_46 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_47
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_48 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_49
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_50 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_51
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_52 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_53
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_54 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_55
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_56 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_57
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_58 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_59
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_60 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_61
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_62 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_63
+ vdd_uq2 vdd_uq3 vdd_uq34 vdd_uq35 vdd_uq27 vdd_uq76 vdd_uq8 gnd_uq8 gnd_uq3 gnd_uq9
+ gnd_uq25 gnd_uq26 gnd_uq20 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_127
+ vdd_uq78 vdd_uq51 vdd_uq4 gnd_uq37 vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_hierarchical_decoder
Xsky130_sram_1kbyte_1rw1r_32x256_8_and2_dec_0_0 wl_en vdd_uq407 vdd_uq405 vdd_uq406
+ gnd rbl_wl sky130_sram_1kbyte_1rw1r_32x256_8_and2_dec_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0 wl_en wl_64 wl_65 wl_66
+ wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80
+ wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94
+ wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107
+ wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119
+ wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_96
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_80 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_97
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_98 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_81
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_99 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_100
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_82 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_101
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_102 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_83
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_103 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_104
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_84 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_105
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_74 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_85
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_86 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_75
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_110 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_87
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_65 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_88
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_76 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_90
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_77 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_91
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_92 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_121
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_78 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_93
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_79 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_95
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_64 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_6
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_7 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_8
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_9 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_10
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_11 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_12
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_13 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_14
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_15 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_16
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_20 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_34
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_35 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_36
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_37 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_38
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_39 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_40
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_41 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_42
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_43 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_44
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_45 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_46
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_47 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_50
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_51 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_62
+ wl_0 wl_32 wl_16 wl_33 wl_8 wl_34 wl_17 wl_35 wl_4 wl_36 wl_18 wl_37 wl_9 wl_38
+ wl_19 wl_39 wl_2 wl_40 wl_20 wl_41 wl_10 wl_42 wl_21 wl_43 wl_5 wl_44 wl_22 wl_45
+ wl_11 wl_46 wl_23 wl_47 wl_1 wl_48 wl_24 wl_49 wl_12 wl_50 wl_25 wl_51 wl_6 wl_52
+ wl_26 wl_53 wl_13 wl_54 wl_27 wl_55 wl_3 wl_56 wl_28 wl_57 wl_14 wl_58 wl_29 wl_59
+ wl_7 wl_60 wl_30 wl_61 wl_15 wl_62 wl_31 wl_63 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_106
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_17 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_107
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_18 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_108
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_48 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_19
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_109 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_49
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_27 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_89
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_111 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_28
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_21 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_122
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_112 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_29
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_22 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_123
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_113 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_52
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_30 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_23
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_124 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_114
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_53 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_2
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_24 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_125
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_54 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_115
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_3 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_25
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_126 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_94
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_55 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_116
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_4 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_26
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_127 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_56
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_117 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_68 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_66
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_57 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_118
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_1 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_69
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_67 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_58
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_119 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_5
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_70 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_31
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_59 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_71
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_120 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_63
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_32 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_60
+ sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_72 vdd_uq406 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_33
+ vdd_uq405 sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_61 gnd sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array_0/in_73
+ gnd sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_array
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_bank rbl_bl_1_1 rbl_bl_0_0 p_en_bar0 s_en0
+ w_en0 wl_en0 s_en1 p_en_bar1 wl_en1 bank_wmask0_0 bank_wmask0_1 bank_wmask0_2 bank_wmask0_3
+ dout1_16 dout1_17 dout1_18 dout1_19 dout1_20 dout1_21 dout1_22 dout1_23 dout1_24
+ dout1_25 dout1_26 dout1_27 dout1_28 dout1_29 dout1_30 dout1_31 dout1_0 dout1_1 dout1_2
+ dout1_3 dout1_4 dout1_5 dout1_6 dout1_7 dout1_8 dout1_9 dout1_10 dout1_11 dout1_12
+ dout1_13 dout1_14 dout1_15 addr0_1 addr0_2 addr0_3 addr0_4 addr0_5 din0_0 din0_1
+ din0_2 din0_3 din0_4 din0_5 din0_6 din0_7 din0_8 din0_9 din0_10 din0_11 din0_12
+ din0_13 din0_14 din0_15 dout0_0 dout0_1 dout0_2 dout0_3 dout0_4 dout0_5 dout0_6
+ dout0_7 dout0_8 dout0_9 dout0_10 dout0_11 dout0_12 dout0_13 dout0_14 dout0_15 din0_23
+ din0_24 din0_25 din0_26 din0_27 din0_28 din0_29 din0_30 din0_31 dout0_16 dout0_17
+ dout0_18 dout0_19 dout0_20 dout0_21 dout0_22 dout0_23 dout0_24 dout0_25 dout0_26
+ dout0_27 dout0_28 dout0_29 dout0_30 dout0_31 din0_16 din0_17 din0_18 din0_19 din0_20
+ din0_22 addr1_1 addr1_2 addr1_3 addr1_4 addr1_5 addr1_6 addr1_7 addr0_0 addr1_0
+ gnd_uq1 gnd_uq2 gnd_uq3 gnd_uq4 gnd_uq5 gnd_uq6 gnd_uq7 gnd_uq8 gnd_uq9 gnd_uq10
+ gnd_uq12 gnd_uq13 gnd_uq14 gnd_uq15 gnd_uq16 gnd_uq17 gnd_uq18 gnd_uq19 gnd_uq20
+ gnd_uq21 gnd_uq22 gnd_uq23 gnd_uq24 gnd_uq25 gnd_uq26 gnd_uq27 gnd_uq28 gnd_uq29
+ gnd_uq30 gnd_uq31 gnd_uq32 gnd_uq194 gnd_uq199 gnd_uq208 gnd_uq220 gnd_uq225 gnd_uq226
+ gnd_uq251 gnd_uq260 gnd_uq278 gnd_uq303 gnd_uq1132 gnd_uq1229 gnd_uq1230 gnd_uq1231
+ gnd_uq1232 vdd vdd_uq9 vdd_uq66 vdd_uq67 vdd_uq68 vdd_uq69 vdd_uq70 vdd_uq71 vdd_uq72
+ vdd_uq73 vdd_uq74 vdd_uq75 vdd_uq76 vdd_uq77 vdd_uq78 vdd_uq79 vdd_uq80 vdd_uq81
+ vdd_uq82 vdd_uq83 vdd_uq84 vdd_uq85 vdd_uq86 vdd_uq87 vdd_uq88 vdd_uq89 vdd_uq90
+ vdd_uq91 vdd_uq92 vdd_uq93 vdd_uq94 vdd_uq95 vdd_uq96 vdd_uq262 vdd_uq263 vdd_uq282
+ vdd_uq289 vdd_uq290 vdd_uq309 vdd_uq328 vdd_uq355 vdd_uq420 vdd_uq422 vdd_uq413
+ vdd_uq998 vdd_uq994 vdd_uq999 vdd_uq996 vdd_uq1075 vdd_uq1241 vdd_uq1242 vdd_uq1243
+ vdd_uq1244 vdd_uq1245 vdd_uq1246 vdd_uq1247 vdd_uq1248 vdd_uq1249 vdd_uq1250 vdd_uq1251
+ vdd_uq1252 vdd_uq1253 vdd_uq1254 vdd_uq1255 vdd_uq1256 vdd_uq1257 vdd_uq1258 vdd_uq1259
+ vdd_uq1260 vdd_uq1261 vdd_uq1262 vdd_uq1263 vdd_uq1264 vdd_uq1265 vdd_uq1266 vdd_uq1267
+ vdd_uq1268 vdd_uq1269 vdd_uq1270 vdd_uq1271 vdd_uq1272 vdd_uq1273 vdd_uq1274 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/gnd_uq26
+ vdd_uq281 din0_21 vdd_uq327 gnd_uq272 vdd_uq336 vdd_uq65 vdd_uq320 vdd_uq335 vdd_uq1208
+ vdd_uq368 addr0_7 addr0_6 gnd_uq11 vdd_uq99 vdd_uq64 vdd_uq274 vdd_uq693 gnd_uq312
+ vdd_uq691 vdd_uq690 vdd_uq1240 vdd_uq193 vdd_uq412 vdd_uq692 vdd_uq259 gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinvbuf_0 gnd_uq1230 sky130_sram_1kbyte_1rw1r_32x256_8_pinvbuf_0/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinvbuf_0/Zb addr0_0 gnd_uq1229 vdd_uq1273 sky130_sram_1kbyte_1rw1r_32x256_8_pinvbuf
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinvbuf_1 gnd_uq1231 sky130_sram_1kbyte_1rw1r_32x256_8_pinvbuf_1/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinvbuf_1/Zb addr1_0 gnd_uq1232 vdd_uq1274 sky130_sram_1kbyte_1rw1r_32x256_8_pinvbuf
Xsky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0 wl_en1 addr1_1 addr1_2 addr1_3
+ addr1_4 addr1_5 addr1_6 addr1_7 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_65
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_66 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_67
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_68 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_69
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_70 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_71
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_72 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_73
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_74 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_75
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_76 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_77
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_78 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_79
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_80 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_81
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_82 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_83
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_84 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_85
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_86 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_87
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_88 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_89
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_90 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_91
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_92 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_93
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_94 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_95
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_96 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_97
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_98 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_99
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_100 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_101
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_102 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_103
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_104 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_105
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_106 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_107
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_108 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_109
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_110 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_111
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_112 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_113
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_114 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_115
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_116 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_117
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_118 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_119
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_120 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_121
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_122 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_123
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_124 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_125
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_126 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_127
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/rbl_wl sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_64
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_0 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_2 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_3
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_4 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_5
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_6 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_7
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_8 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_9
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_10 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_11
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_12 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_13
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_14 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_15
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_16 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_17
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_18 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_19
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_20 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_21
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_22 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_23
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_24 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_25
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_26 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_27
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_28 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_29
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_30 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_31
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_32 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_33
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_34 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_35
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_36 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_37
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_38 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_39
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_40 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_41
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_42 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_43
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_44 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_45
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_46 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_47
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_48 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_49
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_50 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_51
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_52 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_53
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_54 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_55
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_56 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_57
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_58 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_59
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_60 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_61
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_62 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_63
+ vdd_uq282 vdd_uq263 vdd_uq413 vdd_uq999 vdd_uq998 vdd_uq690 vdd_uq1075 gnd_uq220
+ gnd_uq199 gnd_uq251 gnd_uq272 vdd_uq412 vdd_uq327 vdd_uq309 vdd_uq355 gnd_uq303
+ vdd_uq328 vdd_uq281 gnd vdd_uq691 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_port_data_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinvbuf_0/Zb
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinvbuf_0/Z bank_wmask0_0 bank_wmask0_1 bank_wmask0_2
+ bank_wmask0_3 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/wdriver_sel_2 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/wdriver_sel_3
+ din0_16 din0_17 din0_19 din0_20 din0_21 din0_22 din0_23 din0_24 din0_25 din0_26
+ din0_27 din0_28 din0_29 din0_30 din0_31 dout0_16 dout0_17 dout0_18 dout0_19 dout0_20
+ dout0_21 dout0_22 dout0_23 dout0_24 dout0_25 dout0_26 dout0_27 dout0_28 dout0_29
+ dout0_30 dout0_31 din0_12 din0_13 dout0_0 dout0_1 dout0_2 dout0_3 dout0_4 dout0_5
+ dout0_6 dout0_7 dout0_8 dout0_9 dout0_10 dout0_11 dout0_12 dout0_13 dout0_14 dout0_15
+ din0_14 din0_15 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/wdriver_sel_0 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/wdriver_sel_1
+ din0_0 din0_1 din0_2 din0_3 din0_4 din0_5 din0_6 din0_7 din0_8 din0_9 din0_10 din0_11
+ rbl_bl_0_0 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/rbl_br sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_0 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_1 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_2
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_2 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_3
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_3 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_4
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_4 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_5
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_5 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_6
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_6 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_7
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_7 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_8
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_8 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_9
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_9 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_10
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_10 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_11
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_11 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_12
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_12 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_13
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_13 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_14
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_14 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_15
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_15 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_16
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_16 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_17
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_17 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_18
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_18 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_19
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_19 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_20
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_20 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_21
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_21 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_22
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_22 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_23
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_23 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_24
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_24 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_25
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_25 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_26
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_26 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_27
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_27 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_28
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_28 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_29
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_29 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_30
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_30 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_31
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_31 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_32
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_32 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_33
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_33 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_34
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_34 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_35
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_35 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_36
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_36 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_37
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_37 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_38
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_38 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_39
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_39 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_40
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_40 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_41
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_41 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_42
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_42 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_43
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_43 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_44
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_44 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_45
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_45 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_46
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_46 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_47
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_47 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_48
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_48 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_49
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_49 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_50
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_50 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_51
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_51 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_52
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_52 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_53
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_53 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_54
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_54 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_55
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_55 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_56
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_56 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_57
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_57 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_58
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_58 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_59
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_59 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_60
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_60 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_61
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_61 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_62
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_62 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_63
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_63 vdd_uq193 vdd_uq65 vdd_uq66
+ vdd_uq67 vdd_uq69 vdd_uq70 vdd_uq71 vdd_uq72 vdd_uq73 vdd_uq74 vdd_uq75 vdd_uq76
+ vdd_uq77 vdd_uq78 vdd_uq79 vdd_uq80 vdd_uq81 vdd_uq82 vdd_uq83 vdd_uq84 vdd_uq85
+ vdd_uq86 vdd_uq87 vdd_uq88 vdd_uq89 vdd_uq90 vdd_uq91 vdd_uq92 vdd_uq93 vdd_uq94
+ vdd_uq95 vdd_uq96 vdd_uq64 gnd_uq1 gnd_uq2 gnd_uq3 gnd_uq4 gnd_uq5 gnd_uq6 gnd_uq7
+ gnd_uq8 gnd_uq9 gnd_uq10 gnd_uq11 gnd_uq12 gnd_uq13 gnd_uq14 gnd_uq15 gnd_uq16 gnd_uq17
+ gnd_uq18 gnd_uq19 gnd_uq20 gnd_uq21 gnd_uq22 gnd_uq23 gnd_uq24 gnd_uq25 gnd_uq26
+ gnd_uq27 gnd_uq28 gnd_uq29 gnd_uq30 gnd_uq31 gnd_uq32 din0_18 vdd vdd_uq9 vdd_uq99
+ w_en0 s_en0 vdd_uq68 gnd p_en_bar0 sky130_sram_1kbyte_1rw1r_32x256_8_port_data
Xsky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinvbuf_1/Zb
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinvbuf_1/Z dout1_17 dout1_18 dout1_19 dout1_20
+ dout1_21 dout1_22 dout1_23 dout1_24 dout1_25 dout1_26 dout1_27 dout1_28 dout1_29
+ dout1_30 dout1_31 dout1_15 dout1_16 dout1_0 dout1_1 dout1_2 dout1_3 dout1_4 dout1_5
+ dout1_6 dout1_7 dout1_8 dout1_9 dout1_10 dout1_11 dout1_12 dout1_13 dout1_14 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_0 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_1 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_2
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_2 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_3
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_3 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_4
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_4 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_5
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_5 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_6
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_6 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_7
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_7 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_8
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_8 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_9
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_9 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_10
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_10 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_11
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_11 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_12
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_12 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_13
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_13 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_14
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_14 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_15
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_15 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_16
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_16 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_17
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_17 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_18
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_18 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_19
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_19 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_20
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_20 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_21
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_21 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_22
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_22 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_23
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_23 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_24
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_24 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_25
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_25 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_26
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_26 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_27
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_27 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_28
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_28 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_29
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_29 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_30
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_30 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_31
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_31 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_32
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/rbl_br rbl_bl_1_1 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_32
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_33 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_33
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_34 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_34
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_35 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_35
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_36 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_36
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_37 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_37
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_38 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_38
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_39 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_39
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_40 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_40
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_41 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_41
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_42 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_42
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_43 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_43
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_44 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_44
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_45 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_45
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_46 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_46
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_47 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_47
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_48 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_48
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_49 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_49
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_50 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_50
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_51 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_51
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_52 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_52
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_53 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_53
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_54 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_54
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_55 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_55
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_56 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_56
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_57 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_57
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_58 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_58
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_59 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_59
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_60 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_60
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_61 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_61
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_62 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_62
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_63 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_63
+ vdd_uq1208 vdd_uq1241 vdd_uq1242 vdd_uq1243 vdd_uq1245 vdd_uq1246 vdd_uq1247 vdd_uq1248
+ vdd_uq1249 vdd_uq1250 vdd_uq1251 vdd_uq1252 vdd_uq1253 vdd_uq1254 vdd_uq1255 vdd_uq1256
+ vdd_uq1257 vdd_uq1258 vdd_uq1259 vdd_uq1260 vdd_uq1261 vdd_uq1262 vdd_uq1263 vdd_uq1264
+ vdd_uq1265 vdd_uq1266 vdd_uq1267 vdd_uq1268 vdd_uq1269 vdd_uq1270 vdd_uq1271 vdd_uq1272
+ vdd_uq1240 s_en1 p_en_bar1 vdd_uq1244 gnd sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_replica_bitcell_array_0 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_113
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_114 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_114
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_115 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_116
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_116 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_117
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_118 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_119
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_122 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_123
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_125 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_125
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_126 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_127
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/rbl_wl sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_96
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_98 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_101
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_103 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_104
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_105 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_106
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_107 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_107
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_108 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_109
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_110 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_83
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_84 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_85
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_86 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_72
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_87 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_89
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_64 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_91
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_92 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_73
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_74 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_65
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_93 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_94
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_95 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_75
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_69 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_77
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_66 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_78
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_80 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_70
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_81 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_67
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_71 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_82
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_31 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_32
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_34 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_36
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_37 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_37
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_38 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_38
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_39 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_40
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_41 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_42
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_43 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_44
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_45 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_46
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_47 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_48
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_49 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_49
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_50 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_51
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_52 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_53
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_55 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_56
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_58 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_59
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_59 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_60
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_61 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_62
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_63 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_30 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_2 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_13
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_26 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_2
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_14 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_3
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_3 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_15
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_26 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_4
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_16 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_16
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_17 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_17
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_28 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_18
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_28 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_29
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_19 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_19
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/rbl_wl sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_27
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_8 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_20
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_9 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_10 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_22
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_11 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_23
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_25 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_15
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_16 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_16
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_16 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_17
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_17 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_17
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_18 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_18
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_18 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_19
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_19 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_19
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_20 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_20
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_21 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_21
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_22 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_22
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_23 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_23
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_23 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_24
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_24 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_24
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_25 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_25
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_25 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_26
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_26 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_26
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_27 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_27
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_27 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_28
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_28 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_28
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_29 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_29
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_29 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_30
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_30 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_31
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_31 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_12
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_12 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_13
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_13 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_13
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_14 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_14
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_14 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/rbl_br
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_15 sky130_sram_1kbyte_1rw1r_32x256_8_replica_bitcell_array_0/rbl_br_1_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_15 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_0 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_1 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_1 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_2
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_2 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_2
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_3 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_3
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_3 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_4
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_4 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_4
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_5 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_10
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_10 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_11
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_11 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_12
+ rbl_bl_0_0 sky130_sram_1kbyte_1rw1r_32x256_8_replica_bitcell_array_0/rbl_bl_1_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_48 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_48
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_49 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_49
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_49 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_50
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_51 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_51
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_52 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_52
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_53 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_53
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_54 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_54
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_55 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_55
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_56 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_56
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_56 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_57
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_57 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_57
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_58 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_58
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_58 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_59
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_59 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_59
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_60 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_61
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_62 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_62
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_63 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_63
+ sky130_sram_1kbyte_1rw1r_32x256_8_replica_bitcell_array_0/rbl_bl_0_1 sky130_sram_1kbyte_1rw1r_32x256_8_replica_bitcell_array_0/rbl_br_0_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_34 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_34
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_34 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_35
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_35 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_35
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_46 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_48
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_36 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_36
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_36 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_37
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_46 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_37
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_37 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_38
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_38 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_32
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_38 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_32
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_46 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_39
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_39 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_39
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_47 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_47
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_40 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_40
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_41 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_41
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_33 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_47
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_42 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_42
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_43 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_33
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_43 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_44
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_44 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_45
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_45 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_45
+ gnd_uq194 gnd_uq1132 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_3 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_2
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_1 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_0 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_19
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_29 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_18
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_39 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_17
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_28 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_113
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_102 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_124
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_36 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_58
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_47 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_25
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_14 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_38
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_49 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_27
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_16 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_119
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_123 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_112
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_101 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_68
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_57 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_46
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_35 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_24
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_13 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_59
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_48 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_15
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_26 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_37
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_122 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_111
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_100 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_78
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_67 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_56
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_45 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_34
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_23 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_12
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_47 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_58
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_36 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_14
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_25 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_121
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_110 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_99
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_88 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_77
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_66 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_55
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_44 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_33
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_22 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_11
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_57 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_46
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_24 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_35
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_13 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_104
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_120 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_98
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_87 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_54
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_76 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_65
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_43 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_32
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_21 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_10
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_56 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_45
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_23 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_34
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_12 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_90
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_97 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_86
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_75 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_64
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_20 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_53
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_42 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_31
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_44 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_33
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_55 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_11
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_22 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_96
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_74 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_63
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_85 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_30
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_52 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_41
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_32 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_54
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_43 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_21
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_10 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_95
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_84 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_73
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_62 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_51
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_40 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_53
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_42 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_20
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_31 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_94
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_83 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_72
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_50 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_61
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_41 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_52
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_63 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_30
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_115 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_106
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_61 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_50
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_93 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_82
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_71 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_60
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_51 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_62
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_40 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_55
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_33 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_22
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_44 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_11
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_60 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_92
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_81 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_70
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_50 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_61
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_54 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_21
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_43 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_32
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_10 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_5
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_91 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_69
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_80 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_60
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_53 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_31
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_42 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_20
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_118 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_109
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_100 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_90
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_79 rbl_bl_1_1 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_63
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_52 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_41
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_30 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_89
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_127 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_7
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_62 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_51
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_40 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_121
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_112 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_61
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_50 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_103
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_60 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_124
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/rbl_br sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_18
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_9 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_57
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_48 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_39
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_105 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_21
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_12 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_33
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_4 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_117
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_108 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_99
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_9 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_9
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_8 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_9
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_24 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_76
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_15 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_8
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_126 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_6
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_54 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_8
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_9 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_7
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_8 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_120
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_7 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_111
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_102 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_7
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_8 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_6
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_7 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_6
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_6 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_7
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_5 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_35
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_68 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_6
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_88 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_27
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_79 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_97
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0/wl_29 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/br_5
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_5 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0/bl_6
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/br_4 sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0/bl_5
+ gnd vdd_uq259 sky130_sram_1kbyte_1rw1r_32x256_8_replica_bitcell_array
Xsky130_sram_1kbyte_1rw1r_32x256_8_port_address_0 wl_en0 addr0_1 addr0_2 addr0_3 addr0_4
+ addr0_5 addr0_6 addr0_7 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_64 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_65
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_66 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_67
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_68 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_69
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_70 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_71
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_72 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_73
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_74 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_75
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_76 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_77
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_78 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_79
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_80 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_81
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_82 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_83
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_84 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_85
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_86 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_87
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_88 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_89
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_90 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_91
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_92 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_93
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_94 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_95
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_96 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_97
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_98 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_99
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_100 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_101
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_102 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_103
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_104 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_105
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_106 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_107
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_108 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_109
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_110 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_111
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_112 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_113
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_114 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_115
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_116 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_117
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_118 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_119
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_120 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_121
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_122 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_123
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_124 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_125
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_126 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_127
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/rbl_wl sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_2 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_3
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_4 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_5
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_6 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_7
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_8 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_9
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_10 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_11
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_12 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_13
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_14 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_15
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_16 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_17
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_18 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_19
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_20 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_21
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_22 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_23
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_24 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_25
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_26 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_27
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_28 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_29
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_30 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_31
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_32 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_33
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_34 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_35
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_36 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_37
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_38 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_39
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_40 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_41
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_42 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_43
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_44 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_45
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_46 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_47
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_48 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_49
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_50 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_51
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_52 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_53
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_54 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_55
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_56 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_57
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_58 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_59
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_60 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_61
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_62 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_63
+ sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/wl_0 vdd_uq289 vdd_uq290 vdd_uq422
+ vdd_uq420 vdd_uq994 vdd_uq996 vdd_uq693 vdd_uq262 gnd_uq225 gnd_uq226 gnd_uq208
+ gnd_uq260 gnd_uq278 sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/gnd_uq26 vdd_uq336
+ vdd_uq320 vdd_uq368 vdd_uq274 gnd_uq312 vdd_uq335 gnd vdd_uq692 sky130_sram_1kbyte_1rw1r_32x256_8_port_address
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6 Z gnd vdd A VSUBS
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_360_sli_dli_da_p_0 gnd Z A gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_360_sli_dli_da_p
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli_da_p_0 vdd Z A vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli_da_p
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m4_w1_260_sli_dli_da_p S D G S_uq0
+ S_uq1 VSUBS
X0 S_uq0 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X1 D G S_uq1 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X2 D G S VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X3 S G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m4_w2_000_sli_dli_da_p S D G S_uq0
+ S_uq1 w_n59_116#
X0 D G S_uq1 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 D G S w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 S G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 S_uq0 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pinv_17 A Z gnd vdd
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m4_w1_260_sli_dli_da_p_0 gnd Z A gnd gnd gnd
+ sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m4_w1_260_sli_dli_da_p
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m4_w2_000_sli_dli_da_p_0 vdd Z A vdd vdd vdd
+ sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m4_w2_000_sli_dli_da_p
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pinv_11 A Z gnd vdd VSUBS
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m2_w0_740_sli_dli_da_p_0 gnd Z A gnd gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m2_w0_740_sli_dli_da_p
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m2_w1_260_sli_dli_da_p_0 vdd Z A vdd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m2_w1_260_sli_dli_da_p
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m12_w2_000_sli_dli_da_p S D G S_uq0
+ S_uq1 S_uq2 S_uq3 S_uq4 S_uq5 VSUBS
X0 S_uq3 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 S_uq2 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 D G S_uq5 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 S_uq0 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4 D G S_uq4 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 D G S_uq1 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 S_uq4 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7 D G S VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 S_uq1 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9 S G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10 D G S_uq3 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11 D G S_uq2 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m12_w2_000_sli_dli_da_p S D G S_uq0
+ S_uq1 S_uq2 S_uq3 S_uq4 S_uq5 w_n59_116#
X0 D G S_uq5 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 S_uq0 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 D G S_uq4 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 D G S_uq1 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4 S_uq4 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 D G S w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 S_uq1 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7 S G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 D G S_uq3 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9 D G S_uq2 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10 S_uq3 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11 S_uq2 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pinv_18 A Z vdd gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m12_w2_000_sli_dli_da_p_0 gnd Z A gnd gnd
+ gnd gnd gnd gnd gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m12_w2_000_sli_dli_da_p
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m12_w2_000_sli_dli_da_p_0 vdd Z A vdd vdd
+ vdd vdd vdd vdd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m12_w2_000_sli_dli_da_p
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pdriver_5 Z A gnd vdd
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_6_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6_0/Z
+ gnd vdd A sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6_0/VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_17_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_17_0/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_18_0/A gnd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_17
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_11_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6_0/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_17_0/A gnd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_11_0/VSUBS
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_11
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_18_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_18_0/A
+ Z vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_18
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19 A Z gnd vdd
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_360_sli_dli_da_p_0 gnd Z A gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_360_sli_dli_da_p
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli_da_p_0 vdd Z A vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli_da_p
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_delay_chain in out vdd vdd_uq6 vdd_uq2 vdd_uq8
+ vdd_uq4 gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_25 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_38/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_33/A gnd vdd_uq6 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_36 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_38/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_36/Z gnd vdd_uq6 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_14 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_9/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_14/Z gnd vdd_uq2 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_26 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_33/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_26/Z gnd vdd_uq6 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_37 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_38/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_37/Z gnd vdd_uq6 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_15 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_9/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_15/Z gnd vdd_uq2 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_27 out sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_27/Z
+ gnd vdd_uq8 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_38 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_39/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_38/Z gnd vdd_uq6 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_16 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_9/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_16/Z gnd vdd_uq2 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_28 out sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_28/Z
+ gnd vdd_uq8 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_39 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_39/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_39/Z gnd vdd_uq4 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_17 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_9/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_17/Z gnd vdd_uq2 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_29 out sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_29/Z
+ gnd vdd_uq8 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_18 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_7/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_9/A gnd vdd_uq2 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_19 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_7/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_19/Z gnd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_7/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_0/Z gnd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_1 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_7/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_1/Z gnd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_2 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_7/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_2/Z gnd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_3 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_7/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_3/Z gnd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_4 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_7/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_4/Z gnd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_5 in sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_7/A
+ gnd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_6 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_7/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_6/Z gnd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_7 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_7/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_7/Z gnd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_8 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_9/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_8/Z gnd vdd_uq2 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_9 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_9/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_9/Z gnd vdd_uq2 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_40 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_44/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_40/Z gnd vdd_uq4 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_30 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_33/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_30/Z gnd vdd_uq6 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_41 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_44/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_41/Z gnd vdd_uq4 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_31 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_33/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_31/Z gnd vdd_uq6 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_20 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_39/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_20/Z gnd vdd_uq4 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_42 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_44/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_42/Z gnd vdd_uq4 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_32 out sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_32/Z
+ gnd vdd_uq8 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_21 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_39/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_21/Z gnd vdd_uq4 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_43 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_44/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_43/Z gnd vdd_uq4 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_10 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_9/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_10/Z gnd vdd_uq2 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_33 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_33/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_33/Z gnd vdd_uq6 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_34 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_38/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_34/Z gnd vdd_uq6 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_22 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_39/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_22/Z gnd vdd_uq4 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_23 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_44/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_39/A gnd vdd_uq4 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_44 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_9/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_44/Z gnd vdd_uq4 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_11 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_9/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_11/Z gnd vdd_uq2 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_12 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_7/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_12/Z gnd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_24 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_33/A
+ out gnd vdd_uq8 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_35 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_38/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_35/Z gnd vdd_uq6 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_13 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_9/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19_13/Z gnd vdd_uq2 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_19
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pnand2_1 Z vdd A B gnd VSUBS
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sli_dactive_0 gnd A sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sactive_dli_0/a_0_0#
+ sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sli_dactive_0/w_n26_n26# gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sli_dactive
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sactive_dli_0 Z B sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sactive_dli_0/w_n26_n26#
+ sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sactive_dli_0/a_0_0# gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sactive_dli
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli_0 Z vdd B vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli_1 vdd Z A vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m18_w2_000_sli_dli_da_p S D G S_uq0
+ S_uq1 S_uq2 S_uq3 S_uq4 S_uq5 S_uq6 S_uq7 S_uq8 w_n59_116#
X0 D G S_uq8 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 S_uq2 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 D G S_uq7 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 S G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4 D G S_uq4 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 S_uq7 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 D G S_uq3 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7 D G S_uq1 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 S_uq4 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9 S_uq1 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10 S_uq0 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11 S_uq3 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12 D G S_uq6 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13 D G S_uq5 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14 D G S_uq2 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15 D G S w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X16 S_uq6 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X17 S_uq5 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m18_w2_000_sli_dli_da_p S D G S_uq0
+ S_uq1 S_uq2 S_uq3 S_uq4 S_uq5 S_uq6 S_uq7 S_uq8 VSUBS
X0 S_uq6 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 S_uq5 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 D G S_uq8 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 S_uq2 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4 D G S_uq7 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 S G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 D G S_uq4 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7 S_uq7 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 D G S_uq3 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9 D G S_uq1 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10 S_uq4 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11 S_uq1 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12 S_uq0 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13 S_uq3 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14 D G S_uq6 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15 D G S_uq5 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X16 D G S_uq2 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X17 D G S VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pinv_16 A Z gnd vdd
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m18_w2_000_sli_dli_da_p_0 vdd Z A vdd vdd
+ vdd vdd vdd vdd vdd vdd vdd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m18_w2_000_sli_dli_da_p
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m18_w2_000_sli_dli_da_p_0 gnd Z A gnd gnd
+ gnd gnd gnd gnd gnd gnd gnd gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m18_w2_000_sli_dli_da_p
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pdriver_4 Z A vdd gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_16_0 A Z gnd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_16
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pnand3 A B C Z gnd vdd w_n36_679# VSUBS
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sli_dactive_0 gnd A a_154_51# sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sli_dactive_0/w_n26_n26#
+ VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sli_dactive
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sactive_dli_0 Z C sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sli_dactive_0/w_n26_n26#
+ a_244_51# VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sactive_dli
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli_0 vdd Z C w_n36_679# sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli_1 Z vdd B w_n36_679# sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli_2 vdd Z A w_n36_679# sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli
X0 a_244_51# B a_154_51# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pand3_0 Z A B C vdd gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_pdriver_4_0 Z sky130_sram_1kbyte_1rw1r_32x256_8_pnand3_0/Z
+ vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pdriver_4
Xsky130_sram_1kbyte_1rw1r_32x256_8_pnand3_0 A B C sky130_sram_1kbyte_1rw1r_32x256_8_pnand3_0/Z
+ gnd vdd vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pnand3
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m5_w2_000_sli_dli_da_p S D G S_uq0
+ S_uq1 w_n59_116#
X0 D G S_uq1 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 D G S w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 S G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 D G S_uq0 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4 S_uq0 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m5_w1_680_sli_dli_da_p S D G S_uq0
+ S_uq1 VSUBS
X0 S_uq0 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X1 D G S_uq1 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X2 D G S VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X3 S G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X4 D G S_uq0 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pinv_8 A Z vdd gnd VSUBS
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m5_w2_000_sli_dli_da_p_0 vdd Z A vdd vdd vdd
+ sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m5_w2_000_sli_dli_da_p
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m5_w1_680_sli_dli_da_p_0 gnd Z A gnd gnd gnd
+ sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m5_w1_680_sli_dli_da_p
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m13_w2_000_sli_dli_da_p S D G S_uq0
+ S_uq1 S_uq2 S_uq3 S_uq4 S_uq5 w_n59_116#
X0 D G S_uq5 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 S_uq0 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 D G S_uq4 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 D G S_uq1 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4 S_uq4 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 D G S w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 S_uq1 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7 S G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 D G S_uq3 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9 D G S_uq2 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10 D G S_uq0 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11 S_uq3 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12 S_uq2 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m13_w2_000_sli_dli_da_p S D G S_uq0
+ S_uq1 S_uq2 S_uq3 S_uq4 S_uq5 VSUBS
X0 S_uq3 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 S_uq2 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 D G S_uq5 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 S_uq0 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4 D G S_uq4 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 D G S_uq1 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 S_uq4 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7 D G S VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 S_uq1 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9 S G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10 D G S_uq3 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11 D G S_uq2 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12 D G S_uq0 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pinv_9 A Z vdd gnd VSUBS
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m13_w2_000_sli_dli_da_p_0 vdd Z A vdd vdd
+ vdd vdd vdd vdd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m13_w2_000_sli_dli_da_p
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m13_w2_000_sli_dli_da_p_0 gnd Z A gnd gnd
+ gnd gnd gnd gnd gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m13_w2_000_sli_dli_da_p
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m39_w2_000_sli_dli_da_p S D G S_uq0
+ S_uq1 S_uq2 S_uq3 S_uq4 S_uq5 S_uq6 S_uq7 S_uq8 S_uq9 S_uq10 S_uq11 S_uq12 S_uq13
+ S_uq14 S_uq15 S_uq16 S_uq17 S_uq18 w_n59_116#
X0 S_uq7 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 S_uq3 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 S_uq2 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 D G S_uq18 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4 S_uq12 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 S G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 D G S_uq17 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7 S_uq10 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 S_uq5 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9 D G S_uq14 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10 D G S_uq4 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11 D G S_uq0 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12 D G S_uq6 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13 D G S_uq3 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14 D G S_uq1 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15 S_uq17 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X16 D G S_uq13 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X17 D G S_uq11 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X18 D G S_uq8 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X19 S_uq14 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X20 S_uq0 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X21 S_uq11 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X22 S_uq9 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X23 S_uq8 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X24 S_uq6 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X25 S_uq4 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X26 S_uq1 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X27 S_uq13 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X28 D G S_uq16 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X29 D G S_uq15 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X30 D G S_uq5 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X31 D G S w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X32 D G S_uq12 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X33 D G S_uq10 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X34 D G S_uq9 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X35 D G S_uq7 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X36 D G S_uq2 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X37 S_uq16 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X38 S_uq15 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m39_w2_000_sli_dli_da_p S D G S_uq0
+ S_uq1 S_uq2 S_uq3 S_uq4 S_uq5 S_uq6 S_uq7 S_uq8 S_uq9 S_uq10 S_uq11 S_uq12 S_uq13
+ S_uq14 S_uq15 S_uq16 S_uq17 S_uq18 VSUBS
X0 S_uq16 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 S_uq15 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 S_uq3 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 S_uq2 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4 D G S_uq18 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 S_uq12 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 S_uq7 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7 D G S_uq17 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 S_uq10 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9 S_uq5 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10 S G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11 D G S_uq14 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12 D G S_uq4 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13 D G S_uq0 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14 D G S_uq1 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15 S_uq17 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X16 D G S_uq13 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X17 D G S_uq11 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X18 D G S_uq8 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X19 D G S_uq6 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X20 D G S_uq3 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X21 S_uq14 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X22 S_uq0 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X23 S_uq11 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X24 S_uq9 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X25 S_uq6 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X26 S_uq4 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X27 S_uq1 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X28 S_uq13 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X29 S_uq8 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X30 D G S_uq16 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X31 D G S_uq15 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X32 D G S VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X33 D G S_uq12 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X34 D G S_uq10 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X35 D G S_uq9 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X36 D G S_uq7 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X37 D G S_uq5 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X38 D G S_uq2 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pinv_20 A Z vdd gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m39_w2_000_sli_dli_da_p_0 vdd Z A vdd vdd
+ vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m39_w2_000_sli_dli_da_p
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m39_w2_000_sli_dli_da_p_0 gnd Z A gnd gnd
+ gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m39_w2_000_sli_dli_da_p
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m2_w1_260_sli_dli_da_p S D G S_uq0
+ VSUBS
X0 D G S VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X1 S_uq0 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m2_w2_000_sli_dli_da_p S D G S_uq0
+ w_n59_116#
X0 D G S w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 S_uq0 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pinv_7 A Z gnd vdd VSUBS
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m2_w1_260_sli_dli_da_p_0 gnd Z A gnd gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m2_w1_260_sli_dli_da_p
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m2_w2_000_sli_dli_da_p_0 vdd Z A vdd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m2_w2_000_sli_dli_da_p
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pdriver_6 Z A vdd gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_8_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_8_0/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_9_0/A vdd gnd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_8
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_6_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_7_0/A
+ gnd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6_1/Z gnd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_6_1 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6_1/Z
+ gnd vdd A gnd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_9_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_9_0/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_9_0/Z vdd gnd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_9
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_20_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_9_0/Z
+ Z vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_20
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_7_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_7_0/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_8_0/A gnd vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_7
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_dff_buf_0 clk Q Qb vdd D gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_2_0 Qb Q gnd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_2_0/VSUBS
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_2
Xsky130_fd_bd_sram__openram_dff_0 sky130_fd_bd_sram__openram_dff_0/QN D sky130_fd_bd_sram__openram_dff_0/Q
+ clk vdd gnd gnd sky130_fd_bd_sram__openram_dff
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_1_0 sky130_fd_bd_sram__openram_dff_0/Q Qb
+ gnd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_1_0/VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_pinv_1
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_dff_buf_array_0 din_0 dout_0 dout_bar_0
+ clk vdd gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_dff_buf_0_0 clk dout_0 dout_bar_0 vdd din_0 gnd
+ sky130_sram_1kbyte_1rw1r_32x256_8_dff_buf_0
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m24_w2_000_sli_dli_da_p S D G S_uq0
+ S_uq1 S_uq2 S_uq3 S_uq4 S_uq5 S_uq6 S_uq7 S_uq8 S_uq9 S_uq10 S_uq11 VSUBS
X0 S_uq9 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 S_uq8 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 D G S_uq11 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 S_uq5 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4 S G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 D G S_uq10 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 S_uq3 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7 D G S_uq7 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 S_uq10 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9 D G S_uq6 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10 D G S_uq4 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11 D G S_uq1 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12 S_uq7 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13 S_uq4 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14 S_uq2 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15 S_uq0 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X16 S_uq6 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X17 S_uq1 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X18 D G S_uq9 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X19 D G S_uq8 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X20 D G S_uq5 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X21 D G S_uq3 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X22 D G S_uq2 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X23 D G S VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m24_w2_000_sli_dli_da_p S D G S_uq0
+ S_uq1 S_uq2 S_uq3 S_uq4 S_uq5 S_uq6 S_uq7 S_uq8 S_uq9 S_uq10 S_uq11 w_n59_116#
X0 S G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 D G S_uq11 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 S_uq5 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 D G S_uq10 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4 S_uq3 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 D G S_uq7 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 S_uq10 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7 D G S_uq6 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 D G S_uq4 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9 D G S_uq1 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10 S_uq7 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11 S_uq4 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12 S_uq2 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13 S_uq1 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14 S_uq0 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15 S_uq6 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X16 D G S_uq9 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X17 D G S_uq8 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X18 D G S_uq5 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X19 D G S_uq3 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X20 D G S_uq2 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X21 D G S w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X22 S_uq9 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X23 S_uq8 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pinv_14 A Z vdd gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m24_w2_000_sli_dli_da_p_0 gnd Z A gnd gnd
+ gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m24_w2_000_sli_dli_da_p
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m24_w2_000_sli_dli_da_p_0 vdd Z A vdd vdd
+ vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m24_w2_000_sli_dli_da_p
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m3_w2_000_sli_dli_da_p S D G S_uq0
+ VSUBS
X0 D G S VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 D G S_uq0 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 S_uq0 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m3_w2_000_sli_dli_da_p S D G S_uq0
+ w_n59_116#
X0 D G S w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 D G S_uq0 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 S_uq0 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pinv_12 A Z vdd gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m3_w2_000_sli_dli_da_p_0 gnd Z A gnd gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m3_w2_000_sli_dli_da_p
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m3_w2_000_sli_dli_da_p_0 vdd Z A vdd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m3_w2_000_sli_dli_da_p
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m8_w2_000_sli_dli_da_p S D G S_uq0
+ S_uq1 S_uq2 S_uq3 VSUBS
X0 S_uq1 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 S G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 D G S_uq3 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 D G S_uq2 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4 S_uq2 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 S_uq0 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 D G S_uq1 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7 D G S VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m8_w2_000_sli_dli_da_p S D G S_uq0
+ S_uq1 S_uq2 S_uq3 w_n59_116#
X0 D G S_uq3 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 D G S_uq2 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 S_uq2 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 S_uq0 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4 D G S_uq1 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 D G S w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 S_uq1 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7 S G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pinv_13 A Z vdd gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m8_w2_000_sli_dli_da_p_0 gnd Z A gnd gnd gnd
+ gnd gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m8_w2_000_sli_dli_da_p
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m8_w2_000_sli_dli_da_p_0 vdd Z A vdd vdd vdd
+ vdd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m8_w2_000_sli_dli_da_p
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pdriver_2 Z A vdd gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_14_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_14_0/A
+ Z vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_14
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_12_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_12_0/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_13_0/A vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_12
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_6_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6_0/Z
+ gnd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6_1/Z gnd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_6_1 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6_1/Z
+ gnd vdd A gnd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_13_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_13_0/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_14_0/A vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_13
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_11_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6_0/Z
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_12_0/A gnd vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_11
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m7_w1_680_sli_dli_da_p S D G S_uq0
+ S_uq1 S_uq2 VSUBS
X0 S G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X1 S_uq0 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X2 D G S_uq2 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X3 D G S_uq1 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X4 S_uq1 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X5 D G S VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X6 D G S_uq0 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m7_w2_000_sli_dli_da_p S D G S_uq0
+ S_uq1 S_uq2 w_n59_116#
X0 D G S_uq2 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 D G S_uq1 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 S_uq1 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 D G S w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4 D G S_uq0 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 S G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 S_uq0 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pinv_3 A Z gnd vdd
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m7_w1_680_sli_dli_da_p_0 gnd Z A gnd gnd gnd
+ gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m7_w1_680_sli_dli_da_p
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m7_w2_000_sli_dli_da_p_0 vdd Z A vdd vdd vdd
+ vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m7_w2_000_sli_dli_da_p
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pdriver_0 Z A vdd gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_3_0 A Z gnd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_3
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pnand2_0 Z gnd vdd A B w_n36_679# VSUBS
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sli_dactive_0 gnd A sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sactive_dli_0/a_0_0#
+ sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sli_dactive_0/w_n26_n26# VSUBS
+ sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sli_dactive
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sactive_dli_0 Z B sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sli_dactive_0/w_n26_n26#
+ sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sactive_dli_0/a_0_0# VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m1_w0_740_sactive_dli
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli_0 Z vdd B w_n36_679# sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli_1 vdd Z A w_n36_679# sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m1_w1_120_sli_dli
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pand2_0 Z A B vdd gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_pdriver_0_0 Z sky130_sram_1kbyte_1rw1r_32x256_8_pnand2_0_0/Z
+ vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pdriver_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_pnand2_0_0 sky130_sram_1kbyte_1rw1r_32x256_8_pnand2_0_0/Z
+ gnd vdd A B vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pnand2_0
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_control_logic_r csb wl_en s_en rbl_bl p_en_bar
+ clk clk_buf vdd_uq0 vdd vdd_uq3 vdd_uq9 vdd_uq11 vdd_uq12 vdd_uq7 vdd_uq5 gnd vdd_uq10
Xsky130_sram_1kbyte_1rw1r_32x256_8_pdriver_5_0 p_en_bar sky130_sram_1kbyte_1rw1r_32x256_8_pnand2_1_0/Z
+ gnd vdd_uq12 sky130_sram_1kbyte_1rw1r_32x256_8_pdriver_5
Xsky130_sram_1kbyte_1rw1r_32x256_8_delay_chain_0 rbl_bl sky130_sram_1kbyte_1rw1r_32x256_8_pand3_0_0/A
+ vdd_uq9 vdd_uq3 vdd_uq7 vdd vdd_uq5 gnd sky130_sram_1kbyte_1rw1r_32x256_8_delay_chain
Xsky130_sram_1kbyte_1rw1r_32x256_8_pnand2_1_0 sky130_sram_1kbyte_1rw1r_32x256_8_pnand2_1_0/Z
+ vdd_uq12 sky130_sram_1kbyte_1rw1r_32x256_8_pand2_0_0/Z sky130_sram_1kbyte_1rw1r_32x256_8_pand3_0_0/A
+ gnd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pnand2_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_0_0 clk_buf sky130_sram_1kbyte_1rw1r_32x256_8_pinv_0_0/Z
+ gnd vdd_uq10 gnd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_pand3_0_0 s_en sky130_sram_1kbyte_1rw1r_32x256_8_pand3_0_0/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pand3_0_0/B sky130_sram_1kbyte_1rw1r_32x256_8_pand3_0_0/C
+ vdd_uq11 gnd sky130_sram_1kbyte_1rw1r_32x256_8_pand3_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_pdriver_6_0 clk_buf clk vdd_uq10 gnd sky130_sram_1kbyte_1rw1r_32x256_8_pdriver_6
Xsky130_sram_1kbyte_1rw1r_32x256_8_dff_buf_array_0_0 csb sky130_sram_1kbyte_1rw1r_32x256_8_dff_buf_array_0_0/dout_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_pand3_0_0/C clk_buf vdd_uq0 gnd sky130_sram_1kbyte_1rw1r_32x256_8_dff_buf_array_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_pdriver_2_0 wl_en sky130_sram_1kbyte_1rw1r_32x256_8_pand3_0_0/B
+ vdd_uq12 gnd sky130_sram_1kbyte_1rw1r_32x256_8_pdriver_2
Xsky130_sram_1kbyte_1rw1r_32x256_8_pand2_0_0 sky130_sram_1kbyte_1rw1r_32x256_8_pand2_0_0/Z
+ clk_buf sky130_sram_1kbyte_1rw1r_32x256_8_pand3_0_0/C vdd_uq11 gnd sky130_sram_1kbyte_1rw1r_32x256_8_pand2_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_pand2_0_1 sky130_sram_1kbyte_1rw1r_32x256_8_pand3_0_0/B
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_0_0/Z sky130_sram_1kbyte_1rw1r_32x256_8_pand3_0_0/C
+ vdd_uq10 gnd sky130_sram_1kbyte_1rw1r_32x256_8_pand2_0
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m40_w2_000_sli_dli_da_p S D G S_uq0
+ S_uq1 S_uq2 S_uq3 S_uq4 S_uq5 S_uq6 S_uq7 S_uq8 S_uq9 S_uq10 S_uq11 S_uq12 S_uq13
+ S_uq14 S_uq15 S_uq16 S_uq17 S_uq18 S_uq19 w_n59_116#
X0 S_uq8 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 S_uq4 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 S_uq3 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 S_uq0 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4 D G S_uq19 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 S_uq13 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 S_uq1 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7 D G S_uq18 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 S_uq11 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9 S_uq6 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10 D G S_uq15 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11 D G S_uq5 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12 D G S w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13 D G S_uq7 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14 D G S_uq4 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15 D G S_uq2 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X16 S_uq18 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X17 D G S_uq14 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X18 D G S_uq12 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X19 D G S_uq9 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X20 S_uq15 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X21 S G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X22 S_uq12 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X23 S_uq10 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X24 S_uq9 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X25 S_uq7 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X26 S_uq5 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X27 S_uq2 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X28 S_uq14 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X29 D G S_uq17 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X30 D G S_uq16 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X31 D G S_uq6 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X32 D G S_uq1 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X33 D G S_uq13 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X34 D G S_uq11 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X35 D G S_uq10 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X36 D G S_uq8 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X37 D G S_uq3 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X38 S_uq17 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X39 S_uq16 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m40_w2_000_sli_dli_da_p S D G S_uq0
+ S_uq1 S_uq2 S_uq3 S_uq4 S_uq5 S_uq6 S_uq7 S_uq8 S_uq9 S_uq10 S_uq11 S_uq12 S_uq13
+ S_uq14 S_uq15 S_uq16 S_uq17 S_uq18 S_uq19 VSUBS
X0 S_uq17 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 S_uq16 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 S_uq4 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 S_uq3 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4 S_uq0 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 D G S_uq19 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 S_uq13 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7 S_uq8 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 D G S_uq18 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9 S_uq11 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10 S_uq6 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11 S_uq1 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12 D G S_uq15 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13 D G S_uq5 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14 D G S VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15 D G S_uq2 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X16 S_uq18 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X17 D G S_uq14 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X18 D G S_uq12 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X19 D G S_uq9 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X20 D G S_uq7 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X21 D G S_uq4 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X22 S_uq15 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X23 S G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X24 S_uq12 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X25 S_uq10 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X26 S_uq7 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X27 S_uq5 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X28 S_uq2 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X29 S_uq14 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X30 S_uq9 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X31 D G S_uq17 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X32 D G S_uq16 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X33 D G S_uq1 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X34 D G S_uq13 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X35 D G S_uq11 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X36 D G S_uq10 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X37 D G S_uq8 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X38 D G S_uq6 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X39 D G S_uq3 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pinv_10 A Z vdd gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m40_w2_000_sli_dli_da_p_0 vdd Z A vdd vdd
+ vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m40_w2_000_sli_dli_da_p
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m40_w2_000_sli_dli_da_p_0 gnd Z A gnd gnd
+ gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m40_w2_000_sli_dli_da_p
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pdriver_1 Z vdd A gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_8_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_8_0/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_9_0/A vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_8_0/VSUBS
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_8
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_6_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_7_0/A
+ gnd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6_1/Z gnd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_6_1 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6_1/Z
+ gnd vdd A gnd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_10_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_9_0/Z
+ Z vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_10
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_9_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_9_0/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_9_0/Z vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_9_0/VSUBS
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_9
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_7_0 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_7_0/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_8_0/A gnd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_7_0/VSUBS
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_7
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m22_w2_000_sli_dli_da_p S D G S_uq0
+ S_uq1 S_uq2 S_uq3 S_uq4 S_uq5 S_uq6 S_uq7 S_uq8 S_uq9 S_uq10 VSUBS
X0 S_uq8 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 S_uq7 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 D G S_uq10 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 S_uq4 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4 S_uq0 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 D G S_uq9 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 S_uq2 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7 D G S_uq6 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 S_uq9 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9 D G S_uq5 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10 D G S_uq3 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11 D G S VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12 S_uq6 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13 S_uq3 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14 S_uq1 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15 S_uq5 G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X16 S G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X17 D G S_uq8 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X18 D G S_uq7 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X19 D G S_uq4 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X20 D G S_uq2 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X21 D G S_uq1 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m22_w2_000_sli_dli_da_p S D G S_uq0
+ S_uq1 S_uq2 S_uq3 S_uq4 S_uq5 S_uq6 S_uq7 S_uq8 S_uq9 S_uq10 w_n59_116#
X0 S_uq0 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 D G S_uq10 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 S_uq4 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 D G S_uq9 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4 S_uq2 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 D G S_uq6 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6 S_uq9 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7 D G S_uq5 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 D G S_uq3 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9 D G S w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10 S_uq6 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11 S_uq3 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12 S_uq1 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13 S G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14 S_uq5 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15 D G S_uq8 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X16 D G S_uq7 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X17 D G S_uq4 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X18 D G S_uq2 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X19 D G S_uq1 w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X20 S_uq8 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X21 S_uq7 G D w_n59_116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pinv_15 A Z vdd gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_nmos_m22_w2_000_sli_dli_da_p_0 gnd Z A gnd gnd
+ gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m22_w2_000_sli_dli_da_p
Xsky130_sram_1kbyte_1rw1r_32x256_8_pmos_m22_w2_000_sli_dli_da_p_0 vdd Z A vdd vdd
+ vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m22_w2_000_sli_dli_da_p
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pdriver_3 Z A vdd gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_15_0 A Z vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pinv_15
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_pand3 Z A B C vdd gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_pdriver_3_0 Z sky130_sram_1kbyte_1rw1r_32x256_8_pnand3_0/Z
+ vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pdriver_3
Xsky130_sram_1kbyte_1rw1r_32x256_8_pnand3_0 A B C sky130_sram_1kbyte_1rw1r_32x256_8_pnand3_0/Z
+ gnd vdd vdd gnd sky130_sram_1kbyte_1rw1r_32x256_8_pnand3
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_dff_buf_array dout_0 dout_bar_0 dout_1 dout_bar_1
+ clk din_0 din_1 gnd vdd
Xsky130_sram_1kbyte_1rw1r_32x256_8_dff_buf_0_0 clk dout_1 dout_bar_1 vdd din_1 gnd
+ sky130_sram_1kbyte_1rw1r_32x256_8_dff_buf_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_dff_buf_0_1 clk dout_0 dout_bar_0 vdd din_0 gnd
+ sky130_sram_1kbyte_1rw1r_32x256_8_dff_buf_0
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_control_logic_rw web wl_en w_en s_en rbl_bl
+ p_en_bar clk clk_buf vdd_uq0 vdd vdd_uq3 vdd_uq5 vdd_uq9 vdd_uq13 vdd_uq11 csb vdd_uq7
+ vdd_uq12 vdd_uq10 gnd
Xsky130_sram_1kbyte_1rw1r_32x256_8_pdriver_5_0 p_en_bar sky130_sram_1kbyte_1rw1r_32x256_8_pnand2_1_0/Z
+ gnd vdd_uq12 sky130_sram_1kbyte_1rw1r_32x256_8_pdriver_5
Xsky130_sram_1kbyte_1rw1r_32x256_8_pdriver_1_0 clk_buf vdd_uq10 clk gnd sky130_sram_1kbyte_1rw1r_32x256_8_pdriver_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_delay_chain_0 rbl_bl sky130_sram_1kbyte_1rw1r_32x256_8_pinv_0_1/A
+ vdd_uq9 vdd_uq3 vdd_uq7 vdd vdd_uq5 gnd sky130_sram_1kbyte_1rw1r_32x256_8_delay_chain
Xsky130_sram_1kbyte_1rw1r_32x256_8_pnand2_1_0 sky130_sram_1kbyte_1rw1r_32x256_8_pnand2_1_0/Z
+ vdd_uq12 sky130_sram_1kbyte_1rw1r_32x256_8_pand2_0_0/Z sky130_sram_1kbyte_1rw1r_32x256_8_pinv_0_1/A
+ gnd sky130_sram_1kbyte_1rw1r_32x256_8_pnand2_1_0/VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_pnand2_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_0_0 clk_buf sky130_sram_1kbyte_1rw1r_32x256_8_pinv_0_0/Z
+ gnd vdd_uq10 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_0_0/VSUBS sky130_sram_1kbyte_1rw1r_32x256_8_pinv_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_pinv_0_1 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_0_1/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pand3_0/B gnd vdd_uq13 sky130_sram_1kbyte_1rw1r_32x256_8_pinv_0_1/VSUBS
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_pand3_0_0 s_en sky130_sram_1kbyte_1rw1r_32x256_8_pinv_0_1/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pand3_0/C sky130_sram_1kbyte_1rw1r_32x256_8_pand3_0_0/C
+ vdd_uq11 gnd sky130_sram_1kbyte_1rw1r_32x256_8_pand3_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_pdriver_2_0 wl_en sky130_sram_1kbyte_1rw1r_32x256_8_pand3_0/C
+ vdd_uq13 gnd sky130_sram_1kbyte_1rw1r_32x256_8_pdriver_2
Xsky130_sram_1kbyte_1rw1r_32x256_8_pand3_0 w_en sky130_sram_1kbyte_1rw1r_32x256_8_pand3_0/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_pand3_0/B sky130_sram_1kbyte_1rw1r_32x256_8_pand3_0/C
+ vdd_uq12 gnd sky130_sram_1kbyte_1rw1r_32x256_8_pand3
Xsky130_sram_1kbyte_1rw1r_32x256_8_pand2_0_0 sky130_sram_1kbyte_1rw1r_32x256_8_pand2_0_0/Z
+ clk_buf sky130_sram_1kbyte_1rw1r_32x256_8_pand2_0_1/B vdd_uq11 gnd sky130_sram_1kbyte_1rw1r_32x256_8_pand2_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_pand2_0_1 sky130_sram_1kbyte_1rw1r_32x256_8_pand3_0/C
+ sky130_sram_1kbyte_1rw1r_32x256_8_pinv_0_0/Z sky130_sram_1kbyte_1rw1r_32x256_8_pand2_0_1/B
+ vdd_uq10 gnd sky130_sram_1kbyte_1rw1r_32x256_8_pand2_0
Xsky130_sram_1kbyte_1rw1r_32x256_8_dff_buf_array_0 sky130_sram_1kbyte_1rw1r_32x256_8_dff_buf_array_0/dout_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_pand2_0_1/B sky130_sram_1kbyte_1rw1r_32x256_8_pand3_0_0/C
+ sky130_sram_1kbyte_1rw1r_32x256_8_pand3_0/A clk_buf csb web gnd vdd_uq0 sky130_sram_1kbyte_1rw1r_32x256_8_dff_buf_array
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_col_addr_dff vdd gnd clk din_0 dout_0
Xsky130_fd_bd_sram__openram_dff_0 sky130_fd_bd_sram__openram_dff_0/QN din_0 dout_0
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_row_addr_dff vdd clk din_0 dout_0 din_1
+ dout_1 din_2 dout_2 din_3 dout_3 din_4 dout_4 din_5 dout_5 din_6 dout_6 vdd_uq0
+ vdd_uq1 vdd_uq2 gnd
Xsky130_fd_bd_sram__openram_dff_5 sky130_fd_bd_sram__openram_dff_5/QN din_1 dout_1
+ clk vdd_uq0 gnd sky130_fd_bd_sram__openram_dff_5/VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_6 sky130_fd_bd_sram__openram_dff_6/QN din_0 dout_0
+ clk vdd_uq0 gnd sky130_fd_bd_sram__openram_dff_6/VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_0 sky130_fd_bd_sram__openram_dff_0/QN din_6 dout_6
+ clk vdd_uq2 gnd sky130_fd_bd_sram__openram_dff_0/VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_1 sky130_fd_bd_sram__openram_dff_1/QN din_5 dout_5
+ clk vdd_uq1 gnd sky130_fd_bd_sram__openram_dff_1/VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_2 sky130_fd_bd_sram__openram_dff_2/QN din_4 dout_4
+ clk vdd_uq1 gnd sky130_fd_bd_sram__openram_dff_2/VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_4 sky130_fd_bd_sram__openram_dff_4/QN din_2 dout_2
+ clk vdd gnd sky130_fd_bd_sram__openram_dff_4/VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_3 sky130_fd_bd_sram__openram_dff_3/QN din_3 dout_3
+ clk vdd gnd sky130_fd_bd_sram__openram_dff_3/VSUBS sky130_fd_bd_sram__openram_dff
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8_data_dff clk din_0 din_1 dout_1 din_2 dout_2
+ din_3 dout_3 din_4 dout_4 din_5 dout_5 din_6 dout_6 din_7 dout_7 din_8 dout_8 din_9
+ dout_9 din_10 dout_10 din_11 dout_11 din_12 dout_12 din_13 dout_13 dout_14 din_15
+ dout_15 din_16 dout_16 din_17 dout_17 din_18 dout_18 din_19 dout_19 din_20 dout_20
+ din_21 dout_21 din_22 dout_22 din_23 dout_23 din_24 dout_24 din_25 dout_25 din_26
+ dout_26 din_27 dout_27 din_28 dout_28 din_29 dout_29 din_30 dout_30 din_31 dout_31
+ gnd vdd din_14 dout_0
Xsky130_fd_bd_sram__openram_dff_5 sky130_fd_bd_sram__openram_dff_5/QN din_6 dout_6
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_6 sky130_fd_bd_sram__openram_dff_6/QN din_5 dout_5
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_7 sky130_fd_bd_sram__openram_dff_7/QN din_14 dout_14
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_8 sky130_fd_bd_sram__openram_dff_8/QN din_13 dout_13
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_9 sky130_fd_bd_sram__openram_dff_9/QN din_12 dout_12
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_30 sky130_fd_bd_sram__openram_dff_30/QN din_16 dout_16
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_20 sky130_fd_bd_sram__openram_dff_20/QN din_22 dout_22
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_31 sky130_fd_bd_sram__openram_dff_31/QN din_15 dout_15
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_21 sky130_fd_bd_sram__openram_dff_21/QN din_31 dout_31
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_10 sky130_fd_bd_sram__openram_dff_10/QN din_11 dout_11
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_22 sky130_fd_bd_sram__openram_dff_22/QN din_30 dout_30
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_11 sky130_fd_bd_sram__openram_dff_11/QN din_10 dout_10
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_23 sky130_fd_bd_sram__openram_dff_23/QN din_29 dout_29
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_24 sky130_fd_bd_sram__openram_dff_24/QN din_28 dout_28
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_12 sky130_fd_bd_sram__openram_dff_12/QN din_9 dout_9
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_13 sky130_fd_bd_sram__openram_dff_13/QN din_8 dout_8
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_25 sky130_fd_bd_sram__openram_dff_25/QN din_27 dout_27
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_14 sky130_fd_bd_sram__openram_dff_14/QN din_7 dout_7
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_26 sky130_fd_bd_sram__openram_dff_26/QN din_26 dout_26
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_15 sky130_fd_bd_sram__openram_dff_15/QN din_21 dout_21
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_27 sky130_fd_bd_sram__openram_dff_27/QN din_25 dout_25
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_16 sky130_fd_bd_sram__openram_dff_16/QN din_20 dout_20
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_28 sky130_fd_bd_sram__openram_dff_28/QN din_24 dout_24
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_17 sky130_fd_bd_sram__openram_dff_17/QN din_19 dout_19
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_29 sky130_fd_bd_sram__openram_dff_29/QN din_23 dout_23
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_18 sky130_fd_bd_sram__openram_dff_18/QN din_18 dout_18
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_19 sky130_fd_bd_sram__openram_dff_19/QN din_17 dout_17
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_0 sky130_fd_bd_sram__openram_dff_0/QN din_2 dout_2
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_1 sky130_fd_bd_sram__openram_dff_1/QN din_4 dout_4
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_2 sky130_fd_bd_sram__openram_dff_2/QN din_3 dout_3
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_3 sky130_fd_bd_sram__openram_dff_3/QN din_1 dout_1
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_4 sky130_fd_bd_sram__openram_dff_4/QN din_0 dout_0
+ clk vdd gnd VSUBS sky130_fd_bd_sram__openram_dff
.ends

.subckt sky130_sram_1kbyte_1rw1r_32x256_8 csb0 web0 addr0[1] addr0[2] addr0[3] addr0[4]
+ addr0[5] addr0[6] addr0[7] csb1 addr1[1] addr1[2] addr1[3] vccd1 clk1 dout1[16]
+ dout1[17] dout1[18] dout1[19] dout1[20] dout1[21] dout1[22] dout1[23] dout1[24]
+ dout1[25] dout1[26] dout1[27] dout1[28] dout1[29] dout1[30] dout1[31] addr1[0] dout1[1]
+ dout1[2] dout1[3] dout1[4] dout1[5] dout1[6] dout1[7] dout1[8] dout1[9] dout1[10]
+ dout1[11] dout1[12] dout1[13] dout1[14] dout1[15] dout1[0] dout0[10] dout0[11] dout0[12]
+ dout0[13] dout0[14] dout0[15] dout0[16] addr0[0] wmask0[0] wmask0[1] wmask0[2] wmask0[3]
+ clk0 din0[0] din0[1] din0[2] din0[3] din0[4] din0[5] din0[6] din0[7] din0[8] din0[9]
+ din0[10] din0[11] din0[12] din0[13] din0[14] din0[15] din0[16] din0[17] din0[18]
+ din0[19] din0[20] din0[21] din0[22] dout0[0] dout0[1] dout0[2] dout0[3] dout0[4]
+ dout0[5] dout0[6] dout0[7] dout0[8] dout0[9] dout0[25] dout0[26] dout0[27] dout0[28]
+ dout0[29] dout0[30] dout0[31] din0[31] din0[23] din0[24] din0[25] din0[26] din0[27]
+ din0[28] din0[29] din0[30] dout0[17] dout0[18] dout0[19] dout0[20] dout0[21] dout0[22]
+ addr1[4] addr1[5] addr1[6] addr1[7] dout0[23] dout0[24] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/gnd_uq26
+ vssd1
Xsky130_sram_1kbyte_1rw1r_32x256_8_wmask_dff_0 sky130_sram_1kbyte_1rw1r_32x256_8_data_dff_0/clk
+ sky130_sram_1kbyte_1rw1r_32x256_8_wmask_dff_0/dout_0 wmask0[1] sky130_sram_1kbyte_1rw1r_32x256_8_wmask_dff_0/dout_1
+ wmask0[2] sky130_sram_1kbyte_1rw1r_32x256_8_wmask_dff_0/dout_2 wmask0[3] sky130_sram_1kbyte_1rw1r_32x256_8_wmask_dff_0/dout_3
+ vssd1 vccd1 wmask0[0] sky130_sram_1kbyte_1rw1r_32x256_8_wmask_dff
Xsky130_sram_1kbyte_1rw1r_32x256_8_bank_0 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/rbl_bl_1_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/rbl_bl_0_0 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/p_en_bar0
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/s_en0 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/w_en0
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/wl_en0 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/s_en1
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/p_en_bar1 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/wl_en1
+ sky130_sram_1kbyte_1rw1r_32x256_8_wmask_dff_0/dout_0 sky130_sram_1kbyte_1rw1r_32x256_8_wmask_dff_0/dout_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_wmask_dff_0/dout_2 sky130_sram_1kbyte_1rw1r_32x256_8_wmask_dff_0/dout_3
+ dout1[16] dout1[17] dout1[18] dout1[19] dout1[20] dout1[21] dout1[22] dout1[23]
+ dout1[24] dout1[25] dout1[26] dout1[27] dout1[28] dout1[29] dout1[30] dout1[31]
+ dout1[0] dout1[1] dout1[2] dout1[3] dout1[4] dout1[5] dout1[6] dout1[7] dout1[8]
+ dout1[9] dout1[10] dout1[11] dout1[12] dout1[13] dout1[14] dout1[15] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr0_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr0_2 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr0_3
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr0_4 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr0_5
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_0 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_2 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_3
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_4 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_5
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_6 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_7
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_8 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_9
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_10 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_11
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_12 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_13
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_14 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_15
+ dout0[0] dout0[1] dout0[2] dout0[3] dout0[4] dout0[5] dout0[6] dout0[7] dout0[8]
+ dout0[9] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14] dout0[15] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_23
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_24 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_25
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_26 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_27
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_28 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_29
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_30 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_31
+ dout0[16] dout0[17] dout0[18] dout0[19] dout0[20] dout0[21] dout0[22] dout0[23]
+ dout0[24] dout0[25] dout0[26] dout0[27] dout0[28] dout0[29] dout0[30] dout0[31]
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_16 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_17
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_18 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_19
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_20 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_22
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr1_1 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr1_2
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr1_3 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr1_4
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr1_5 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr1_6
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr1_7 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr0_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr1_0 vssd1 vssd1 vssd1 vssd1 vssd1 vssd1
+ vssd1 vssd1 vssd1 vssd1 vssd1 vssd1 vssd1 vssd1 vssd1 vssd1 vssd1 vssd1 vssd1 vssd1
+ vssd1 vssd1 vssd1 vssd1 vssd1 vssd1 vssd1 vssd1 vssd1 vssd1 vssd1 vssd1 vssd1 vssd1
+ vssd1 vssd1 vssd1 vssd1 vssd1 vssd1 vssd1 vssd1 vssd1 vssd1 vssd1 vssd1 vccd1 vccd1
+ vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1
+ vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1
+ vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1
+ vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1
+ vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1
+ vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/gnd_uq26
+ vccd1 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_21 vccd1 vssd1 vccd1 vccd1 vccd1
+ vccd1 vccd1 vccd1 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr0_7 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr0_6
+ vssd1 vccd1 vccd1 vccd1 vccd1 vssd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vssd1
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank
Xsky130_sram_1kbyte_1rw1r_32x256_8_control_logic_r_0 csb1 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/wl_en1
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/s_en1 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/rbl_bl_1_1
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/p_en_bar1 clk1 sky130_sram_1kbyte_1rw1r_32x256_8_row_addr_dff_0/clk
+ vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 vssd1 vccd1 sky130_sram_1kbyte_1rw1r_32x256_8_control_logic_r
Xsky130_sram_1kbyte_1rw1r_32x256_8_control_logic_rw_0 web0 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/wl_en0
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/w_en0 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/s_en0
+ sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/rbl_bl_0_0 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/p_en_bar0
+ clk0 sky130_sram_1kbyte_1rw1r_32x256_8_data_dff_0/clk vccd1 vccd1 vccd1 vccd1 vccd1
+ vccd1 vccd1 csb0 vccd1 vccd1 vccd1 vssd1 sky130_sram_1kbyte_1rw1r_32x256_8_control_logic_rw
Xsky130_sram_1kbyte_1rw1r_32x256_8_col_addr_dff_0 vccd1 vssd1 sky130_sram_1kbyte_1rw1r_32x256_8_data_dff_0/clk
+ addr0[0] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr0_0 sky130_sram_1kbyte_1rw1r_32x256_8_col_addr_dff
Xsky130_sram_1kbyte_1rw1r_32x256_8_col_addr_dff_1 vccd1 vssd1 sky130_sram_1kbyte_1rw1r_32x256_8_row_addr_dff_0/clk
+ addr1[0] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr1_0 sky130_sram_1kbyte_1rw1r_32x256_8_col_addr_dff
Xsky130_sram_1kbyte_1rw1r_32x256_8_row_addr_dff_0 vccd1 sky130_sram_1kbyte_1rw1r_32x256_8_row_addr_dff_0/clk
+ addr1[1] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr1_1 addr1[2] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr1_2
+ addr1[3] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr1_3 addr1[4] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr1_4
+ addr1[5] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr1_5 addr1[6] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr1_6
+ addr1[7] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr1_7 vccd1 vccd1 vccd1 vssd1
+ sky130_sram_1kbyte_1rw1r_32x256_8_row_addr_dff
Xsky130_sram_1kbyte_1rw1r_32x256_8_row_addr_dff_1 vccd1 sky130_sram_1kbyte_1rw1r_32x256_8_data_dff_0/clk
+ addr0[1] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr0_1 addr0[2] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr0_2
+ addr0[3] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr0_3 addr0[4] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr0_4
+ addr0[5] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr0_5 addr0[6] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr0_6
+ addr0[7] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/addr0_7 vccd1 vccd1 vccd1 vssd1
+ sky130_sram_1kbyte_1rw1r_32x256_8_row_addr_dff
Xsky130_sram_1kbyte_1rw1r_32x256_8_data_dff_0 sky130_sram_1kbyte_1rw1r_32x256_8_data_dff_0/clk
+ din0[0] din0[1] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_1 din0[2] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_2
+ din0[3] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_3 din0[4] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_4
+ din0[5] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_5 din0[6] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_6
+ din0[7] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_7 din0[8] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_8
+ din0[9] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_9 din0[10] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_10
+ din0[11] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_11 din0[12] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_12
+ din0[13] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_13 sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_14
+ din0[15] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_15 din0[16] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_16
+ din0[17] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_17 din0[18] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_18
+ din0[19] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_19 din0[20] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_20
+ din0[21] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_21 din0[22] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_22
+ din0[23] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_23 din0[24] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_24
+ din0[25] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_25 din0[26] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_26
+ din0[27] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_27 din0[28] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_28
+ din0[29] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_29 din0[30] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_30
+ din0[31] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_31 vssd1 vccd1 din0[14] sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/din0_0
+ sky130_sram_1kbyte_1rw1r_32x256_8_data_dff
.ends

.subckt sky130_fd_sc_hd__a22o_1 A1 A2 X B2 B1 VPWR VGND VNB VPB
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21oi_2 B1 A2 A1 Y VGND VPWR VNB VPB
X0 VGND A2 a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A1 a_114_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_114_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_285_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_8 A X VGND VPWR VNB VPB
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_12 A Y VGND VPWR VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_8 A Y VGND VPWR VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__bufbuf_8 A X VGND VPWR VNB VPB
X0 a_318_47# a_206_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_318_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_206_47# a_318_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_318_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_318_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_318_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_318_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_206_47# a_318_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR a_318_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_318_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_318_47# a_206_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_318_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_206_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X a_318_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_206_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR a_318_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND a_206_47# a_318_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND a_318_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND a_318_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VGND a_318_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 X a_318_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VGND a_318_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VPWR a_206_47# a_318_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 X a_318_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__bufinv_8 A Y VGND VPWR VNB VPB
X0 VPWR a_215_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_109_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND a_109_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND a_215_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_215_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR a_215_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND a_215_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND a_215_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR a_109_47# a_215_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_215_47# a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR a_215_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_215_47# a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR a_109_47# a_215_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR a_215_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 Y a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux2_8 S A1 VPWR VGND A0 X VNB VPB
X0 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_79_21# A0 a_792_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_1259_199# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_1302_47# A0 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_792_297# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_1259_199# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND a_1259_199# a_1302_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 a_79_21# A1 a_792_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15 a_79_21# A0 a_1302_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X16 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VPWR S a_792_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_792_297# A0 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1302_47# a_1259_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 VPWR a_1259_199# a_1302_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_1302_297# a_1259_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_792_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X27 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_1302_297# A1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND S a_792_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X30 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_79_21# A1 a_1302_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 a_792_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hd__fah_1 COUT B A SUM CI VPWR VGND VNB VPB
X0 a_508_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_1332_297# a_719_47# a_1262_49# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_27_47# a_508_297# a_719_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 VGND CI a_1262_49# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_67_199# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_508_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A a_310_49# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_310_49# B a_1008_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 a_508_297# a_1008_47# a_1332_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 a_1332_297# a_719_47# a_508_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X10 a_719_47# B a_310_49# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 a_1640_380# a_719_47# a_1617_49# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_1008_47# a_508_297# a_310_49# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 VGND a_1332_297# COUT VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_719_47# B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X15 a_1262_49# a_719_47# a_1617_49# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X16 SUM a_1617_49# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_1640_380# a_1262_49# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_1617_49# a_1008_47# a_1640_380# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X19 VPWR a_1332_297# COUT VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR a_67_199# a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_310_49# a_508_297# a_719_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22 a_67_199# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 VGND A a_310_49# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 a_27_47# B a_1008_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X25 a_1617_49# a_1008_47# a_1262_49# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X26 a_1640_380# a_1262_49# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X27 SUM a_1617_49# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 VPWR CI a_1262_49# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_1008_47# a_508_297# a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X30 VGND a_67_199# a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_1262_49# a_1008_47# a_1332_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_4 Y A B VGND VPWR VNB VPB
X0 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21a_1 X A1 B1 A2 VGND VPWR VNB VPB
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2b_2 B Y A_N VGND VPWR VNB VPB
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND B a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y a_27_93# a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_229_47# a_27_93# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y a_27_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_229_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand4_1 C B Y D A VPWR VGND VNB VPB
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_193_47# C a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y A a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_277_47# B a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o22ai_1 A2 B1 Y A1 B2 VGND VPWR VNB VPB
X0 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR A1 a_307_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_307_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 X A VGND VPWR VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_6 Y A VPWR VGND VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor4b_1 C B A D_N Y VGND VPWR VNB VPB
X0 Y a_91_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_91_199# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR A a_341_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_245_297# C a_161_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_341_297# B a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_91_199# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_161_297# a_91_199# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_2 Y A B VGND VPWR VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
.ends

.subckt sky130_fd_sc_hd__and3_4 A B C X VGND VPWR VNB VPB
X0 VPWR A a_94_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_294_47# B a_185_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_185_47# A a_94_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_94_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND C a_294_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_94_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_94_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_94_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR C a_94_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_94_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND a_94_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR a_94_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND a_94_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X a_94_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_4 VPWR VGND X A VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_2 Y A VPWR VGND VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfxtp_4 VGND VPWR D CLK Q VNB VPB
X0 Q a_1062_300# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_1020_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2 a_572_47# a_193_47# a_475_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 VPWR a_1062_300# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_634_183# a_475_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_475_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8 VGND a_1062_300# a_1020_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR a_634_183# a_568_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 Q a_1062_300# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_568_413# a_27_47# a_475_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_634_183# a_475_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X13 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_891_413# a_27_47# a_634_183# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 Q a_1062_300# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND a_891_413# a_1062_300# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR a_1062_300# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND a_1062_300# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 Q a_1062_300# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 VGND a_1062_300# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 VPWR a_891_413# a_1062_300# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_891_413# a_193_47# a_634_183# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X26 a_475_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 VGND a_634_183# a_572_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 VPWR a_1062_300# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2b_2 B_N A Y VGND VPWR VNB VPB
X0 Y a_251_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y a_251_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND a_251_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR B_N a_251_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND B_N a_251_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_27_297# a_251_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2b_1 Y A_N B VGND VPWR VNB VPB
X0 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 Y a_27_93# a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_206_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux2_4 X S A0 A1 VPWR VGND VNB VPB
X0 a_204_297# A1 a_396_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_396_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_396_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR S a_314_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_204_297# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_396_47# A0 a_314_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_206_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_396_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_396_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR a_396_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_490_47# A1 a_396_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND S a_490_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND a_396_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_396_47# A0 a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND a_396_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR S a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X a_396_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND S a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor3_2 C Y A B VGND VPWR VNB VPB
X0 Y C a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_281_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31o_1 A2 B1 A1 A3 X VGND VPWR VNB VPB
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2_1 A X B VGND VPWR VNB VPB
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__sdlclkp_2 SCE CLK GCLK GATE VGND VPWR VNB VPB
X0 GCLK a_1020_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_109_369# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_465_315# a_287_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_257_147# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_1102_47# a_465_315# a_1020_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND a_1020_47# GCLK VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_287_413# a_257_147# a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X7 VGND a_257_147# a_257_243# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR a_465_315# a_383_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND CLK a_1102_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_27_47# GATE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR CLK a_1020_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 GCLK a_1020_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_287_413# a_257_243# a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_383_413# a_257_147# a_287_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_257_147# CLK VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_27_47# GATE a_109_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 VPWR a_257_147# a_257_243# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X18 a_1020_47# a_465_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 a_395_47# a_257_243# a_287_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20 VGND a_465_315# a_395_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VPWR a_1020_47# GCLK VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND SCE a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_465_315# a_287_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfxtp_2 Q CLK D VPWR VGND VNB VPB
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2 VPWR a_1059_315# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND a_1059_315# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X14 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X19 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__bufbuf_16 A X VGND VPWR VNB VPB
X0 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_215_47# a_549_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND a_109_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_109_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_215_47# a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_549_47# a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND a_215_47# a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_549_47# a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_549_47# a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_549_47# a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_215_47# a_549_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_549_47# a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 VGND a_215_47# a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 VPWR a_109_47# a_215_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 a_215_47# a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X40 a_215_47# a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X41 VPWR a_109_47# a_215_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X42 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X43 VPWR a_215_47# a_549_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X44 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X45 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X46 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X47 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X48 a_549_47# a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X49 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X50 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X51 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__edfxbp_1 VPWR VGND CLK Q_N DE D Q VNB VPB
X0 a_381_369# D a_299_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 Q a_1591_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR DE a_423_343# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_1591_413# a_193_47# a_1514_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X5 Q_N a_791_264# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_986_413# a_193_47# a_299_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_1101_47# a_193_47# a_986_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8 VGND DE a_423_343# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_1500_413# a_1150_159# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_1514_47# a_1150_159# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 Q a_1591_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_1675_413# a_193_47# a_1591_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VPWR a_1591_413# a_791_264# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_1591_413# a_27_47# a_1500_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_729_47# a_423_343# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_729_369# DE VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X18 a_1077_413# a_27_47# a_986_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR a_791_264# a_1675_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_299_47# a_791_264# a_729_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND a_791_264# a_1717_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 a_1717_47# a_27_47# a_1591_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24 VPWR a_1150_159# a_1077_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_1150_159# a_986_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X26 a_986_413# a_27_47# a_299_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X27 a_299_47# a_791_264# a_729_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X28 VGND a_1591_413# a_791_264# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_381_47# D a_299_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 VGND a_1150_159# a_1101_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VPWR a_423_343# a_381_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X32 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VGND DE a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 a_1150_159# a_986_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X35 Q_N a_791_264# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_4 Y A B VGND VPWR VNB VPB
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__xor2_2 VPWR VGND X B A VNB VPB
X0 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_470_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_470_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_470_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_470_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR B a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND A a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X a_112_47# a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_470_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X B a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22o_4 B1 B2 X A2 A1 VGND VPWR VNB VPB
X0 a_484_297# B2 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND B2 a_566_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_96_21# B1 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_484_297# B1 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_484_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A2 a_918_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_96_21# B2 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_96_21# B1 a_566_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_484_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A1 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_96_21# A1 a_918_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VPWR A2 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_566_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_918_47# A1 a_96_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_566_47# B1 a_96_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_918_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3_1 Y A C B VGND VPWR VNB VPB
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_193_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__xor3_1 X C B A VGND VPWR VNB VPB
X0 a_112_21# C a_404_49# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_1198_49# a_931_365# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_386_325# B a_1198_49# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_404_49# a_266_93# a_112_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4 a_931_365# a_827_297# a_404_49# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X5 VPWR a_112_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_827_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_1198_49# a_827_297# a_404_49# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND A a_931_365# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 a_112_21# C a_386_325# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X10 a_1198_49# a_827_297# a_386_325# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 a_266_93# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_1198_49# a_931_365# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_931_365# a_827_297# a_386_325# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X14 VPWR A a_931_365# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_827_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND a_112_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_386_325# B a_931_365# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X18 a_266_93# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_404_49# B a_931_365# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X20 a_386_325# a_266_93# a_112_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 a_404_49# B a_1198_49# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2bb2ai_1 Y A1_N A2_N B2 B1 VGND VPWR VNB VPB
X0 VPWR A2_N a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y a_112_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND B2 a_394_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_112_297# A2_N a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_112_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_112_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR B1 a_478_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_394_47# a_112_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_394_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_478_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o32ai_1 A2 Y A1 A3 B2 B1 VGND VPWR VNB VPB
X0 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_333_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A1 a_461_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_461_297# A2 a_333_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22o_2 A1 A2 X B2 B1 VPWR VGND VNB VPB
X0 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_381_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor3b_1 C_N Y A B VGND VPWR VNB VPB
X0 VGND a_91_199# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR A a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_91_199# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_245_297# B a_161_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_91_199# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_161_297# a_91_199# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
.ends

.subckt sky130_fd_sc_hd__o31ai_1 Y A2 A1 A3 B1 VPWR VGND VNB VPB
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y A3 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_193_297# A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 X A VGND VPWR VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor4_1 D C Y A B VGND VPWR VNB VPB
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_191_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_297_297# B a_191_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2_4 X B A VGND VPWR VNB VPB
X0 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND B a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_110_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a211oi_1 A1 C1 B1 Y A2 VPWR VGND VNB VPB
X0 a_56_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A2 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_139_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_311_297# B1 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y C1 a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y A1 a_139_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
.ends

.subckt sky130_fd_sc_hd__nor2_2 B Y A VGND VPWR VNB VPB
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__xnor2_2 VGND VPWR Y A B VNB VPB
X0 a_27_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_560_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND B a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y a_27_297# a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_474_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_27_47# B a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_297# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_474_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_560_47# a_27_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR A a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR a_27_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_560_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__maj3_1 C X B A VGND VPWR VNB VPB
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_109_341# C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_27_47# B a_265_341# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_265_341# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR A a_109_341# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_421_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_265_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND C a_421_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_27_47# B a_265_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR C a_421_341# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_421_341# B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_109_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor4b_2 D_N Y C A B VGND VPWR VNB VPB
X0 VPWR D_N a_694_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_27_297# B a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_474_297# a_694_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_277_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y a_694_21# a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND D_N a_694_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_474_297# C a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y a_694_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_277_297# C a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND a_694_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2b_2 A B_N X VPWR VGND VNB VPB
X0 VPWR A a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_218_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_300_297# a_27_53# a_218_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_218_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR a_218_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_218_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_218_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND A a_218_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4_1 C A X B D VPWR VGND VNB VPB
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a221oi_1 Y C1 A1 A2 B2 B1 VGND VPWR VNB VPB
X0 a_465_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_204_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y B1 a_204_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_109_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a32oi_1 A2 Y A1 B2 B1 A3 VGND VPWR VNB VPB
X0 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A3 a_383_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_309_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_383_47# A2 a_309_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31oi_1 VGND VPWR Y B1 A2 A1 A3 VNB VPB
X0 Y A1 a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_181_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21o_2 X B1 A1 A2 VGND VPWR VNB VPB
X0 VPWR a_80_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_80_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_80_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_386_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_80_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_80_199# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_386_297# B1 a_80_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_458_47# A1 a_80_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A1 a_386_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A2 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor3_1 C Y A B VGND VPWR VNB VPB
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a221o_1 X B1 A1 B2 A2 VGND VPWR C1 VNB VPB
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__sdlclkp_1 SCE CLK GCLK GATE VGND VPWR VNB VPB
X0 a_1094_47# a_464_315# a_1012_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_464_315# a_286_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_464_315# a_286_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR CLK a_1012_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_1012_47# a_464_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_109_369# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 VPWR a_464_315# a_382_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_382_413# a_256_147# a_286_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_286_413# a_256_243# a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_27_47# GATE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_256_147# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 VGND a_256_147# a_256_243# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 GCLK a_1012_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_27_47# GATE a_109_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 a_256_147# CLK VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 GCLK a_1012_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR a_256_147# a_256_243# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 a_286_413# a_256_147# a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X18 VGND CLK a_1094_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_394_47# a_256_243# a_286_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20 VGND a_464_315# a_394_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND SCE a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and3_1 VGND VPWR X B A C VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_1 Y A VGND VPWR VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__bufinv_16 A Y VGND VPWR VNB VPB
X0 a_361_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_361_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_27_47# a_361_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_361_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_361_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR a_27_47# a_361_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_361_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 VGND a_27_47# a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 VPWR a_27_47# a_361_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 VGND a_27_47# a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X38 VGND a_27_47# a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 a_361_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X41 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X42 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X43 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X44 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X45 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X46 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X47 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X48 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X49 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o31ai_2 A1 Y B1 A3 A2 VGND VPWR VNB VPB
X0 a_281_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_281_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y A3 a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_297# A2 a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt user_proj_example la_data_in[127] la_data_in[126] la_data_in[125] la_data_in[124]
+ la_data_in[123] la_data_in[122] la_data_in[121] la_data_in[120] la_data_in[119]
+ la_data_in[118] la_data_in[117] la_data_in[116] la_data_in[115] la_data_in[114]
+ la_data_in[113] la_data_in[112] la_data_in[111] la_data_in[110] la_data_in[109]
+ la_data_in[108] la_data_in[107] la_data_in[106] la_data_in[105] la_data_in[104]
+ la_data_in[103] la_data_in[102] la_data_in[101] la_data_in[100] la_data_in[99] la_data_in[98]
+ la_data_in[97] la_data_in[96] la_data_in[95] la_data_in[94] la_data_in[93] la_data_in[92]
+ la_data_in[91] la_data_in[90] la_data_in[89] la_data_in[88] la_data_in[87] la_data_in[86]
+ la_data_in[85] la_data_in[84] la_data_in[83] la_data_in[82] la_data_in[81] la_data_in[80]
+ la_data_in[79] la_data_in[78] la_data_in[77] la_data_in[76] la_data_in[75] la_data_in[74]
+ la_data_in[73] la_data_in[72] la_data_in[71] la_data_in[70] la_data_in[69] la_data_in[68]
+ la_data_in[67] la_data_in[66] la_data_in[65] la_data_in[64] la_data_in[63] la_data_in[62]
+ la_data_in[61] la_data_in[60] la_data_in[59] la_data_in[58] la_data_in[57] la_data_in[56]
+ la_data_in[55] la_data_in[54] la_data_in[53] la_data_in[52] la_data_in[51] la_data_in[50]
+ la_data_in[49] la_data_in[48] la_data_in[47] la_data_in[46] la_data_in[45] la_data_in[44]
+ la_data_in[43] la_data_in[42] la_data_in[41] la_data_in[40] la_data_in[39] la_data_in[38]
+ la_data_in[37] la_data_in[36] la_data_in[35] la_data_in[34] la_data_in[33] la_data_in[32]
+ la_data_in[31] la_data_in[30] la_data_in[29] la_data_in[28] la_data_in[27] la_data_in[26]
+ la_data_in[25] la_data_in[24] la_data_in[23] la_data_in[22] la_data_in[21] la_data_in[20]
+ la_data_in[19] la_data_in[18] la_data_in[17] la_data_in[16] la_data_in[15] la_data_in[14]
+ la_data_in[13] la_data_in[12] la_data_in[11] la_data_in[10] la_data_in[9] la_data_in[8]
+ la_data_in[7] la_data_in[6] la_data_in[5] la_data_in[4] la_data_in[3] la_data_in[2]
+ la_data_in[1] la_data_in[0] la_data_out[127] la_data_out[126] la_data_out[125] la_data_out[124]
+ la_data_out[123] la_data_out[122] la_data_out[121] la_data_out[120] la_data_out[119]
+ la_data_out[118] la_data_out[117] la_data_out[116] la_data_out[115] la_data_out[114]
+ la_data_out[113] la_data_out[112] la_data_out[111] la_data_out[110] la_data_out[109]
+ la_data_out[108] la_data_out[107] la_data_out[106] la_data_out[105] la_data_out[104]
+ la_data_out[103] la_data_out[102] la_data_out[101] la_data_out[100] la_data_out[99]
+ la_data_out[98] la_data_out[97] la_data_out[96] la_data_out[95] la_data_out[94]
+ la_data_out[93] la_data_out[92] la_data_out[91] la_data_out[90] la_data_out[89]
+ la_data_out[88] la_data_out[87] la_data_out[86] la_data_out[85] la_data_out[84]
+ la_data_out[83] la_data_out[82] la_data_out[81] la_data_out[80] la_data_out[79]
+ la_data_out[78] la_data_out[77] la_data_out[76] la_data_out[75] la_data_out[74]
+ la_data_out[73] la_data_out[72] la_data_out[71] la_data_out[70] la_data_out[69]
+ la_data_out[68] la_data_out[67] la_data_out[66] la_data_out[65] la_data_out[64]
+ la_data_out[63] la_data_out[62] la_data_out[61] la_data_out[60] la_data_out[59]
+ la_data_out[58] la_data_out[57] la_data_out[56] la_data_out[55] la_data_out[54]
+ la_data_out[53] la_data_out[52] la_data_out[51] la_data_out[50] la_data_out[49]
+ la_data_out[48] la_data_out[47] la_data_out[46] la_data_out[45] la_data_out[44]
+ la_data_out[43] la_data_out[42] la_data_out[41] la_data_out[40] la_data_out[39]
+ la_data_out[38] la_data_out[37] la_data_out[36] la_data_out[35] la_data_out[34]
+ la_data_out[33] la_data_out[32] la_data_out[31] la_data_out[30] la_data_out[29]
+ la_data_out[28] la_data_out[27] la_data_out[26] la_data_out[25] la_data_out[24]
+ la_data_out[23] la_data_out[22] la_data_out[21] la_data_out[20] la_data_out[19]
+ la_data_out[18] la_data_out[17] la_data_out[16] la_data_out[15] la_data_out[14]
+ la_data_out[13] la_data_out[12] la_data_out[11] la_data_out[10] la_data_out[9] la_data_out[8]
+ la_data_out[7] la_data_out[6] la_data_out[5] la_data_out[4] la_data_out[3] la_data_out[2]
+ la_data_out[1] la_data_out[0] la_oenb[127] la_oenb[126] la_oenb[125] la_oenb[124]
+ la_oenb[123] la_oenb[122] la_oenb[121] la_oenb[120] la_oenb[119] la_oenb[118] la_oenb[117]
+ la_oenb[116] la_oenb[115] la_oenb[114] la_oenb[113] la_oenb[112] la_oenb[111] la_oenb[110]
+ la_oenb[109] la_oenb[108] la_oenb[107] la_oenb[106] la_oenb[105] la_oenb[104] la_oenb[103]
+ la_oenb[102] la_oenb[101] la_oenb[100] la_oenb[99] la_oenb[98] la_oenb[97] la_oenb[96]
+ la_oenb[95] la_oenb[94] la_oenb[93] la_oenb[92] la_oenb[91] la_oenb[90] la_oenb[89]
+ la_oenb[88] la_oenb[87] la_oenb[86] la_oenb[85] la_oenb[84] la_oenb[83] la_oenb[82]
+ la_oenb[81] la_oenb[80] la_oenb[79] la_oenb[78] la_oenb[77] la_oenb[76] la_oenb[75]
+ la_oenb[74] la_oenb[73] la_oenb[72] la_oenb[71] la_oenb[70] la_oenb[69] la_oenb[68]
+ la_oenb[67] la_oenb[66] la_oenb[65] la_oenb[64] la_oenb[63] la_oenb[62] la_oenb[61]
+ la_oenb[60] la_oenb[59] la_oenb[58] la_oenb[57] la_oenb[56] la_oenb[55] la_oenb[54]
+ la_oenb[53] la_oenb[52] la_oenb[51] la_oenb[50] la_oenb[49] la_oenb[48] la_oenb[47]
+ la_oenb[46] la_oenb[45] la_oenb[44] la_oenb[43] la_oenb[42] la_oenb[41] la_oenb[40]
+ la_oenb[39] la_oenb[38] la_oenb[37] la_oenb[36] la_oenb[35] la_oenb[34] la_oenb[33]
+ la_oenb[32] la_oenb[31] la_oenb[30] la_oenb[29] la_oenb[28] la_oenb[27] la_oenb[26]
+ la_oenb[25] la_oenb[24] la_oenb[23] la_oenb[22] la_oenb[21] la_oenb[20] la_oenb[19]
+ la_oenb[18] la_oenb[17] la_oenb[16] la_oenb[15] la_oenb[14] la_oenb[13] la_oenb[12]
+ la_oenb[11] la_oenb[10] la_oenb[9] la_oenb[8] la_oenb[7] la_oenb[6] la_oenb[5] la_oenb[4]
+ la_oenb[3] la_oenb[2] la_oenb[1] la_oenb[0] io_in[37] io_in[36] io_in[35] io_in[34]
+ io_in[33] io_in[32] io_in[31] io_in[30] io_in[29] io_in[28] io_in[27] io_in[26]
+ io_in[25] io_in[24] io_in[23] io_in[22] io_in[21] io_in[20] io_in[19] io_in[18]
+ io_in[17] io_in[16] io_in[15] io_in[14] io_in[13] io_in[12] io_in[11] io_in[10]
+ io_in[9] io_in[8] io_in[7] io_in[6] io_in[5] io_in[4] io_in[3] io_in[2] io_in[1]
+ io_in[0] io_out[37] io_out[36] io_out[35] io_out[34] io_out[33] io_out[32] io_out[31]
+ io_out[30] io_out[29] io_out[28] io_out[27] io_out[26] io_out[25] io_out[24] io_out[23]
+ io_out[22] io_out[21] io_out[20] io_out[19] io_out[18] io_out[17] io_out[16] io_out[15]
+ io_out[14] io_out[13] io_out[12] io_out[11] io_out[10] io_out[9] io_out[8] io_out[7]
+ io_out[6] io_out[5] io_out[4] io_out[3] io_out[2] io_out[1] io_out[0] io_oeb[37]
+ io_oeb[36] io_oeb[35] io_oeb[34] io_oeb[33] io_oeb[32] io_oeb[31] io_oeb[30] io_oeb[29]
+ io_oeb[28] io_oeb[27] io_oeb[26] io_oeb[25] io_oeb[24] io_oeb[23] io_oeb[22] io_oeb[21]
+ io_oeb[20] io_oeb[19] io_oeb[18] io_oeb[17] io_oeb[16] io_oeb[15] io_oeb[14] io_oeb[13]
+ io_oeb[12] io_oeb[11] io_oeb[10] io_oeb[9] io_oeb[8] io_oeb[7] io_oeb[6] io_oeb[5]
+ io_oeb[4] io_oeb[3] io_oeb[2] io_oeb[1] io_oeb[0] user_irq[2] user_irq[1] user_irq[0]
+ user_clock2 analog_io[28] analog_io[27] analog_io[26] analog_io[25] analog_io[24]
+ analog_io[23] analog_io[22] analog_io[21] analog_io[20] analog_io[19] analog_io[18]
+ analog_io[17] analog_io[16] analog_io[15] analog_io[14] analog_io[13] analog_io[12]
+ analog_io[11] analog_io[10] analog_io[9] analog_io[8] analog_io[7] analog_io[6]
+ analog_io[5] analog_io[4] analog_io[3] analog_io[2] analog_io[1] analog_io[0] wb_clk_i
+ wb_rst_i wbs_stb_i wbs_cyc_i wbs_we_i wbs_sel_i[3] wbs_sel_i[2] wbs_sel_i[1] wbs_sel_i[0]
+ wbs_dat_i[31] wbs_dat_i[30] wbs_dat_i[29] wbs_dat_i[28] wbs_dat_i[27] wbs_dat_i[26]
+ wbs_dat_i[25] wbs_dat_i[24] wbs_dat_i[23] wbs_dat_i[22] wbs_dat_i[21] wbs_dat_i[20]
+ wbs_dat_i[19] wbs_dat_i[18] wbs_dat_i[17] wbs_dat_i[16] wbs_dat_i[15] wbs_dat_i[14]
+ wbs_dat_i[13] wbs_dat_i[12] wbs_dat_i[11] wbs_dat_i[10] wbs_dat_i[9] wbs_dat_i[8]
+ wbs_dat_i[7] wbs_dat_i[6] wbs_dat_i[5] wbs_dat_i[4] wbs_dat_i[3] wbs_dat_i[2] wbs_dat_i[1]
+ wbs_dat_i[0] wbs_adr_i[31] wbs_adr_i[30] wbs_adr_i[29] wbs_adr_i[28] wbs_adr_i[27]
+ wbs_adr_i[26] wbs_adr_i[25] wbs_adr_i[24] wbs_adr_i[23] wbs_adr_i[22] wbs_adr_i[21]
+ wbs_adr_i[20] wbs_adr_i[19] wbs_adr_i[18] wbs_adr_i[17] wbs_adr_i[16] wbs_adr_i[15]
+ wbs_adr_i[14] wbs_adr_i[13] wbs_adr_i[12] wbs_adr_i[11] wbs_adr_i[10] wbs_adr_i[9]
+ wbs_adr_i[8] wbs_adr_i[7] wbs_adr_i[6] wbs_adr_i[5] wbs_adr_i[4] wbs_adr_i[3] wbs_adr_i[2]
+ wbs_adr_i[1] wbs_adr_i[0] wbs_ack_o wbs_dat_o[31] wbs_dat_o[30] wbs_dat_o[29] wbs_dat_o[28]
+ wbs_dat_o[27] wbs_dat_o[26] wbs_dat_o[25] wbs_dat_o[24] wbs_dat_o[23] wbs_dat_o[22]
+ wbs_dat_o[21] wbs_dat_o[20] wbs_dat_o[19] wbs_dat_o[18] wbs_dat_o[17] wbs_dat_o[16]
+ wbs_dat_o[15] wbs_dat_o[14] wbs_dat_o[13] wbs_dat_o[12] wbs_dat_o[11] wbs_dat_o[10]
+ wbs_dat_o[9] wbs_dat_o[8] wbs_dat_o[7] wbs_dat_o[6] wbs_dat_o[5] wbs_dat_o[4] wbs_dat_o[3]
+ wbs_dat_o[2] wbs_dat_o[1] wbs_dat_o[0] vssd1 vccd1
Xsky130_fd_sc_hd__decap_12_1780 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1791 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_90 sky130_fd_sc_hd__inv_2_90/A sky130_fd_sc_hd__inv_2_90/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__ha_2_11 vssd1 vccd1 sky130_fd_sc_hd__ha_2_11/A sky130_fd_sc_hd__fa_2_429/B
+ sky130_fd_sc_hd__ha_2_11/SUM sky130_fd_sc_hd__ha_2_11/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_22 vssd1 vccd1 la_data_out[61] sky130_fd_sc_hd__ha_2_21/B sky130_fd_sc_hd__ha_2_22/SUM
+ sky130_fd_sc_hd__ha_2_22/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_33 vssd1 vccd1 sky130_fd_sc_hd__ha_2_33/A sky130_fd_sc_hd__xor2_1_691/A
+ sky130_fd_sc_hd__ha_2_33/SUM sky130_fd_sc_hd__ha_2_33/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_44 vssd1 vccd1 sky130_fd_sc_hd__or4_1_3/D sky130_fd_sc_hd__ha_2_43/B
+ sky130_fd_sc_hd__ha_2_44/SUM sky130_fd_sc_hd__ha_2_44/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__and2b_4_6 sky130_fd_sc_hd__nor2_4_14/A sky130_fd_sc_hd__and2b_4_6/X
+ sky130_fd_sc_hd__and3_4_12/C vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__and2b_4
Xsky130_fd_sc_hd__ha_2_55 vssd1 vccd1 sky130_fd_sc_hd__ha_2_55/A sky130_fd_sc_hd__ha_2_54/B
+ sky130_fd_sc_hd__ha_2_55/SUM sky130_fd_sc_hd__ha_2_55/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_7 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_7/X sky130_fd_sc_hd__xnor2_2_0/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__sdlclkp_4_40 sky130_fd_sc_hd__conb_1_145/LO sky130_fd_sc_hd__clkinv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_392/CLK sky130_fd_sc_hd__o21ai_1_892/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_51 sky130_fd_sc_hd__conb_1_148/LO sky130_fd_sc_hd__clkinv_2_48/Y
+ sky130_fd_sc_hd__dfxtp_1_498/CLK sky130_fd_sc_hd__o21ai_2_18/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_120 sky130_fd_sc_hd__or2_0_61/A sky130_fd_sc_hd__nor2_1_120/Y
+ sky130_fd_sc_hd__or2_0_60/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_131 sky130_fd_sc_hd__nor2_1_73/B sky130_fd_sc_hd__nor2_1_131/Y
+ sky130_fd_sc_hd__buf_6_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_142 sky130_fd_sc_hd__nor2_1_142/B sky130_fd_sc_hd__nor2_1_142/Y
+ sky130_fd_sc_hd__nor2_1_142/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_153 sky130_fd_sc_hd__nor2_2_16/Y sky130_fd_sc_hd__nor2_1_153/Y
+ sky130_fd_sc_hd__nor2_2_17/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_1_7 la_data_out[120] sky130_fd_sc_hd__clkinv_1_7/A vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_164 sky130_fd_sc_hd__nor2_1_164/B sky130_fd_sc_hd__nor2_1_164/Y
+ sky130_fd_sc_hd__nor2_1_164/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_40 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__clkbuf_1_25/X
+ sky130_fd_sc_hd__nand2_1_79/B sky130_fd_sc_hd__dfxtp_1_131/Q sky130_fd_sc_hd__a22oi_1_40/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_175 sky130_fd_sc_hd__nor2_1_175/B sky130_fd_sc_hd__nor2_1_175/Y
+ sky130_fd_sc_hd__nor2_1_177/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_51 sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__dfxtp_1_104/Q sky130_fd_sc_hd__dfxtp_1_72/Q sky130_fd_sc_hd__a22oi_1_51/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_186 sky130_fd_sc_hd__and3_4_25/A sky130_fd_sc_hd__nor2_1_186/Y
+ sky130_fd_sc_hd__and3_4_25/C vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_62 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__nor2_4_3/Y
+ sky130_fd_sc_hd__nand2_1_68/B sky130_fd_sc_hd__dfxtp_1_142/Q sky130_fd_sc_hd__a22oi_1_62/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_73 sky130_fd_sc_hd__clkbuf_1_24/X sky130_fd_sc_hd__clkbuf_1_23/X
+ sky130_fd_sc_hd__dfxtp_1_115/Q sky130_fd_sc_hd__dfxtp_1_83/Q sky130_fd_sc_hd__a22oi_1_73/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_197 sky130_fd_sc_hd__nor2_1_202/Y sky130_fd_sc_hd__nor2_1_197/Y
+ sky130_fd_sc_hd__nor2_1_199/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_84 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__nor2_4_3/Y
+ sky130_fd_sc_hd__nand2_1_56/B sky130_fd_sc_hd__dfxtp_1_153/Q sky130_fd_sc_hd__a22oi_1_84/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_95 sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__dfxtp_1_126/Q sky130_fd_sc_hd__dfxtp_1_94/Q sky130_fd_sc_hd__a22oi_1_95/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_360 sky130_fd_sc_hd__buf_12_71/X sky130_fd_sc_hd__buf_12_566/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_371 sky130_fd_sc_hd__buf_12_72/X sky130_fd_sc_hd__buf_12_541/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_382 sky130_fd_sc_hd__buf_12_382/A sky130_fd_sc_hd__buf_12_464/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_393 sky130_fd_sc_hd__buf_12_393/A sky130_fd_sc_hd__buf_12_646/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xnor2_1_101 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_383/B sky130_fd_sc_hd__nor2_2_19/A
+ sky130_fd_sc_hd__xnor2_1_99/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_112 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_112/B sky130_fd_sc_hd__inv_2_31/A
+ sky130_fd_sc_hd__xnor2_1_112/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_560 sky130_fd_sc_hd__nor2_1_181/B sky130_fd_sc_hd__nand2_1_569/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_123 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_123/B sky130_fd_sc_hd__xnor2_1_123/Y
+ sky130_fd_sc_hd__xnor2_1_123/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_571 sky130_fd_sc_hd__nand2_1_577/A sky130_fd_sc_hd__nor2_1_185/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_134 vssd1 vccd1 sky130_fd_sc_hd__fa_2_310/A sky130_fd_sc_hd__nor2_1_167/B
+ sky130_fd_sc_hd__xnor2_1_134/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_582 sky130_fd_sc_hd__xnor2_1_166/B sky130_fd_sc_hd__o21ai_2_16/A2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_145 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_145/B sky130_fd_sc_hd__inv_2_55/A
+ sky130_fd_sc_hd__xnor2_1_145/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_593 sky130_fd_sc_hd__nand2_1_619/A sky130_fd_sc_hd__nor2_1_204/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_156 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_156/B sky130_fd_sc_hd__xnor2_1_156/Y
+ sky130_fd_sc_hd__xnor2_1_156/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_167 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_167/B sky130_fd_sc_hd__inv_2_47/A
+ sky130_fd_sc_hd__xnor2_1_167/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_178 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_180/A sky130_fd_sc_hd__and3_4_21/C
+ sky130_fd_sc_hd__xor2_1_622/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_4_40 sky130_fd_sc_hd__clkinv_4_40/A sky130_fd_sc_hd__clkinv_8_23/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__xnor2_1_189 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_189/B sky130_fd_sc_hd__and2_0_275/A
+ sky130_fd_sc_hd__xnor2_1_189/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_4_51 sky130_fd_sc_hd__clkinv_4_51/A sky130_fd_sc_hd__clkinv_4_51/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_62 sky130_fd_sc_hd__clkinv_4_62/A sky130_fd_sc_hd__clkinv_4_62/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_73 sky130_fd_sc_hd__clkinv_4_73/A sky130_fd_sc_hd__clkinv_4_73/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_84 wbs_dat_i[22] sky130_fd_sc_hd__clkinv_4_84/Y vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_1010 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_4_95 sky130_fd_sc_hd__nand2_1_17/Y sky130_fd_sc_hd__clkinv_4_95/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_1021 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1032 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1043 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1054 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1065 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__decap_12_1076 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_507 vssd1 vccd1 sky130_fd_sc_hd__buf_2_8/X sky130_fd_sc_hd__nand2b_1_8/Y
+ sky130_fd_sc_hd__o21ai_1_507/B1 sky130_fd_sc_hd__xor2_1_306/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1087 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_518 vssd1 vccd1 sky130_fd_sc_hd__inv_2_27/Y sky130_fd_sc_hd__nand2b_1_13/Y
+ sky130_fd_sc_hd__nand2_1_325/Y sky130_fd_sc_hd__xor2_1_316/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1098 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_529 vssd1 vccd1 sky130_fd_sc_hd__inv_2_29/Y sky130_fd_sc_hd__nand2b_1_8/Y
+ sky130_fd_sc_hd__o21ai_1_529/B1 sky130_fd_sc_hd__xor2_1_328/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__and2b_4_10 sky130_fd_sc_hd__nor2_4_18/A sky130_fd_sc_hd__and2b_4_10/X
+ sky130_fd_sc_hd__and3_4_22/C vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__and2b_4
Xsky130_fd_sc_hd__xor2_1_301 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__fa_2_207/A
+ sky130_fd_sc_hd__xor2_1_301/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_312 sky130_fd_sc_hd__dfxtp_2_5/Q sky130_fd_sc_hd__fa_2_209/A
+ sky130_fd_sc_hd__xor2_1_312/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_323 sky130_fd_sc_hd__dfxtp_2_5/Q sky130_fd_sc_hd__xor2_1_323/X
+ sky130_fd_sc_hd__xor2_1_323/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_334 sky130_fd_sc_hd__fa_2_262/A sky130_fd_sc_hd__xor2_1_334/X
+ sky130_fd_sc_hd__xor2_1_334/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_345 sky130_fd_sc_hd__dfxtp_2_5/Q sky130_fd_sc_hd__fa_2_235/A
+ sky130_fd_sc_hd__xor2_1_345/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_356 sky130_fd_sc_hd__dfxtp_2_5/Q sky130_fd_sc_hd__fah_1_4/A
+ sky130_fd_sc_hd__xor2_1_356/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_367 sky130_fd_sc_hd__xor2_1_367/B sky130_fd_sc_hd__xor2_1_367/X
+ sky130_fd_sc_hd__xor2_1_367/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_378 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__xor2_1_378/X
+ sky130_fd_sc_hd__xor2_1_378/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_389 sky130_fd_sc_hd__xor2_1_389/B sky130_fd_sc_hd__xor2_1_389/X
+ sky130_fd_sc_hd__xor2_1_389/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_305 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_305/X sky130_fd_sc_hd__buf_12_81/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_316 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_316/X sky130_fd_sc_hd__clkinv_1_899/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_327 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_275/A sky130_fd_sc_hd__nor4b_1_0/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_338 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1_7/D sky130_fd_sc_hd__dfxtp_1_8/Q
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_409 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__or2_0_60/B
+ sky130_fd_sc_hd__or2_0_60/A sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__or2_0_61/A
+ sky130_fd_sc_hd__o21ai_1_677/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_349 vssd1 vccd1 sky130_fd_sc_hd__inv_4_2/A sky130_fd_sc_hd__a222oi_1_7/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_20 sky130_fd_sc_hd__dfxtp_1_20/Q sky130_fd_sc_hd__dfxtp_1_20/CLK
+ la_data_out[36] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_31 sky130_fd_sc_hd__nand2_1_81/B sky130_fd_sc_hd__dfxtp_1_46/CLK
+ sky130_fd_sc_hd__dfxtp_1_31/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_42 sky130_fd_sc_hd__nand2_1_72/B sky130_fd_sc_hd__dfxtp_1_43/CLK
+ sky130_fd_sc_hd__dfxtp_1_42/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_53 sky130_fd_sc_hd__nand2_1_61/B sky130_fd_sc_hd__dfxtp_1_57/CLK
+ sky130_fd_sc_hd__dfxtp_1_53/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_64 sky130_fd_sc_hd__dfxtp_1_64/Q sky130_fd_sc_hd__dfxtp_1_65/CLK
+ sky130_fd_sc_hd__dfxtp_1_64/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_75 sky130_fd_sc_hd__dfxtp_1_75/Q sky130_fd_sc_hd__dfxtp_1_81/CLK
+ sky130_fd_sc_hd__dfxtp_1_75/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_86 sky130_fd_sc_hd__dfxtp_1_86/Q sky130_fd_sc_hd__dfxtp_1_89/CLK
+ sky130_fd_sc_hd__dfxtp_1_86/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_97 sky130_fd_sc_hd__dfxtp_1_97/Q sky130_fd_sc_hd__dfxtp_1_97/CLK
+ sky130_fd_sc_hd__dfxtp_1_97/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_303 vccd1 vssd1 sky130_fd_sc_hd__and2_0_303/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_303/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_314 vccd1 vssd1 sky130_fd_sc_hd__and2_0_314/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_314/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_325 vccd1 vssd1 sky130_fd_sc_hd__and2_0_325/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_325/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_336 vccd1 vssd1 sky130_fd_sc_hd__and2_0_397/A sky130_fd_sc_hd__ha_2_41/SUM
+ sky130_fd_sc_hd__and2_0_342/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_347 vccd1 vssd1 sky130_fd_sc_hd__and2_0_347/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__buf_2_43/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_358 vccd1 vssd1 sky130_fd_sc_hd__and2_0_358/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__buf_2_47/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_369 vccd1 vssd1 sky130_fd_sc_hd__and2_0_369/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_61/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__inv_2_103 sky130_fd_sc_hd__inv_2_199/Y sky130_fd_sc_hd__inv_2_103/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_114 sky130_fd_sc_hd__inv_2_114/A sky130_fd_sc_hd__inv_2_114/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__or2_0_5 sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__or2_0_5/X sky130_fd_sc_hd__or2_0_5/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__inv_2_125 sky130_fd_sc_hd__inv_2_125/A sky130_fd_sc_hd__inv_2_125/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_136 sky130_fd_sc_hd__inv_2_136/A sky130_fd_sc_hd__inv_2_136/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_147 sky130_fd_sc_hd__inv_2_147/A sky130_fd_sc_hd__buf_8_44/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_158 sky130_fd_sc_hd__inv_12_1/Y sky130_fd_sc_hd__inv_2_158/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_169 sky130_fd_sc_hd__inv_2_169/A sky130_fd_sc_hd__inv_2_170/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_12_190 sky130_fd_sc_hd__buf_4_36/X sky130_fd_sc_hd__buf_12_407/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_390 sky130_fd_sc_hd__a21oi_1_61/B1 sky130_fd_sc_hd__nand2_1_295/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a211o_1_4 vssd1 vccd1 sky130_fd_sc_hd__fa_2_280/A sky130_fd_sc_hd__dfxtp_1_67/Q
+ sky130_fd_sc_hd__nor2_1_8/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_4/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__o21ai_1_304 vssd1 vccd1 sky130_fd_sc_hd__inv_2_17/Y sky130_fd_sc_hd__nand2b_2_0/Y
+ sky130_fd_sc_hd__o21ai_1_304/B1 sky130_fd_sc_hd__xor2_1_124/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_315 vssd1 vccd1 sky130_fd_sc_hd__inv_2_18/Y sky130_fd_sc_hd__nand2b_2_0/Y
+ sky130_fd_sc_hd__o21ai_1_315/B1 sky130_fd_sc_hd__xor2_1_135/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_326 vssd1 vccd1 sky130_fd_sc_hd__inv_2_11/Y sky130_fd_sc_hd__nand2_1_245/Y
+ sky130_fd_sc_hd__a21oi_1_51/Y sky130_fd_sc_hd__xnor2_1_37/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_337 vssd1 vccd1 sky130_fd_sc_hd__inv_2_9/Y sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__o21ai_1_337/B1 sky130_fd_sc_hd__xor2_1_156/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_348 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_171/A sky130_fd_sc_hd__nor2_1_88/Y
+ sky130_fd_sc_hd__nand2_1_271/Y sky130_fd_sc_hd__xnor2_1_44/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_359 vssd1 vccd1 sky130_fd_sc_hd__inv_2_18/Y sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__o21ai_1_359/B1 sky130_fd_sc_hd__xor2_1_175/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nand2_1_708 sky130_fd_sc_hd__xor2_1_651/B sky130_fd_sc_hd__nand2_1_709/Y
+ sky130_fd_sc_hd__nand2_1_708/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_719 sky130_fd_sc_hd__o22ai_1_98/B2 sky130_fd_sc_hd__xnor2_2_6/Y
+ sky130_fd_sc_hd__xor2_1_668/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_17 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_17/A1 sky130_fd_sc_hd__buf_2_77/X
+ sky130_fd_sc_hd__mux2_8_0/S sky130_fd_sc_hd__or2_0_74/B vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_28 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_28/A1 sky130_fd_sc_hd__buf_4_23/X
+ sky130_fd_sc_hd__mux2_8_1/S sky130_fd_sc_hd__or2_0_78/B vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_39 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_39/A1 sky130_fd_sc_hd__buf_2_95/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__mux2_2_39/X vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__conb_1_103 sky130_fd_sc_hd__conb_1_103/LO sky130_fd_sc_hd__conb_1_103/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_114 sky130_fd_sc_hd__conb_1_114/LO sky130_fd_sc_hd__conb_1_114/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_125 sky130_fd_sc_hd__conb_1_125/LO sky130_fd_sc_hd__conb_1_125/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_136 sky130_fd_sc_hd__conb_1_136/LO sky130_fd_sc_hd__clkinv_1_6/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_147 sky130_fd_sc_hd__conb_1_147/LO sky130_fd_sc_hd__conb_1_147/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__xor2_1_120 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__fa_2_87/CIN
+ sky130_fd_sc_hd__xor2_1_120/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_131 sky130_fd_sc_hd__fa_2_97/A sky130_fd_sc_hd__and3_4_6/A
+ sky130_fd_sc_hd__xor2_1_131/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_142 sky130_fd_sc_hd__xor2_1_6/B sky130_fd_sc_hd__fa_2_104/B
+ sky130_fd_sc_hd__xor2_1_142/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_153 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__fa_2_109/A
+ sky130_fd_sc_hd__xor2_1_153/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_504 sky130_fd_sc_hd__ha_2_43/A sky130_fd_sc_hd__dfxtp_1_509/CLK
+ sky130_fd_sc_hd__and2_0_390/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_164 sky130_fd_sc_hd__fa_2_122/A sky130_fd_sc_hd__fa_2_118/B
+ sky130_fd_sc_hd__xor2_1_164/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_515 sky130_fd_sc_hd__ha_2_55/A sky130_fd_sc_hd__dfxtp_1_515/CLK
+ sky130_fd_sc_hd__and2_0_348/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_175 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__fa_2_126/A
+ sky130_fd_sc_hd__xor2_1_175/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_526 wbs_dat_o[5] sky130_fd_sc_hd__dfxtp_1_533/CLK sky130_fd_sc_hd__nor2b_1_152/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_186 sky130_fd_sc_hd__xor2_1_186/B sky130_fd_sc_hd__inv_2_19/A
+ sky130_fd_sc_hd__inv_2_11/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_537 wbs_dat_o[16] sky130_fd_sc_hd__dfxtp_1_538/CLK sky130_fd_sc_hd__nor2b_1_141/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_197 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__nor2_4_9/B
+ sky130_fd_sc_hd__xor2_1_197/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_548 wbs_dat_o[27] sky130_fd_sc_hd__dfxtp_1_552/CLK sky130_fd_sc_hd__nor2b_1_130/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_102 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_51/A1 sky130_fd_sc_hd__clkbuf_1_102/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_113 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_113/X sky130_fd_sc_hd__clkinv_1_976/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_124 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_124/X sky130_fd_sc_hd__buf_2_133/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_135 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_197/A sky130_fd_sc_hd__buf_6_19/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_206 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__buf_8_0/X sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__buf_4_6/X
+ sky130_fd_sc_hd__o21ai_1_378/B1 sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_146 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_27/A1 sky130_fd_sc_hd__clkbuf_1_146/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_217 vccd1 vssd1 sky130_fd_sc_hd__and3_4_15/X sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__nor2_1_87/A sky130_fd_sc_hd__nor2_1_130/Y sky130_fd_sc_hd__and2_0_49/A
+ sky130_fd_sc_hd__o21ai_1_406/B1 sky130_fd_sc_hd__nor2b_1_11/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_157 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_55/A1 sky130_fd_sc_hd__clkbuf_1_157/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_4 sky130_fd_sc_hd__dfxtp_1_4/Q sky130_fd_sc_hd__dfxtp_1_8/CLK
+ sky130_fd_sc_hd__dfxtp_1_4/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a222oi_1_228 vccd1 vssd1 sky130_fd_sc_hd__and3_4_11/X sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__or2_0_60/B sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__or2_0_60/A
+ sky130_fd_sc_hd__o21ai_1_419/B1 sky130_fd_sc_hd__and2b_4_8/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_168 vssd1 vccd1 sky130_fd_sc_hd__buf_8_40/A sky130_fd_sc_hd__inv_2_150/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o21ai_1_860 vssd1 vccd1 sky130_fd_sc_hd__nand2_2_13/Y sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__a22oi_1_222/Y sky130_fd_sc_hd__xor2_1_635/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_239 vccd1 vssd1 sky130_fd_sc_hd__and3_4_10/X sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__buf_4_2/X sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__o21ai_1_433/B1 sky130_fd_sc_hd__and2b_4_7/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_179 vssd1 vccd1 sky130_fd_sc_hd__a22o_1_24/B2 sky130_fd_sc_hd__clkbuf_1_179/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o21ai_1_871 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_649/A sky130_fd_sc_hd__nor2_1_230/Y
+ sky130_fd_sc_hd__nand2_1_701/Y sky130_fd_sc_hd__xnor2_1_197/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_882 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_662/A sky130_fd_sc_hd__nor2_1_247/Y
+ sky130_fd_sc_hd__nand2_1_776/Y sky130_fd_sc_hd__xnor2_1_214/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_409 sky130_fd_sc_hd__nor2_1_209/A sky130_fd_sc_hd__nor2_1_211/B
+ sky130_fd_sc_hd__fa_2_409/A sky130_fd_sc_hd__fa_2_409/B sky130_fd_sc_hd__xor2_1_617/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o21ai_1_893 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_676/A sky130_fd_sc_hd__nor2_1_254/Y
+ sky130_fd_sc_hd__nand2_1_793/Y sky130_fd_sc_hd__xnor2_1_290/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__inv_4_14 sky130_fd_sc_hd__inv_4_14/Y sky130_fd_sc_hd__inv_4_14/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__and2_0_100 vccd1 vssd1 sky130_fd_sc_hd__and2_0_100/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__or2_0_9/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_111 vccd1 vssd1 sky130_fd_sc_hd__and2_0_111/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_111/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_122 vccd1 vssd1 sky130_fd_sc_hd__and2_0_122/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_122/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_30 la_data_out[97] sky130_fd_sc_hd__conb_1_112/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_8_2 sky130_fd_sc_hd__nand2_8_2/A sky130_fd_sc_hd__nand2_8_2/B
+ sky130_fd_sc_hd__nor2_1_85/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_8
Xsky130_fd_sc_hd__and2_0_133 vccd1 vssd1 sky130_fd_sc_hd__and2_0_133/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_133/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_41 la_data_out[22] sky130_fd_sc_hd__conb_1_101/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_144 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_71/D sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_144/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_52 la_data_out[11] sky130_fd_sc_hd__conb_1_90/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_155 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_73/D sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_155/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_63 la_data_out[0] sky130_fd_sc_hd__conb_1_79/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_166 vccd1 vssd1 sky130_fd_sc_hd__and2_0_166/X sky130_fd_sc_hd__o21ai_2_0/B1
+ sky130_fd_sc_hd__and2_0_166/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_74 io_out[27] sky130_fd_sc_hd__conb_1_68/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_177 vccd1 vssd1 sky130_fd_sc_hd__and2_0_177/X sky130_fd_sc_hd__o21ai_2_0/B1
+ sky130_fd_sc_hd__and2_0_177/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_85 io_out[16] sky130_fd_sc_hd__conb_1_57/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_188 vccd1 vssd1 sky130_fd_sc_hd__and2_0_188/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_92/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_96 io_out[5] sky130_fd_sc_hd__conb_1_46/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_199 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_50/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_83/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o21ai_1_101 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_99/A2 sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__a22oi_1_161/Y sky130_fd_sc_hd__and2_0_176/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_112 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_113/A2 sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__a22oi_1_166/Y sky130_fd_sc_hd__and2_0_163/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_123 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_125/A2 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_129/Y sky130_fd_sc_hd__and2_0_149/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_134 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_137/A2 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_134/Y sky130_fd_sc_hd__and2_0_135/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_145 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_145/A2 sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__a22oi_1_183/Y sky130_fd_sc_hd__and2_0_122/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_156 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_157/A2 sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__a22oi_1_188/Y sky130_fd_sc_hd__and2_0_108/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_167 vssd1 vccd1 sky130_fd_sc_hd__inv_2_14/Y sky130_fd_sc_hd__nand2b_2_0/Y
+ sky130_fd_sc_hd__a222oi_1_49/Y sky130_fd_sc_hd__xor2_1_1/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_178 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_2/X sky130_fd_sc_hd__or2_0_5/X
+ sky130_fd_sc_hd__o21a_1_0/X sky130_fd_sc_hd__xnor2_1_6/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_189 vssd1 vccd1 sky130_fd_sc_hd__inv_2_10/Y sky130_fd_sc_hd__nand2b_2_0/Y
+ sky130_fd_sc_hd__a222oi_1_66/Y sky130_fd_sc_hd__xor2_1_18/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nand2_1_505 sky130_fd_sc_hd__nand2_1_602/B sky130_fd_sc_hd__nor2_1_196/A
+ sky130_fd_sc_hd__fah_1_9/SUM vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_516 sky130_fd_sc_hd__nand2_1_516/Y sky130_fd_sc_hd__or2_0_9/A
+ sky130_fd_sc_hd__or2_0_9/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_527 sky130_fd_sc_hd__xor2_1_468/B sky130_fd_sc_hd__o21ai_2_12/B1
+ sky130_fd_sc_hd__nand2_1_527/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_538 sky130_fd_sc_hd__xor2_1_489/B sky130_fd_sc_hd__o21ai_2_13/B1
+ sky130_fd_sc_hd__nand2_1_538/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_549 sky130_fd_sc_hd__xor2_1_509/B sky130_fd_sc_hd__nand2_1_550/Y
+ sky130_fd_sc_hd__nand2_1_549/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_7 sky130_fd_sc_hd__xnor2_1_71/Y sky130_fd_sc_hd__nor2b_1_7/Y
+ sky130_fd_sc_hd__nor2b_1_7/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1107 sky130_fd_sc_hd__clkinv_4_50/A sky130_fd_sc_hd__a22o_1_27/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1118 sky130_fd_sc_hd__clkinv_4_61/A sky130_fd_sc_hd__a22o_1_38/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1129 sky130_fd_sc_hd__clkinv_4_72/A sky130_fd_sc_hd__a22o_1_49/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_90 sky130_fd_sc_hd__nand2_1_90/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__xnor2_1_73/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_301 sky130_fd_sc_hd__dfxtp_1_301/Q sky130_fd_sc_hd__clkinv_8_6/Y
+ sky130_fd_sc_hd__and2_0_277/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1609 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_312 sky130_fd_sc_hd__nor2_1_240/A sky130_fd_sc_hd__dfxtp_1_319/CLK
+ sky130_fd_sc_hd__and2_0_289/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_323 sky130_fd_sc_hd__nor2_1_234/A sky130_fd_sc_hd__dfxtp_1_323/CLK
+ sky130_fd_sc_hd__and2_0_300/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_334 sky130_fd_sc_hd__dfxtp_1_334/Q sky130_fd_sc_hd__dfxtp_1_339/CLK
+ sky130_fd_sc_hd__and2_0_327/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_345 sky130_fd_sc_hd__dfxtp_1_345/Q sky130_fd_sc_hd__dfxtp_1_356/CLK
+ sky130_fd_sc_hd__and2_0_312/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_356 sky130_fd_sc_hd__dfxtp_1_356/Q sky130_fd_sc_hd__dfxtp_1_356/CLK
+ sky130_fd_sc_hd__and2_0_305/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_367 sky130_fd_sc_hd__dfxtp_1_367/Q sky130_fd_sc_hd__dfxtp_1_371/CLK
+ sky130_fd_sc_hd__nor2b_1_116/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_378 sky130_fd_sc_hd__dfxtp_1_378/Q sky130_fd_sc_hd__dfxtp_1_380/CLK
+ sky130_fd_sc_hd__nor2b_1_105/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_389 sky130_fd_sc_hd__dfxtp_1_389/Q sky130_fd_sc_hd__dfxtp_1_395/CLK
+ sky130_fd_sc_hd__nor2b_1_94/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_9 sky130_fd_sc_hd__nand2_1_9/Y sky130_fd_sc_hd__nand2_1_9/B
+ sky130_fd_sc_hd__nand2_1_9/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__fa_2_206 sky130_fd_sc_hd__fa_2_200/CIN sky130_fd_sc_hd__fa_2_203/B
+ sky130_fd_sc_hd__fa_2_206/A sky130_fd_sc_hd__fa_2_206/B sky130_fd_sc_hd__xor2_1_303/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o21ai_1_690 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_751/A2 sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__o21ai_1_690/B1 sky130_fd_sc_hd__xor2_1_470/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_217 sky130_fd_sc_hd__fa_2_214/CIN sky130_fd_sc_hd__fa_2_220/A
+ sky130_fd_sc_hd__fa_2_217/A sky130_fd_sc_hd__fa_2_217/B sky130_fd_sc_hd__xor2_1_316/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_228 sky130_fd_sc_hd__nor2_1_124/A sky130_fd_sc_hd__or2_0_34/B
+ sky130_fd_sc_hd__fa_2_228/A sky130_fd_sc_hd__fa_2_228/B sky130_fd_sc_hd__fa_2_228/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_239 sky130_fd_sc_hd__fa_2_232/CIN sky130_fd_sc_hd__fa_2_236/A
+ sky130_fd_sc_hd__fa_2_239/A sky130_fd_sc_hd__fa_2_239/B sky130_fd_sc_hd__xor2_1_343/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_20 sky130_fd_sc_hd__fa_2_16/B sky130_fd_sc_hd__fa_2_26/B sky130_fd_sc_hd__fa_2_20/A
+ sky130_fd_sc_hd__fa_2_20/B sky130_fd_sc_hd__xor2_1_32/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_31 sky130_fd_sc_hd__fa_2_24/A sky130_fd_sc_hd__fa_2_32/B sky130_fd_sc_hd__fa_2_31/A
+ sky130_fd_sc_hd__fa_2_31/B sky130_fd_sc_hd__xor2_1_51/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_42 sky130_fd_sc_hd__fa_2_35/A sky130_fd_sc_hd__fa_2_43/A sky130_fd_sc_hd__fa_2_42/A
+ sky130_fd_sc_hd__fa_2_42/B sky130_fd_sc_hd__fa_2_42/CIN vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_53 sky130_fd_sc_hd__fa_2_46/CIN sky130_fd_sc_hd__fa_2_52/A
+ sky130_fd_sc_hd__fa_2_53/A sky130_fd_sc_hd__fa_2_53/B sky130_fd_sc_hd__xor2_1_80/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_64 sky130_fd_sc_hd__fa_2_58/CIN sky130_fd_sc_hd__fa_2_61/B
+ sky130_fd_sc_hd__fa_2_64/A sky130_fd_sc_hd__fa_2_64/B sky130_fd_sc_hd__xor2_1_90/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_75 sky130_fd_sc_hd__fa_2_72/CIN sky130_fd_sc_hd__fa_2_78/A
+ sky130_fd_sc_hd__fa_2_75/A sky130_fd_sc_hd__fa_2_75/B sky130_fd_sc_hd__fa_2_75/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_86 sky130_fd_sc_hd__nor2_1_65/A sky130_fd_sc_hd__or2_0_7/B
+ sky130_fd_sc_hd__fa_2_86/A sky130_fd_sc_hd__fa_2_86/B sky130_fd_sc_hd__fa_2_86/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_97 sky130_fd_sc_hd__fa_2_90/CIN sky130_fd_sc_hd__fa_2_94/A
+ sky130_fd_sc_hd__fa_2_97/A sky130_fd_sc_hd__fa_2_97/B sky130_fd_sc_hd__fa_2_97/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_201 vccd1 vssd1 la_data_out[87] sky130_fd_sc_hd__nand2_2_6/Y
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_212 vccd1 vssd1 la_data_out[69] sky130_fd_sc_hd__or2_0_82/B
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__or3_1_0 wbs_adr_i[4] sky130_fd_sc_hd__or3_1_0/X wbs_adr_i[3] wbs_adr_i[2]
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__or3_1
Xsky130_fd_sc_hd__a21oi_1_14 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_43/Y
+ sky130_fd_sc_hd__a21oi_1_14/Y sky130_fd_sc_hd__dfxtp_1_83/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_25 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_54/Y
+ sky130_fd_sc_hd__a21oi_1_25/Y sky130_fd_sc_hd__dfxtp_1_72/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_570 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_400/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_432/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_767/A sky130_fd_sc_hd__dfxtp_1_368/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a21oi_1_36 sky130_fd_sc_hd__inv_2_11/A sky130_fd_sc_hd__o21ai_1_314/Y
+ sky130_fd_sc_hd__xnor2_1_0/A sky130_fd_sc_hd__nor2_1_74/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_581 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_412/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_444/Q sky130_fd_sc_hd__clkbuf_1_32/X
+ sky130_fd_sc_hd__clkinv_1_778/A sky130_fd_sc_hd__dfxtp_1_380/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a21oi_1_47 sky130_fd_sc_hd__o21ai_1_281/Y sky130_fd_sc_hd__nor2_1_63/A
+ sky130_fd_sc_hd__a21oi_1_47/Y sky130_fd_sc_hd__or2_0_17/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_592 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_400/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_432/Q sky130_fd_sc_hd__clkbuf_1_32/X
+ sky130_fd_sc_hd__clkinv_1_789/A sky130_fd_sc_hd__dfxtp_1_368/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a21oi_1_58 sky130_fd_sc_hd__nand2_1_272/Y sky130_fd_sc_hd__a21oi_1_58/B1
+ sky130_fd_sc_hd__a21oi_1_58/Y sky130_fd_sc_hd__nand2_1_273/A vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_69 sky130_fd_sc_hd__xnor2_2_1/B sky130_fd_sc_hd__a21oi_1_69/B1
+ sky130_fd_sc_hd__a21oi_1_69/Y sky130_fd_sc_hd__or2_0_27/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__decap_12_10 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_21 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_32 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_43 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_54 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_65 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_76 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_87 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_98 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_10 vccd1 vssd1 sky130_fd_sc_hd__buf_6_10/X sky130_fd_sc_hd__buf_6_9/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_21 vccd1 vssd1 sky130_fd_sc_hd__buf_6_21/X sky130_fd_sc_hd__inv_12_1/Y
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_32 vccd1 vssd1 sky130_fd_sc_hd__buf_6_32/X sky130_fd_sc_hd__buf_8_66/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_43 vccd1 vssd1 sky130_fd_sc_hd__buf_6_43/X sky130_fd_sc_hd__buf_8_94/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_54 vccd1 vssd1 sky130_fd_sc_hd__buf_6_54/X sky130_fd_sc_hd__buf_8_85/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_65 vccd1 vssd1 sky130_fd_sc_hd__buf_6_65/X sky130_fd_sc_hd__buf_8_81/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_76 vccd1 vssd1 sky130_fd_sc_hd__buf_6_76/X sky130_fd_sc_hd__buf_6_76/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_87 vccd1 vssd1 sky130_fd_sc_hd__buf_6_87/X sky130_fd_sc_hd__inv_16_4/Y
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_12 la_data_out[62] vssd1 vccd1 vccd1 vssd1 sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_23 sky130_fd_sc_hd__clkinv_4_61/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_34 sky130_fd_sc_hd__clkinv_4_46/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_45 sky130_fd_sc_hd__buf_2_189/A vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_56 sky130_fd_sc_hd__buf_2_192/A vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_67 la_data_out[62] vssd1 vccd1 vccd1 vssd1 sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__decap_12_407 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_418 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_302 sky130_fd_sc_hd__xnor2_1_56/A sky130_fd_sc_hd__nand2_1_303/Y
+ sky130_fd_sc_hd__nand2_1_302/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_429 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_901 sky130_fd_sc_hd__clkinv_1_901/Y sky130_fd_sc_hd__clkinv_1_901/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_313 sky130_fd_sc_hd__xor2_1_207/A sky130_fd_sc_hd__nand2_1_314/Y
+ sky130_fd_sc_hd__nand2_1_313/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_912 sky130_fd_sc_hd__clkinv_1_912/Y sky130_fd_sc_hd__inv_2_107/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_324 sky130_fd_sc_hd__nand2_1_324/Y sky130_fd_sc_hd__nor2_1_121/Y
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_923 sky130_fd_sc_hd__inv_2_111/A sky130_fd_sc_hd__inv_4_10/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_335 sky130_fd_sc_hd__nor2_1_107/A sky130_fd_sc_hd__or2_0_36/X
+ sky130_fd_sc_hd__or2_0_38/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_934 sky130_fd_sc_hd__inv_2_124/A sky130_fd_sc_hd__buf_2_54/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_346 sky130_fd_sc_hd__nand2_1_346/Y sky130_fd_sc_hd__nor2_1_112/Y
+ sky130_fd_sc_hd__nand2_1_374/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_945 sky130_fd_sc_hd__buf_8_86/A sky130_fd_sc_hd__inv_2_141/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_357 sky130_fd_sc_hd__nand2_1_357/Y sky130_fd_sc_hd__nor2_1_115/Y
+ sky130_fd_sc_hd__nand2_1_374/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_956 sky130_fd_sc_hd__clkinv_1_956/Y sky130_fd_sc_hd__inv_2_151/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_368 sky130_fd_sc_hd__nand2_1_368/Y sky130_fd_sc_hd__nand2_1_368/B
+ sky130_fd_sc_hd__nand2_1_374/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_967 sky130_fd_sc_hd__clkinv_1_967/Y sky130_fd_sc_hd__clkinv_2_32/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_379 sky130_fd_sc_hd__or2_0_32/B sky130_fd_sc_hd__nor2_1_123/Y
+ sky130_fd_sc_hd__nor2_1_128/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_978 sky130_fd_sc_hd__clkinv_1_978/Y sky130_fd_sc_hd__clkinv_4_26/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_989 sky130_fd_sc_hd__clkinv_1_989/Y sky130_fd_sc_hd__clkinv_2_35/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1406 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1417 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_120 sky130_fd_sc_hd__dfxtp_1_120/Q sky130_fd_sc_hd__dfxtp_1_122/CLK
+ sky130_fd_sc_hd__and2_0_228/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1428 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_131 sky130_fd_sc_hd__dfxtp_1_131/Q sky130_fd_sc_hd__dfxtp_1_138/CLK
+ sky130_fd_sc_hd__and2_0_126/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1439 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_142 sky130_fd_sc_hd__dfxtp_1_142/Q sky130_fd_sc_hd__dfxtp_1_146/CLK
+ sky130_fd_sc_hd__and2_0_185/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_153 sky130_fd_sc_hd__dfxtp_1_153/Q sky130_fd_sc_hd__dfxtp_1_154/CLK
+ sky130_fd_sc_hd__and2_0_236/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_164 sky130_fd_sc_hd__dfxtp_1_164/Q sky130_fd_sc_hd__dfxtp_1_170/CLK
+ sky130_fd_sc_hd__and2_0_128/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_175 sky130_fd_sc_hd__dfxtp_1_175/Q sky130_fd_sc_hd__dfxtp_1_176/CLK
+ sky130_fd_sc_hd__and2_0_172/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_186 sky130_fd_sc_hd__dfxtp_1_186/Q sky130_fd_sc_hd__dfxtp_1_190/CLK
+ sky130_fd_sc_hd__and2_0_237/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_197 sky130_fd_sc_hd__xnor2_1_176/A sky130_fd_sc_hd__dfxtp_2_1/CLK
+ sky130_fd_sc_hd__and2_0_55/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_930 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_941 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_952 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_963 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_974 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_985 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_996 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o211ai_1_17 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_46/B1
+ sky130_fd_sc_hd__o211ai_1_17/Y sky130_fd_sc_hd__a22oi_1_66/Y sky130_fd_sc_hd__a22oi_1_67/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_28 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_33/B1
+ sky130_fd_sc_hd__o211ai_1_28/Y sky130_fd_sc_hd__a22oi_1_88/Y sky130_fd_sc_hd__a22oi_1_89/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_39 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o21ai_1_9/A2
+ sky130_fd_sc_hd__xor3_1_25/A sky130_fd_sc_hd__nand2_1_59/Y sky130_fd_sc_hd__a21oi_1_10/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o21ai_1_80 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_81/A2 sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_80/B1 sky130_fd_sc_hd__o21ai_1_80/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_91 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_93/A2 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__o21ai_1_91/B1 sky130_fd_sc_hd__o21ai_1_91/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkinv_1_208 sky130_fd_sc_hd__o22ai_1_51/B1 sky130_fd_sc_hd__dfxtp_1_171/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_219 sky130_fd_sc_hd__o22ai_1_9/B1 sky130_fd_sc_hd__dfxtp_1_104/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_2_8 sky130_fd_sc_hd__o21ai_2_8/B1 sky130_fd_sc_hd__o21ai_2_8/Y
+ sky130_fd_sc_hd__a21oi_2_5/Y sky130_fd_sc_hd__nor2_1_69/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__o21ai_2
Xsky130_fd_sc_hd__a21oi_1_105 sky130_fd_sc_hd__nand2_1_503/Y sky130_fd_sc_hd__nand2_1_643/Y
+ sky130_fd_sc_hd__o21ai_2_17/A2 sky130_fd_sc_hd__nor2_1_215/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_116 sky130_fd_sc_hd__nand2_1_572/Y sky130_fd_sc_hd__o21ai_1_735/Y
+ sky130_fd_sc_hd__o21a_1_4/A2 sky130_fd_sc_hd__nor2_1_180/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_127 sky130_fd_sc_hd__nor2_1_197/Y sky130_fd_sc_hd__nand2_1_603/Y
+ sky130_fd_sc_hd__a21oi_1_127/Y sky130_fd_sc_hd__nand2_1_614/Y vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_138 sky130_fd_sc_hd__xnor2_1_188/B sky130_fd_sc_hd__clkinv_1_625/Y
+ sky130_fd_sc_hd__a21oi_1_138/Y sky130_fd_sc_hd__or2_0_73/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_149 sky130_fd_sc_hd__xnor2_1_199/B sky130_fd_sc_hd__clkinv_1_647/Y
+ sky130_fd_sc_hd__xor2_1_650/A sky130_fd_sc_hd__or2_0_82/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_520 sky130_fd_sc_hd__buf_12_520/A sky130_fd_sc_hd__buf_12_520/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_531 sky130_fd_sc_hd__buf_12_531/A sky130_fd_sc_hd__buf_12_531/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_542 sky130_fd_sc_hd__buf_12_542/A sky130_fd_sc_hd__buf_12_542/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_553 sky130_fd_sc_hd__buf_12_553/A sky130_fd_sc_hd__buf_12_553/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_564 sky130_fd_sc_hd__buf_12_564/A sky130_fd_sc_hd__buf_12_564/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_8_1 sky130_fd_sc_hd__buf_6_23/A sky130_fd_sc_hd__clkbuf_8_1/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_8
Xsky130_fd_sc_hd__buf_12_575 sky130_fd_sc_hd__buf_12_575/A sky130_fd_sc_hd__buf_12_575/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_204 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_586 sky130_fd_sc_hd__buf_12_586/A sky130_fd_sc_hd__buf_12_586/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_215 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_597 sky130_fd_sc_hd__buf_12_597/A sky130_fd_sc_hd__buf_12_597/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_226 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_110 sky130_fd_sc_hd__o21ai_1_86/B1 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__xnor2_1_95/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_237 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_121 sky130_fd_sc_hd__nand2_1_121/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__xnor2_1_104/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_248 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_720 sky130_fd_sc_hd__nor2b_1_99/A sky130_fd_sc_hd__xnor2_1_293/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_132 sky130_fd_sc_hd__nand2_1_132/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_133/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_259 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_731 sky130_fd_sc_hd__nor2b_1_110/A sky130_fd_sc_hd__xor2_1_684/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_143 sky130_fd_sc_hd__nand2_1_143/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__xor2_1_419/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_742 sky130_fd_sc_hd__fa_2_463/A sky130_fd_sc_hd__clkinv_1_742/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_305 vssd1 vccd1 sky130_fd_sc_hd__ha_2_49/SUM sky130_fd_sc_hd__nand4_1_2/C
+ la_data_out[42] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_154 sky130_fd_sc_hd__nand2_1_154/Y sky130_fd_sc_hd__nor2_1_61/Y
+ sky130_fd_sc_hd__clkbuf_1_3/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_753 sky130_fd_sc_hd__fa_2_476/A sky130_fd_sc_hd__clkinv_1_753/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_165 sky130_fd_sc_hd__xnor2_1_6/A sky130_fd_sc_hd__nand2_1_166/Y
+ sky130_fd_sc_hd__or2_0_4/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_764 sky130_fd_sc_hd__fa_2_487/A sky130_fd_sc_hd__clkinv_1_764/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_176 sky130_fd_sc_hd__nor2_1_50/A sky130_fd_sc_hd__or2_0_12/X
+ sky130_fd_sc_hd__nand2_1_188/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_775 sky130_fd_sc_hd__and2_0_332/A sky130_fd_sc_hd__clkinv_1_775/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_187 sky130_fd_sc_hd__nor2_1_54/A sky130_fd_sc_hd__nand2_1_199/A
+ sky130_fd_sc_hd__or2_0_15/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_786 sky130_fd_sc_hd__and2_0_321/A sky130_fd_sc_hd__clkinv_1_786/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_198 sky130_fd_sc_hd__nor2_1_57/B sky130_fd_sc_hd__or2_0_14/X
+ sky130_fd_sc_hd__or2_0_13/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_797 sky130_fd_sc_hd__and2_0_310/A sky130_fd_sc_hd__clkinv_1_797/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1203 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_3 sky130_fd_sc_hd__fa_2_28/A sky130_fd_sc_hd__xor3_1_4/B
+ sky130_fd_sc_hd__xor2_1_3/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1214 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1225 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1236 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1247 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1258 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1269 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_8_1 sky130_fd_sc_hd__clkinv_8_1/Y sky130_fd_sc_hd__clkinv_8_1/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__xor2_1_18 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__fa_2_3/CIN
+ sky130_fd_sc_hd__xor2_1_18/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_29 sky130_fd_sc_hd__xor2_1_9/B sky130_fd_sc_hd__xor2_1_29/X
+ sky130_fd_sc_hd__xor2_1_29/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_760 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_771 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_782 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_793 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_505 sky130_fd_sc_hd__fah_1_14/A sky130_fd_sc_hd__fa_2_339/A
+ sky130_fd_sc_hd__xor2_1_505/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_516 sky130_fd_sc_hd__fa_2_357/A sky130_fd_sc_hd__xor2_1_516/X
+ sky130_fd_sc_hd__xor2_1_516/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_527 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__xor2_1_527/X
+ sky130_fd_sc_hd__xor2_1_527/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_538 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__fa_2_365/A
+ sky130_fd_sc_hd__xor2_1_538/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_549 sky130_fd_sc_hd__fa_2_379/A sky130_fd_sc_hd__fa_2_372/B
+ sky130_fd_sc_hd__xor2_1_549/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1770 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1781 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_80 la_data_out[46] sky130_fd_sc_hd__inv_2_81/A vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1792 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_91 sky130_fd_sc_hd__inv_2_92/A sky130_fd_sc_hd__inv_2_91/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__ha_2_12 vssd1 vccd1 sky130_fd_sc_hd__ha_2_12/A sky130_fd_sc_hd__fa_2_433/A
+ sky130_fd_sc_hd__fa_2_435/B sky130_fd_sc_hd__ha_2_12/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_23 vssd1 vccd1 sky130_fd_sc_hd__ha_2_23/A sky130_fd_sc_hd__ha_2_22/B
+ sky130_fd_sc_hd__ha_2_23/SUM sky130_fd_sc_hd__ha_2_23/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_34 vssd1 vccd1 sky130_fd_sc_hd__ha_2_34/A sky130_fd_sc_hd__ha_2_33/B
+ sky130_fd_sc_hd__ha_2_34/SUM sky130_fd_sc_hd__ha_2_34/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_45 vssd1 vccd1 sky130_fd_sc_hd__ha_2_45/A sky130_fd_sc_hd__ha_2_44/B
+ sky130_fd_sc_hd__ha_2_45/SUM sky130_fd_sc_hd__ha_2_45/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__and2b_4_7 sky130_fd_sc_hd__nor2_4_12/A sky130_fd_sc_hd__and2b_4_7/X
+ sky130_fd_sc_hd__and3_4_10/C vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__and2b_4
Xsky130_fd_sc_hd__ha_2_56 vssd1 vccd1 sky130_fd_sc_hd__ha_2_56/A sky130_fd_sc_hd__ha_2_55/B
+ sky130_fd_sc_hd__maj3_1_3/A sky130_fd_sc_hd__ha_2_56/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__sdlclkp_4_30 sky130_fd_sc_hd__conb_1_144/LO sky130_fd_sc_hd__clkinv_4_99/Y
+ sky130_fd_sc_hd__dfxtp_1_323/CLK sky130_fd_sc_hd__nand2_1_713/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__clkbuf_1_8 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_548/B sky130_fd_sc_hd__fa_2_389/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__sdlclkp_4_41 sky130_fd_sc_hd__conb_1_145/LO sky130_fd_sc_hd__clkinv_4_11/Y
+ sky130_fd_sc_hd__dfxtp_1_410/CLK sky130_fd_sc_hd__o21ai_1_891/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_52 sky130_fd_sc_hd__conb_1_149/LO sky130_fd_sc_hd__clkinv_4_119/A
+ sky130_fd_sc_hd__dfxtp_1_538/CLK sky130_fd_sc_hd__or2_0_113/X vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_110 sky130_fd_sc_hd__nor2_1_110/B sky130_fd_sc_hd__nor2_1_110/Y
+ sky130_fd_sc_hd__nor2_1_110/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_121 sky130_fd_sc_hd__and3_4_13/A sky130_fd_sc_hd__nor2_1_121/Y
+ sky130_fd_sc_hd__and3_4_13/C vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_132 sky130_fd_sc_hd__nor2_1_132/B sky130_fd_sc_hd__nor2_1_132/Y
+ sky130_fd_sc_hd__nor2_1_132/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_143 sky130_fd_sc_hd__nor2_1_148/Y sky130_fd_sc_hd__nor2_1_143/Y
+ sky130_fd_sc_hd__nor2_1_146/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_154 sky130_fd_sc_hd__nor2_1_154/B sky130_fd_sc_hd__nor2_1_154/Y
+ sky130_fd_sc_hd__nor2_1_154/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_30 sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__dfxtp_1_276/Q sky130_fd_sc_hd__o211ai_1_0/Y sky130_fd_sc_hd__nand2_2_7/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_8 la_data_out[119] sky130_fd_sc_hd__clkinv_1_8/A vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_165 sky130_fd_sc_hd__nor2_1_169/A sky130_fd_sc_hd__nor2_1_165/Y
+ sky130_fd_sc_hd__nor2_1_165/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_41 sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__dfxtp_1_99/Q sky130_fd_sc_hd__dfxtp_1_67/Q sky130_fd_sc_hd__a22oi_1_41/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_176 sky130_fd_sc_hd__nor2_1_176/B sky130_fd_sc_hd__nor2_1_176/Y
+ sky130_fd_sc_hd__nor2_1_176/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_52 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__nor2_4_3/Y
+ sky130_fd_sc_hd__nand2_1_73/B sky130_fd_sc_hd__dfxtp_1_137/Q sky130_fd_sc_hd__a22oi_1_52/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_187 sky130_fd_sc_hd__nor2_1_73/B sky130_fd_sc_hd__nor2_1_187/Y
+ sky130_fd_sc_hd__buf_6_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_63 sky130_fd_sc_hd__clkbuf_1_24/X sky130_fd_sc_hd__clkbuf_1_23/X
+ sky130_fd_sc_hd__dfxtp_1_110/Q sky130_fd_sc_hd__dfxtp_1_78/Q sky130_fd_sc_hd__a22oi_1_63/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_198 sky130_fd_sc_hd__nor2_1_85/B sky130_fd_sc_hd__nor2_1_198/Y
+ sky130_fd_sc_hd__nor2_1_87/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_74 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__nor2_4_3/Y
+ sky130_fd_sc_hd__nand2_1_62/B sky130_fd_sc_hd__dfxtp_1_148/Q sky130_fd_sc_hd__a22oi_1_74/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_85 sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__dfxtp_1_121/Q sky130_fd_sc_hd__dfxtp_1_89/Q sky130_fd_sc_hd__a22oi_1_85/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_96 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_188/Q sky130_fd_sc_hd__dfxtp_1_156/Q sky130_fd_sc_hd__o21ai_1_2/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_350 sky130_fd_sc_hd__buf_12_36/X sky130_fd_sc_hd__buf_12_617/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_361 sky130_fd_sc_hd__buf_12_48/X sky130_fd_sc_hd__buf_12_662/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_220 sky130_fd_sc_hd__or2_0_72/B sky130_fd_sc_hd__or2_0_72/A
+ sky130_fd_sc_hd__nor2b_2_5/Y sky130_fd_sc_hd__nor2_2_32/Y sky130_fd_sc_hd__a22oi_1_220/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_372 sky130_fd_sc_hd__buf_12_69/X sky130_fd_sc_hd__buf_12_472/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_383 sky130_fd_sc_hd__buf_12_383/A sky130_fd_sc_hd__buf_12_499/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_394 sky130_fd_sc_hd__buf_12_394/A sky130_fd_sc_hd__buf_12_540/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xnor2_1_102 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_102/B sky130_fd_sc_hd__inv_2_35/A
+ sky130_fd_sc_hd__xnor2_1_102/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_550 sky130_fd_sc_hd__nand2_1_546/A sky130_fd_sc_hd__or2_0_55/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_113 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_113/B sky130_fd_sc_hd__xnor2_1_113/Y
+ sky130_fd_sc_hd__xnor2_1_113/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_561 sky130_fd_sc_hd__o21ai_1_752/A1 sky130_fd_sc_hd__nor2_1_182/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_124 vssd1 vccd1 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__nor2_4_14/A
+ sky130_fd_sc_hd__xnor2_1_124/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_572 sky130_fd_sc_hd__nand2_1_579/A sky130_fd_sc_hd__nor2_2_27/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_135 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_135/B sky130_fd_sc_hd__xnor2_1_135/Y
+ sky130_fd_sc_hd__xnor2_1_135/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_583 sky130_fd_sc_hd__nand2_1_605/A sky130_fd_sc_hd__nor2_1_198/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_146 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_146/B sky130_fd_sc_hd__xnor2_1_146/Y
+ sky130_fd_sc_hd__xnor2_1_146/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_594 sky130_fd_sc_hd__nand2_1_621/A sky130_fd_sc_hd__nor2_1_206/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_157 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_557/A sky130_fd_sc_hd__and3_4_25/B
+ sky130_fd_sc_hd__xnor2_1_160/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_168 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_596/A sky130_fd_sc_hd__nor2b_2_5/A
+ sky130_fd_sc_hd__xnor2_1_171/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_4_30 sky130_fd_sc_hd__nand2_2_1/Y sky130_fd_sc_hd__inv_2_155/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__xnor2_1_179 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_179/B sky130_fd_sc_hd__xnor2_1_179/Y
+ sky130_fd_sc_hd__xnor2_1_179/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_4_41 sky130_fd_sc_hd__clkinv_8_25/A sky130_fd_sc_hd__clkinv_8_24/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_52 sky130_fd_sc_hd__clkinv_4_52/A sky130_fd_sc_hd__clkinv_4_52/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_63 sky130_fd_sc_hd__clkinv_4_63/A sky130_fd_sc_hd__clkinv_4_63/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_74 sky130_fd_sc_hd__clkinv_4_74/A sky130_fd_sc_hd__clkinv_4_74/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_1000 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_4_85 wbs_dat_i[21] sky130_fd_sc_hd__clkinv_4_85/Y vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_1011 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_4_96 sky130_fd_sc_hd__clkinv_8_47/Y sky130_fd_sc_hd__clkinv_8_48/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_1022 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1033 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1044 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1055 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1066 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_16_4 sky130_fd_sc_hd__inv_16_4/Y sky130_fd_sc_hd__inv_16_4/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__decap_12_1077 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_508 vssd1 vccd1 sky130_fd_sc_hd__inv_2_28/Y sky130_fd_sc_hd__nand2b_1_14/Y
+ sky130_fd_sc_hd__o21ai_1_508/B1 sky130_fd_sc_hd__xor2_1_307/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1088 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_519 vssd1 vccd1 sky130_fd_sc_hd__inv_2_32/Y sky130_fd_sc_hd__nand2b_2_3/Y
+ sky130_fd_sc_hd__o21ai_1_519/B1 sky130_fd_sc_hd__xor2_1_318/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1099 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__and2b_4_11 sky130_fd_sc_hd__nor2_4_16/A sky130_fd_sc_hd__and2b_4_11/X
+ sky130_fd_sc_hd__and3_4_20/C vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__and2b_4
Xsky130_fd_sc_hd__decap_12_590 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_302 sky130_fd_sc_hd__xor2_1_383/B sky130_fd_sc_hd__xor2_1_302/X
+ sky130_fd_sc_hd__xor2_1_302/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_313 sky130_fd_sc_hd__xor2_1_313/B sky130_fd_sc_hd__xor2_1_313/X
+ sky130_fd_sc_hd__xor2_1_313/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_324 sky130_fd_sc_hd__fa_2_262/A sky130_fd_sc_hd__fa_2_225/B
+ sky130_fd_sc_hd__xor2_1_324/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_335 sky130_fd_sc_hd__fa_2_250/A sky130_fd_sc_hd__fa_2_233/B
+ sky130_fd_sc_hd__xor2_1_335/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_346 sky130_fd_sc_hd__xor2_1_346/B sky130_fd_sc_hd__xor2_1_346/X
+ sky130_fd_sc_hd__xor2_1_346/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_357 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__xor2_1_357/X
+ sky130_fd_sc_hd__xor2_1_357/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_368 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__fa_2_254/B
+ sky130_fd_sc_hd__xor2_1_368/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_379 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__fa_2_261/B
+ sky130_fd_sc_hd__xor2_1_379/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_306 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_306/X sky130_fd_sc_hd__buf_8_19/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_317 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_317/X sky130_fd_sc_hd__clkinv_1_878/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_328 vssd1 vccd1 la_data_out[49] sky130_fd_sc_hd__ha_2_39/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_339 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1_9/D sky130_fd_sc_hd__dfxtp_1_10/Q
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_10 sky130_fd_sc_hd__dfxtp_1_10/Q sky130_fd_sc_hd__dfxtp_1_8/CLK
+ la_data_out[61] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_21 sky130_fd_sc_hd__ha_2_5/A sky130_fd_sc_hd__dfxtp_1_29/CLK
+ sky130_fd_sc_hd__or4_1_3/B vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_32 sky130_fd_sc_hd__nand2_1_82/B sky130_fd_sc_hd__dfxtp_1_46/CLK
+ sky130_fd_sc_hd__dfxtp_1_32/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_43 sky130_fd_sc_hd__nand2_1_71/B sky130_fd_sc_hd__dfxtp_1_43/CLK
+ sky130_fd_sc_hd__dfxtp_1_43/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_54 sky130_fd_sc_hd__nand2_1_60/B sky130_fd_sc_hd__dfxtp_1_57/CLK
+ sky130_fd_sc_hd__dfxtp_1_54/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_65 sky130_fd_sc_hd__dfxtp_1_65/Q sky130_fd_sc_hd__dfxtp_1_65/CLK
+ sky130_fd_sc_hd__dfxtp_1_65/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_76 sky130_fd_sc_hd__dfxtp_1_76/Q sky130_fd_sc_hd__dfxtp_1_78/CLK
+ sky130_fd_sc_hd__dfxtp_1_76/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_87 sky130_fd_sc_hd__dfxtp_1_87/Q sky130_fd_sc_hd__dfxtp_1_89/CLK
+ sky130_fd_sc_hd__dfxtp_1_87/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_98 sky130_fd_sc_hd__dfxtp_1_98/Q sky130_fd_sc_hd__dfxtp_1_99/CLK
+ sky130_fd_sc_hd__dfxtp_1_98/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_304 vccd1 vssd1 sky130_fd_sc_hd__and2_0_304/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_304/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_315 vccd1 vssd1 sky130_fd_sc_hd__and2_0_315/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_315/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_326 vccd1 vssd1 sky130_fd_sc_hd__and2_0_326/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_326/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_337 vccd1 vssd1 sky130_fd_sc_hd__and2_0_396/A sky130_fd_sc_hd__ha_2_46/SUM
+ sky130_fd_sc_hd__and2_0_342/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_348 vccd1 vssd1 sky130_fd_sc_hd__and2_0_348/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__buf_2_41/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_359 vccd1 vssd1 sky130_fd_sc_hd__and2_0_359/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__buf_2_45/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__inv_2_104 sky130_fd_sc_hd__inv_4_21/Y sky130_fd_sc_hd__inv_2_104/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_115 sky130_fd_sc_hd__inv_2_115/A sky130_fd_sc_hd__buf_4_26/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__or2_0_6 sky130_fd_sc_hd__or2_0_6/A sky130_fd_sc_hd__or2_0_6/X sky130_fd_sc_hd__or2_0_6/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__inv_2_126 sky130_fd_sc_hd__inv_2_126/A sky130_fd_sc_hd__inv_2_126/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_137 sky130_fd_sc_hd__buf_8_5/A sky130_fd_sc_hd__inv_2_138/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_148 sky130_fd_sc_hd__inv_2_148/A sky130_fd_sc_hd__buf_8_34/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_159 sky130_fd_sc_hd__inv_2_159/A sky130_fd_sc_hd__buf_12_9/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_sram_1kbyte_1rw1r_32x256_8_0 sky130_fd_sc_hd__clkinv_2_30/Y sky130_fd_sc_hd__clkinv_2_30/Y
+ sky130_fd_sc_hd__buf_12_672/X sky130_fd_sc_hd__buf_12_617/X sky130_fd_sc_hd__buf_12_671/X
+ sky130_fd_sc_hd__buf_12_624/X sky130_fd_sc_hd__buf_12_378/X sky130_fd_sc_hd__buf_12_629/X
+ sky130_fd_sc_hd__buf_12_583/X sky130_fd_sc_hd__clkinv_2_32/Y sky130_fd_sc_hd__buf_12_576/X
+ sky130_fd_sc_hd__buf_12_567/X sky130_fd_sc_hd__buf_12_579/X vccd1 sky130_fd_sc_hd__clkinv_8_30/Y
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[16] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[17]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[18] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[19]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[20] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[21]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[22] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[23]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[24] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[25]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[26] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[27]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[28] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[29]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[30] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[31]
+ sky130_fd_sc_hd__buf_12_554/X sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[1] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[2]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[3] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[4]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[5] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[6]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[7] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[8]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[9] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[10]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[11] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[12]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[13] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[14]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[15] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout1[0]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[10] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[11]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[12] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[13]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[14] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[15]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[16] sky130_fd_sc_hd__buf_12_549/X sky130_fd_sc_hd__buf_12_307/X
+ sky130_fd_sc_hd__buf_12_127/X sky130_fd_sc_hd__buf_12_309/X sky130_fd_sc_hd__buf_12_164/X
+ sky130_fd_sc_hd__dfxtp_1_3/CLK sky130_fd_sc_hd__buf_6_9/X sky130_fd_sc_hd__buf_6_9/X
+ sky130_fd_sc_hd__buf_6_9/X sky130_fd_sc_hd__buf_6_9/X sky130_fd_sc_hd__buf_6_9/X
+ sky130_fd_sc_hd__buf_6_9/X sky130_fd_sc_hd__buf_6_9/X sky130_fd_sc_hd__buf_6_9/X
+ sky130_fd_sc_hd__buf_6_9/X sky130_fd_sc_hd__buf_6_9/X sky130_fd_sc_hd__buf_6_9/X
+ sky130_fd_sc_hd__buf_6_9/X sky130_fd_sc_hd__buf_6_10/X sky130_fd_sc_hd__buf_6_10/X
+ sky130_fd_sc_hd__buf_6_10/X sky130_fd_sc_hd__buf_6_10/X sky130_fd_sc_hd__buf_6_10/X
+ sky130_fd_sc_hd__buf_6_10/X sky130_fd_sc_hd__buf_6_10/X sky130_fd_sc_hd__buf_6_10/X
+ sky130_fd_sc_hd__buf_6_10/X sky130_fd_sc_hd__buf_6_10/X sky130_fd_sc_hd__buf_6_10/X
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[0] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[1]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[2] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[3]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[4] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[5]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[6] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[7]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[8] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[9]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[25] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[26]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[27] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[28]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[29] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[30]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[31] sky130_fd_sc_hd__clkbuf_4_22/X sky130_fd_sc_hd__buf_6_10/X
+ sky130_fd_sc_hd__buf_6_10/X sky130_fd_sc_hd__clkbuf_4_22/X sky130_fd_sc_hd__clkbuf_4_22/X
+ sky130_fd_sc_hd__clkbuf_4_22/X sky130_fd_sc_hd__clkbuf_4_22/X sky130_fd_sc_hd__clkbuf_4_22/X
+ sky130_fd_sc_hd__clkbuf_4_22/X sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[17] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[18]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[19] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[20]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[21] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[22]
+ sky130_fd_sc_hd__buf_12_569/X sky130_fd_sc_hd__buf_12_524/X sky130_fd_sc_hd__buf_12_197/X
+ sky130_fd_sc_hd__buf_12_464/X sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[23] sky130_sram_1kbyte_1rw1r_32x256_8_0/dout0[24]
+ sky130_sram_1kbyte_1rw1r_32x256_8_0/sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/gnd_uq26
+ vssd1 sky130_sram_1kbyte_1rw1r_32x256_8
Xsky130_fd_sc_hd__buf_12_180 sky130_fd_sc_hd__buf_8_106/X sky130_fd_sc_hd__buf_12_354/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_191 sky130_fd_sc_hd__buf_4_33/X sky130_fd_sc_hd__buf_12_322/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_380 sky130_fd_sc_hd__nand2_1_270/A sky130_fd_sc_hd__nor2_1_88/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_391 sky130_fd_sc_hd__nand2_1_289/A sky130_fd_sc_hd__nor2_1_98/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a211o_1_5 vssd1 vccd1 sky130_fd_sc_hd__fa_2_279/A sky130_fd_sc_hd__dfxtp_1_68/Q
+ sky130_fd_sc_hd__nor2_1_9/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_5/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__o21ai_1_305 vssd1 vccd1 sky130_fd_sc_hd__inv_2_20/Y sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__o21ai_1_305/B1 sky130_fd_sc_hd__xor2_1_125/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_316 vssd1 vccd1 sky130_fd_sc_hd__inv_2_9/Y sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__o21ai_1_316/B1 sky130_fd_sc_hd__xor2_1_136/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_327 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_327/A2 sky130_fd_sc_hd__nor2_2_10/Y
+ sky130_fd_sc_hd__nand2_1_253/Y sky130_fd_sc_hd__o21ai_1_327/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_338 vssd1 vccd1 sky130_fd_sc_hd__inv_2_11/Y sky130_fd_sc_hd__nand2_1_256/Y
+ sky130_fd_sc_hd__a21oi_1_54/Y sky130_fd_sc_hd__xnor2_1_40/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_349 vssd1 vccd1 sky130_fd_sc_hd__inv_2_20/Y sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__o21ai_1_349/B1 sky130_fd_sc_hd__xor2_1_165/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nand2_1_709 sky130_fd_sc_hd__nand2_1_709/Y la_data_out[68] sky130_fd_sc_hd__mux2_4_4/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_18 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_18/A1 sky130_fd_sc_hd__buf_2_144/X
+ sky130_fd_sc_hd__mux2_8_0/S sky130_fd_sc_hd__mux2_2_18/X vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_29 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_29/A1 sky130_fd_sc_hd__buf_2_71/X
+ sky130_fd_sc_hd__mux2_8_1/S sky130_fd_sc_hd__fa_2_416/B vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__conb_1_104 sky130_fd_sc_hd__conb_1_104/LO sky130_fd_sc_hd__conb_1_104/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_115 sky130_fd_sc_hd__conb_1_115/LO sky130_fd_sc_hd__conb_1_115/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_126 sky130_fd_sc_hd__conb_1_126/LO sky130_fd_sc_hd__conb_1_126/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_137 sky130_fd_sc_hd__conb_1_137/LO sky130_fd_sc_hd__clkinv_1_5/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_148 sky130_fd_sc_hd__conb_1_148/LO sky130_fd_sc_hd__conb_1_148/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__xor2_1_110 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__fa_2_83/CIN
+ sky130_fd_sc_hd__xor2_1_110/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_121 sky130_fd_sc_hd__xor2_1_9/B sky130_fd_sc_hd__fa_2_91/CIN
+ sky130_fd_sc_hd__xor2_1_121/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_132 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__fa_2_93/A
+ sky130_fd_sc_hd__xor2_1_132/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_143 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__fa_2_106/A
+ sky130_fd_sc_hd__xor2_1_143/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_154 sky130_fd_sc_hd__xor2_1_154/B sky130_fd_sc_hd__xor2_1_154/X
+ sky130_fd_sc_hd__xor2_1_154/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_505 sky130_fd_sc_hd__ha_2_42/A sky130_fd_sc_hd__dfxtp_1_509/CLK
+ sky130_fd_sc_hd__and2_0_398/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_165 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__xor2_1_165/X
+ sky130_fd_sc_hd__xor2_1_165/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_516 sky130_fd_sc_hd__ha_2_54/A sky130_fd_sc_hd__dfxtp_1_520/CLK
+ sky130_fd_sc_hd__and2_0_343/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_176 sky130_fd_sc_hd__xor2_1_176/B sky130_fd_sc_hd__xor2_1_176/X
+ sky130_fd_sc_hd__xor2_1_176/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_527 wbs_dat_o[6] sky130_fd_sc_hd__dfxtp_1_532/CLK sky130_fd_sc_hd__nor2b_1_151/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_187 sky130_fd_sc_hd__xor2_1_187/B sky130_fd_sc_hd__xor2_1_187/X
+ sky130_fd_sc_hd__xor2_1_187/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_538 wbs_dat_o[17] sky130_fd_sc_hd__dfxtp_1_538/CLK sky130_fd_sc_hd__nor2b_1_140/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_198 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__or2_0_16/A
+ sky130_fd_sc_hd__xor2_1_198/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_549 wbs_dat_o[28] sky130_fd_sc_hd__dfxtp_1_552/CLK sky130_fd_sc_hd__nor2b_1_129/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_103 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_48/A1 sky130_fd_sc_hd__clkbuf_1_103/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_114 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_114/X sky130_fd_sc_hd__clkinv_1_977/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_125 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_125/X sky130_fd_sc_hd__inv_4_2/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_136 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_136/X sky130_fd_sc_hd__clkinv_1_904/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_207 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__buf_2_32/X sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__o21ai_1_380/B1 sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_147 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_36/A1 sky130_fd_sc_hd__clkbuf_1_147/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_218 vccd1 vssd1 sky130_fd_sc_hd__and3_4_14/X sky130_fd_sc_hd__buf_2_31/X
+ sky130_fd_sc_hd__buf_2_19/X sky130_fd_sc_hd__nor2_1_127/Y sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__o21ai_1_407/B1 sky130_fd_sc_hd__nor2b_1_10/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_158 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_25/A1 sky130_fd_sc_hd__clkbuf_1_158/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_5 sky130_fd_sc_hd__dfxtp_1_5/Q sky130_fd_sc_hd__dfxtp_1_9/CLK
+ sky130_fd_sc_hd__dfxtp_1_5/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_850 vssd1 vccd1 sky130_fd_sc_hd__nand2_1_640/Y sky130_fd_sc_hd__a21oi_1_136/Y
+ sky130_fd_sc_hd__a21oi_1_134/Y sky130_fd_sc_hd__xnor2_1_179/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_229 vccd1 vssd1 sky130_fd_sc_hd__and3_4_17/X sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__nor2_1_73/B sky130_fd_sc_hd__nor2_2_20/Y sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__o21ai_1_420/B1 sky130_fd_sc_hd__nor2b_2_4/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_169 vssd1 vccd1 sky130_fd_sc_hd__a22o_1_35/B2 sky130_fd_sc_hd__clkbuf_1_169/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o21ai_1_861 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_861/A2 sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__nand2_1_501/Y sky130_fd_sc_hd__xor2_1_636/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_872 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_650/A sky130_fd_sc_hd__nor2_1_231/Y
+ sky130_fd_sc_hd__nand2_1_705/Y sky130_fd_sc_hd__xnor2_1_198/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_883 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_664/A sky130_fd_sc_hd__nor2_1_252/Y
+ sky130_fd_sc_hd__nand2_1_781/Y sky130_fd_sc_hd__xnor2_1_216/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_894 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_677/A sky130_fd_sc_hd__nor2_1_255/Y
+ sky130_fd_sc_hd__nand2_1_797/Y sky130_fd_sc_hd__xnor2_1_291/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__inv_4_15 sky130_fd_sc_hd__inv_4_15/Y wbs_dat_i[19] vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__and2_0_101 vccd1 vssd1 sky130_fd_sc_hd__and2_0_101/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__or2_0_9/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_112 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_97/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_112/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_20 la_data_out[107] sky130_fd_sc_hd__conb_1_122/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_123 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_99/D sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_123/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_31 la_data_out[96] sky130_fd_sc_hd__conb_1_111/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_8_3 sky130_fd_sc_hd__nand2_8_3/A sky130_fd_sc_hd__nand2_8_3/B
+ sky130_fd_sc_hd__nor2_1_87/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_8
Xsky130_fd_sc_hd__and2_0_134 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_69/D sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_134/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_42 la_data_out[21] sky130_fd_sc_hd__conb_1_100/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_145 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_39/D sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_145/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_53 la_data_out[10] sky130_fd_sc_hd__conb_1_89/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_156 vccd1 vssd1 sky130_fd_sc_hd__and2_0_156/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_156/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_64 io_out[37] sky130_fd_sc_hd__conb_1_78/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_167 vccd1 vssd1 sky130_fd_sc_hd__and2_0_167/X sky130_fd_sc_hd__o21ai_2_0/B1
+ sky130_fd_sc_hd__and2_0_167/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_75 io_out[26] sky130_fd_sc_hd__conb_1_67/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_178 vccd1 vssd1 sky130_fd_sc_hd__and2_0_178/X sky130_fd_sc_hd__o21ai_2_0/B1
+ sky130_fd_sc_hd__o21ai_1_99/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_86 io_out[15] sky130_fd_sc_hd__conb_1_56/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_189 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_80/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_91/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_97 io_out[4] sky130_fd_sc_hd__conb_1_45/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_0 sky130_fd_sc_hd__nand2_1_7/B sky130_fd_sc_hd__or2_0_75/B
+ sky130_fd_sc_hd__buf_4_5/A sky130_fd_sc_hd__or2_0_75/A sky130_fd_sc_hd__nand2_1_8/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__o21ai_1_102 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_105/A2 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_118/Y sky130_fd_sc_hd__and2_0_174/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_113 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_113/A2 sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__a22oi_1_167/Y sky130_fd_sc_hd__and2_0_162/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_124 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_125/A2 sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__a22oi_1_172/Y sky130_fd_sc_hd__and2_0_147/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_135 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_137/A2 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_135/Y sky130_fd_sc_hd__and2_0_134/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_146 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_149/A2 sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__a22oi_1_184/Y sky130_fd_sc_hd__and2_0_119/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_157 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_157/A2 sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__a22oi_1_189/Y sky130_fd_sc_hd__and2_0_107/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_168 vssd1 vccd1 sky130_fd_sc_hd__buf_2_5/X sky130_fd_sc_hd__nand2b_1_4/Y
+ sky130_fd_sc_hd__a222oi_1_50/Y sky130_fd_sc_hd__xor2_1_2/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_179 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_49/Y sky130_fd_sc_hd__nor2_1_46/A
+ sky130_fd_sc_hd__nor2_1_45/Y sky130_fd_sc_hd__o21ai_1_179/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nand2_1_506 sky130_fd_sc_hd__nand2_2_13/B sky130_fd_sc_hd__or2_0_72/A
+ sky130_fd_sc_hd__or2_0_72/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_517 sky130_fd_sc_hd__xor2_1_447/B sky130_fd_sc_hd__nand2_1_517/B
+ sky130_fd_sc_hd__nand2_1_517/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_528 sky130_fd_sc_hd__o21ai_2_12/B1 sky130_fd_sc_hd__nor2_2_21/A
+ sky130_fd_sc_hd__nor2_2_21/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_539 sky130_fd_sc_hd__o21ai_2_13/B1 sky130_fd_sc_hd__nor2_2_24/A
+ sky130_fd_sc_hd__nor2_2_24/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_8 sky130_fd_sc_hd__and3_1_1/C sky130_fd_sc_hd__nor2b_1_8/Y
+ sky130_fd_sc_hd__and3_1_1/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1108 sky130_fd_sc_hd__clkinv_4_51/A sky130_fd_sc_hd__a22o_1_28/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1119 sky130_fd_sc_hd__clkinv_4_62/A sky130_fd_sc_hd__a22o_1_39/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_80 sky130_fd_sc_hd__nand2_1_80/Y sky130_fd_sc_hd__nand2_1_80/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_91 sky130_fd_sc_hd__nand2_1_91/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__xnor2_1_73/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_302 sky130_fd_sc_hd__dfxtp_1_302/Q sky130_fd_sc_hd__clkinv_8_6/Y
+ sky130_fd_sc_hd__and2_0_278/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_313 sky130_fd_sc_hd__or2_0_91/A sky130_fd_sc_hd__dfxtp_1_319/CLK
+ sky130_fd_sc_hd__and2_0_290/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_324 sky130_fd_sc_hd__nor2_4_19/A sky130_fd_sc_hd__dfxtp_2_7/CLK
+ sky130_fd_sc_hd__nand2_1_789/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_335 sky130_fd_sc_hd__dfxtp_1_335/Q sky130_fd_sc_hd__dfxtp_1_339/CLK
+ sky130_fd_sc_hd__and2_0_330/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_346 sky130_fd_sc_hd__dfxtp_1_346/Q sky130_fd_sc_hd__dfxtp_1_354/CLK
+ sky130_fd_sc_hd__and2_0_311/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_357 sky130_fd_sc_hd__nor2_4_19/B sky130_fd_sc_hd__dfxtp_2_7/CLK
+ sky130_fd_sc_hd__ha_2_9/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_368 sky130_fd_sc_hd__dfxtp_1_368/Q sky130_fd_sc_hd__dfxtp_1_371/CLK
+ sky130_fd_sc_hd__nor2b_1_115/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_379 sky130_fd_sc_hd__dfxtp_1_379/Q sky130_fd_sc_hd__dfxtp_1_380/CLK
+ sky130_fd_sc_hd__nor2b_1_104/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_680 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_10/X sky130_fd_sc_hd__nand2_1_524/Y
+ sky130_fd_sc_hd__a21oi_1_111/Y sky130_fd_sc_hd__xnor2_1_137/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_691 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_691/A2 sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_691/B1 sky130_fd_sc_hd__xor2_1_471/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_207 sky130_fd_sc_hd__fa_2_194/B sky130_fd_sc_hd__fa_2_202/B
+ sky130_fd_sc_hd__fa_2_207/A sky130_fd_sc_hd__fa_2_207/B sky130_fd_sc_hd__xor2_1_299/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_218 sky130_fd_sc_hd__fa_2_212/A sky130_fd_sc_hd__fa_2_219/B
+ sky130_fd_sc_hd__fa_2_218/A sky130_fd_sc_hd__fa_2_218/B sky130_fd_sc_hd__xor2_1_314/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_229 sky130_fd_sc_hd__fa_2_226/CIN sky130_fd_sc_hd__fa_2_234/A
+ sky130_fd_sc_hd__fa_2_229/A sky130_fd_sc_hd__fa_2_229/B sky130_fd_sc_hd__xor2_1_333/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_10 sky130_fd_sc_hd__fa_2_1/B sky130_fd_sc_hd__fa_2_16/CIN sky130_fd_sc_hd__fa_2_10/A
+ sky130_fd_sc_hd__fa_2_10/B sky130_fd_sc_hd__fa_2_9/SUM vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_21 sky130_fd_sc_hd__fa_2_16/A sky130_fd_sc_hd__fa_2_26/A sky130_fd_sc_hd__fa_2_21/A
+ sky130_fd_sc_hd__fa_2_21/B sky130_fd_sc_hd__xor2_1_35/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_32 sky130_fd_sc_hd__fa_2_25/A sky130_fd_sc_hd__fa_2_33/B sky130_fd_sc_hd__fa_2_32/A
+ sky130_fd_sc_hd__fa_2_32/B sky130_fd_sc_hd__fa_2_32/CIN vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_43 sky130_fd_sc_hd__nor2_1_52/A sky130_fd_sc_hd__or2_0_2/B
+ sky130_fd_sc_hd__fa_2_43/A sky130_fd_sc_hd__fa_2_43/B sky130_fd_sc_hd__fa_2_43/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_54 sky130_fd_sc_hd__fa_2_47/A sky130_fd_sc_hd__fa_2_55/B sky130_fd_sc_hd__fa_2_54/A
+ sky130_fd_sc_hd__fa_2_54/B sky130_fd_sc_hd__fa_2_54/CIN vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_65 sky130_fd_sc_hd__fa_2_52/B sky130_fd_sc_hd__fa_2_60/B sky130_fd_sc_hd__fa_2_65/A
+ sky130_fd_sc_hd__fa_2_65/B sky130_fd_sc_hd__xor2_1_86/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_76 sky130_fd_sc_hd__fa_2_70/A sky130_fd_sc_hd__fa_2_77/B sky130_fd_sc_hd__fa_2_76/A
+ sky130_fd_sc_hd__fa_2_76/B sky130_fd_sc_hd__fa_2_76/CIN vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_87 sky130_fd_sc_hd__fa_2_84/CIN sky130_fd_sc_hd__fa_2_92/A
+ sky130_fd_sc_hd__fa_2_87/A sky130_fd_sc_hd__fa_2_87/B sky130_fd_sc_hd__fa_2_87/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_98 sky130_fd_sc_hd__nor2_1_69/A sky130_fd_sc_hd__or2_0_8/B
+ sky130_fd_sc_hd__fa_2_98/A sky130_fd_sc_hd__fa_2_98/B sky130_fd_sc_hd__fa_2_98/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_202 vccd1 vssd1 la_data_out[86] sky130_fd_sc_hd__nand2_2_7/Y
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_213 vccd1 vssd1 la_data_out[70] sky130_fd_sc_hd__buf_4_41/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__a21oi_1_15 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_44/Y
+ sky130_fd_sc_hd__a21oi_1_15/Y sky130_fd_sc_hd__dfxtp_1_82/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_560 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_410/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_442/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_757/A sky130_fd_sc_hd__dfxtp_1_378/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a21oi_1_26 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_55/Y
+ sky130_fd_sc_hd__a21oi_1_26/Y sky130_fd_sc_hd__dfxtp_1_71/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_571 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_399/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_431/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_768/A sky130_fd_sc_hd__dfxtp_1_367/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a21oi_1_37 sky130_fd_sc_hd__o21ai_1_221/Y sky130_fd_sc_hd__o21ai_1_179/Y
+ sky130_fd_sc_hd__o21a_1_0/B1 sky130_fd_sc_hd__nor2_1_46/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_582 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_414/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_446/Q sky130_fd_sc_hd__nor2_4_19/B
+ sky130_fd_sc_hd__clkinv_1_779/A sky130_fd_sc_hd__dfxtp_1_382/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a21oi_1_48 sky130_fd_sc_hd__nand2_1_229/Y sky130_fd_sc_hd__nor2_1_66/A
+ sky130_fd_sc_hd__a21oi_1_48/Y sky130_fd_sc_hd__or2_0_18/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_593 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_397/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_429/Q sky130_fd_sc_hd__clkbuf_1_32/X
+ sky130_fd_sc_hd__clkinv_1_790/A sky130_fd_sc_hd__dfxtp_1_365/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a21oi_1_59 sky130_fd_sc_hd__nor2_1_93/Y sky130_fd_sc_hd__o21ai_1_366/Y
+ sky130_fd_sc_hd__xor2_1_176/A sky130_fd_sc_hd__o21ai_1_372/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__decap_12_11 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_22 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_33 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_44 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_55 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_66 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_77 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_88 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_99 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_11 vccd1 vssd1 sky130_fd_sc_hd__buf_6_11/X sky130_fd_sc_hd__buf_6_11/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_22 vccd1 vssd1 sky130_fd_sc_hd__buf_6_22/X sky130_fd_sc_hd__buf_6_22/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_33 vccd1 vssd1 sky130_fd_sc_hd__buf_6_33/X sky130_fd_sc_hd__buf_8_92/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_44 vccd1 vssd1 sky130_fd_sc_hd__buf_6_44/X sky130_fd_sc_hd__buf_8_5/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_55 vccd1 vssd1 sky130_fd_sc_hd__buf_6_55/X sky130_fd_sc_hd__buf_6_55/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_66 vccd1 vssd1 sky130_fd_sc_hd__buf_6_66/X sky130_fd_sc_hd__buf_8_90/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_77 vccd1 vssd1 sky130_fd_sc_hd__buf_6_77/X sky130_fd_sc_hd__buf_6_77/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_88 vccd1 vssd1 sky130_fd_sc_hd__buf_6_88/X sky130_fd_sc_hd__buf_6_88/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_13 la_data_out[62] vssd1 vccd1 vccd1 vssd1 sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_24 sky130_fd_sc_hd__clkinv_4_61/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_35 sky130_fd_sc_hd__clkinv_4_51/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_46 sky130_fd_sc_hd__buf_2_189/A vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_57 sky130_fd_sc_hd__buf_2_192/A vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_68 la_data_out[62] vssd1 vccd1 vccd1 vssd1 sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__decap_12_408 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_419 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_303 sky130_fd_sc_hd__nand2_1_303/Y sky130_fd_sc_hd__buf_4_6/X
+ sky130_fd_sc_hd__buf_4_1/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_902 sky130_fd_sc_hd__clkinv_1_902/Y sky130_fd_sc_hd__clkinv_4_90/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_314 sky130_fd_sc_hd__nand2_1_314/Y sky130_fd_sc_hd__o21ai_1_33/Y
+ sky130_fd_sc_hd__xor2_1_208/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_913 sky130_fd_sc_hd__clkinv_1_913/Y sky130_fd_sc_hd__inv_2_107/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_325 sky130_fd_sc_hd__nand2_1_325/Y sky130_fd_sc_hd__nor2_1_127/Y
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_924 sky130_fd_sc_hd__inv_2_116/A sky130_fd_sc_hd__buf_8_99/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_336 sky130_fd_sc_hd__xnor2_1_69/A sky130_fd_sc_hd__nand2_1_337/Y
+ sky130_fd_sc_hd__or2_0_31/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_935 sky130_fd_sc_hd__inv_2_125/A sky130_fd_sc_hd__buf_8_91/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_347 sky130_fd_sc_hd__nor2_1_112/A sky130_fd_sc_hd__or2_0_39/X
+ sky130_fd_sc_hd__nand2_1_359/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_946 sky130_fd_sc_hd__inv_2_145/A sky130_fd_sc_hd__dfxtp_1_17/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_358 sky130_fd_sc_hd__nor2_1_115/A sky130_fd_sc_hd__nand2_1_370/A
+ sky130_fd_sc_hd__or2_0_42/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_957 sky130_fd_sc_hd__clkinv_1_959/A sky130_fd_sc_hd__buf_2_143/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_369 sky130_fd_sc_hd__nor2_1_118/B sky130_fd_sc_hd__or2_0_40/X
+ sky130_fd_sc_hd__or2_0_41/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_968 sky130_fd_sc_hd__clkinv_1_968/Y sky130_fd_sc_hd__clkinv_4_22/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_979 sky130_fd_sc_hd__clkinv_1_979/Y sky130_fd_sc_hd__clkinv_4_26/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1407 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_110 sky130_fd_sc_hd__dfxtp_1_110/Q sky130_fd_sc_hd__dfxtp_1_99/CLK
+ sky130_fd_sc_hd__and2_0_179/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1418 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_121 sky130_fd_sc_hd__dfxtp_1_121/Q sky130_fd_sc_hd__dfxtp_1_122/CLK
+ sky130_fd_sc_hd__and2_0_233/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1429 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_132 sky130_fd_sc_hd__dfxtp_1_132/Q sky130_fd_sc_hd__dfxtp_1_138/CLK
+ sky130_fd_sc_hd__and2_0_131/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_143 sky130_fd_sc_hd__dfxtp_1_143/Q sky130_fd_sc_hd__dfxtp_1_146/CLK
+ sky130_fd_sc_hd__and2_0_184/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_154 sky130_fd_sc_hd__dfxtp_1_154/Q sky130_fd_sc_hd__dfxtp_1_154/CLK
+ sky130_fd_sc_hd__and2_0_241/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_165 sky130_fd_sc_hd__dfxtp_1_165/Q sky130_fd_sc_hd__dfxtp_1_170/CLK
+ sky130_fd_sc_hd__and2_0_133/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_176 sky130_fd_sc_hd__dfxtp_1_176/Q sky130_fd_sc_hd__dfxtp_1_176/CLK
+ sky130_fd_sc_hd__and2_0_187/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_187 sky130_fd_sc_hd__dfxtp_1_187/Q sky130_fd_sc_hd__dfxtp_1_190/CLK
+ sky130_fd_sc_hd__and2_0_242/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_198 sky130_fd_sc_hd__xor2_1_609/A sky130_fd_sc_hd__dfxtp_2_1/CLK
+ sky130_fd_sc_hd__and2_0_43/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_920 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_931 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_942 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_953 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_964 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_975 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_986 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_997 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o211ai_1_18 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_45/B1
+ sky130_fd_sc_hd__o211ai_1_18/Y sky130_fd_sc_hd__a22oi_1_68/Y sky130_fd_sc_hd__a22oi_1_69/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_29 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_32/B1
+ sky130_fd_sc_hd__o211ai_1_29/Y sky130_fd_sc_hd__a22oi_1_90/Y sky130_fd_sc_hd__a22oi_1_91/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o21ai_1_70 vssd1 vccd1 sky130_fd_sc_hd__inv_2_57/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__o21ai_1_70/B1 sky130_fd_sc_hd__o21ai_1_70/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_81 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_81/A2 sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__o21ai_1_81/B1 sky130_fd_sc_hd__o21ai_1_81/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_92 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_93/A2 sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_92/B1 sky130_fd_sc_hd__o21ai_1_92/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_390 vccd1 vssd1 sky130_fd_sc_hd__and3_4_23/X sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__buf_4_7/X sky130_fd_sc_hd__nor2_1_178/Y sky130_fd_sc_hd__buf_4_0/X
+ sky130_fd_sc_hd__o21ai_1_653/B1 sky130_fd_sc_hd__nor2b_1_15/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkinv_1_209 sky130_fd_sc_hd__nor2_1_16/A sky130_fd_sc_hd__dfxtp_1_139/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_2_9 sky130_fd_sc_hd__o21ai_2_9/B1 sky130_fd_sc_hd__o21ai_2_9/Y
+ sky130_fd_sc_hd__xor2_1_346/A sky130_fd_sc_hd__nor2_2_14/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__o21ai_2
Xsky130_fd_sc_hd__a21oi_1_106 sky130_fd_sc_hd__clkinv_1_615/Y sky130_fd_sc_hd__o21ai_1_786/Y
+ sky130_fd_sc_hd__xnor2_1_126/A sky130_fd_sc_hd__nor2_1_188/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_117 sky130_fd_sc_hd__o21ai_1_753/Y sky130_fd_sc_hd__nor2_1_179/A
+ sky130_fd_sc_hd__a21oi_1_117/Y sky130_fd_sc_hd__or2_0_65/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_128 sky130_fd_sc_hd__nand2_1_614/Y sky130_fd_sc_hd__clkinv_1_585/Y
+ sky130_fd_sc_hd__a21oi_1_128/Y sky130_fd_sc_hd__nand2_1_615/A vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_139 sky130_fd_sc_hd__xnor2_1_189/B sky130_fd_sc_hd__clkinv_1_627/Y
+ sky130_fd_sc_hd__xor2_1_640/A sky130_fd_sc_hd__or2_0_74/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_510 sky130_fd_sc_hd__buf_12_510/A sky130_fd_sc_hd__buf_12_551/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_521 sky130_fd_sc_hd__buf_12_521/A sky130_fd_sc_hd__buf_12_521/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_532 sky130_fd_sc_hd__buf_12_532/A sky130_fd_sc_hd__buf_12_532/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_543 sky130_fd_sc_hd__buf_12_543/A sky130_fd_sc_hd__buf_12_543/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_554 sky130_fd_sc_hd__buf_12_554/A sky130_fd_sc_hd__buf_12_554/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_565 sky130_fd_sc_hd__buf_12_565/A sky130_fd_sc_hd__buf_12_565/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_8_2 sky130_fd_sc_hd__buf_12_65/A sky130_fd_sc_hd__buf_12_9/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_8
Xsky130_fd_sc_hd__buf_12_576 sky130_fd_sc_hd__buf_12_576/A sky130_fd_sc_hd__buf_12_576/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_205 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_587 sky130_fd_sc_hd__buf_12_587/A sky130_fd_sc_hd__buf_12_587/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_216 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_598 sky130_fd_sc_hd__buf_12_598/A sky130_fd_sc_hd__buf_12_598/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__nand2_1_100 sky130_fd_sc_hd__o21ai_1_66/B1 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__xor2_1_296/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_227 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_111 sky130_fd_sc_hd__o21ai_1_87/B1 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__xnor2_1_95/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_238 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_710 sky130_fd_sc_hd__nor2b_1_89/A sky130_fd_sc_hd__xor2_1_674/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_122 sky130_fd_sc_hd__nand2_1_122/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_123/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_249 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_721 sky130_fd_sc_hd__nor2b_1_100/A sky130_fd_sc_hd__xor2_1_679/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_133 sky130_fd_sc_hd__nand2_1_133/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_133/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_732 sky130_fd_sc_hd__nor2b_1_111/A sky130_fd_sc_hd__xnor2_1_299/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_144 sky130_fd_sc_hd__nand2_1_144/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__xor2_1_421/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_743 sky130_fd_sc_hd__fa_2_465/A sky130_fd_sc_hd__clkinv_1_743/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_306 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_306/B sky130_fd_sc_hd__nand4_1_2/B
+ la_data_out[39] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_155 sky130_fd_sc_hd__nand2_1_155/Y sky130_fd_sc_hd__nor2_1_68/Y
+ sky130_fd_sc_hd__clkbuf_1_3/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_754 sky130_fd_sc_hd__fa_2_477/A sky130_fd_sc_hd__clkinv_1_754/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_166 sky130_fd_sc_hd__nand2_1_166/Y sky130_fd_sc_hd__or2_0_9/A
+ sky130_fd_sc_hd__or2_0_4/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_765 sky130_fd_sc_hd__fa_2_488/A sky130_fd_sc_hd__clkinv_1_765/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_177 sky130_fd_sc_hd__xnor2_1_9/A sky130_fd_sc_hd__nand2_1_178/Y
+ sky130_fd_sc_hd__or2_0_10/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_776 sky130_fd_sc_hd__and2_0_331/A sky130_fd_sc_hd__clkinv_1_776/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_188 sky130_fd_sc_hd__xnor2_1_13/A sky130_fd_sc_hd__nand2_1_189/Y
+ sky130_fd_sc_hd__nand2_1_188/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_787 sky130_fd_sc_hd__and2_0_320/A sky130_fd_sc_hd__clkinv_1_787/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_199 sky130_fd_sc_hd__xnor2_1_17/A sky130_fd_sc_hd__nand2_1_200/Y
+ sky130_fd_sc_hd__nand2_1_199/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_798 sky130_fd_sc_hd__and2_0_309/A sky130_fd_sc_hd__clkinv_1_798/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1204 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_4 sky130_fd_sc_hd__fa_2_97/A sky130_fd_sc_hd__xor3_1_3/A
+ sky130_fd_sc_hd__xor2_1_4/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1215 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1226 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1237 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1248 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1259 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_8_2 sky130_fd_sc_hd__clkinv_8_3/A sky130_fd_sc_hd__clkinv_8_2/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__xor2_1_19 sky130_fd_sc_hd__fa_2_28/A sky130_fd_sc_hd__fa_2_6/B sky130_fd_sc_hd__xor2_1_19/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_750 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_761 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_772 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_783 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_794 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_506 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__xor2_1_506/X
+ sky130_fd_sc_hd__xor2_1_506/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_517 sky130_fd_sc_hd__fa_2_379/A sky130_fd_sc_hd__fa_2_343/A
+ sky130_fd_sc_hd__xor2_1_517/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_528 sky130_fd_sc_hd__fa_2_379/A sky130_fd_sc_hd__fa_2_360/B
+ sky130_fd_sc_hd__xor2_1_528/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_539 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__xor2_1_539/X
+ sky130_fd_sc_hd__xor2_1_539/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1760 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1771 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_70 sky130_fd_sc_hd__inv_2_70/A sky130_fd_sc_hd__inv_2_70/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1782 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_81 sky130_fd_sc_hd__inv_2_81/A sky130_fd_sc_hd__inv_2_81/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1793 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_92 sky130_fd_sc_hd__inv_2_92/A sky130_fd_sc_hd__inv_2_92/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__ha_2_13 vssd1 vccd1 sky130_fd_sc_hd__ha_2_13/A sky130_fd_sc_hd__ha_2_13/COUT
+ sky130_fd_sc_hd__fa_2_439/A sky130_fd_sc_hd__ha_2_13/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_24 vssd1 vccd1 sky130_fd_sc_hd__ha_2_24/A sky130_fd_sc_hd__ha_2_23/B
+ sky130_fd_sc_hd__ha_2_24/SUM sky130_fd_sc_hd__ha_2_24/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_35 vssd1 vccd1 sky130_fd_sc_hd__ha_2_35/A sky130_fd_sc_hd__ha_2_34/B
+ sky130_fd_sc_hd__ha_2_35/SUM sky130_fd_sc_hd__ha_2_35/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_46 vssd1 vccd1 sky130_fd_sc_hd__ha_2_46/A sky130_fd_sc_hd__ha_2_45/B
+ sky130_fd_sc_hd__ha_2_46/SUM sky130_fd_sc_hd__ha_2_46/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__and2b_4_8 sky130_fd_sc_hd__nor2_4_13/A sky130_fd_sc_hd__and2b_4_8/X
+ sky130_fd_sc_hd__and3_4_11/C vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__and2b_4
Xsky130_fd_sc_hd__ha_2_57 vssd1 vccd1 sky130_fd_sc_hd__ha_2_57/A sky130_fd_sc_hd__ha_2_60/B
+ sky130_fd_sc_hd__ha_2_57/SUM sky130_fd_sc_hd__ha_2_57/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__sdlclkp_4_20 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_8_1/Y
+ sky130_fd_sc_hd__dfxtp_2_0/CLK sky130_fd_sc_hd__o21ai_2_2/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_390 sky130_fd_sc_hd__fa_2_387/B sky130_fd_sc_hd__fah_1_16/CI
+ sky130_fd_sc_hd__fa_2_390/A sky130_fd_sc_hd__fa_2_390/B sky130_fd_sc_hd__fa_2_390/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_31 sky130_fd_sc_hd__conb_1_144/LO sky130_fd_sc_hd__clkinv_4_99/Y
+ sky130_fd_sc_hd__dfxtp_1_319/CLK sky130_fd_sc_hd__nand2_1_713/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__clkbuf_1_9 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_9/X sky130_fd_sc_hd__clkbuf_1_9/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__sdlclkp_4_42 sky130_fd_sc_hd__conb_1_145/LO sky130_fd_sc_hd__clkinv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_427/CLK sky130_fd_sc_hd__o21ai_1_891/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_53 sky130_fd_sc_hd__conb_1_149/LO sky130_fd_sc_hd__clkinv_4_117/A
+ sky130_fd_sc_hd__dfxtp_1_544/CLK sky130_fd_sc_hd__or2_0_113/X vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_100 sky130_fd_sc_hd__nor2_2_6/Y sky130_fd_sc_hd__nor2_1_100/Y
+ sky130_fd_sc_hd__nor2_1_102/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_111 sky130_fd_sc_hd__nor2_1_111/B sky130_fd_sc_hd__nor2_1_111/Y
+ sky130_fd_sc_hd__nor2_1_111/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_122 sky130_fd_sc_hd__nor2_1_122/B sky130_fd_sc_hd__nor2_1_122/Y
+ sky130_fd_sc_hd__nor2_1_122/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_133 sky130_fd_sc_hd__nor2_1_137/Y sky130_fd_sc_hd__nor2_1_133/Y
+ sky130_fd_sc_hd__nor2_1_135/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_144 sky130_fd_sc_hd__nor2_1_85/B sky130_fd_sc_hd__nor2_1_144/Y
+ sky130_fd_sc_hd__nor2_1_87/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_20 sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__dfxtp_1_281/Q sky130_fd_sc_hd__o211ai_1_5/Y sky130_fd_sc_hd__nand2_1_15/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_155 sky130_fd_sc_hd__nor2_1_155/B sky130_fd_sc_hd__nor2_1_155/Y
+ sky130_fd_sc_hd__nor2_1_155/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_31 sky130_fd_sc_hd__nor2_4_0/Y sky130_fd_sc_hd__nor2_2_0/Y
+ sky130_fd_sc_hd__dfxtp_1_325/Q sky130_fd_sc_hd__or2_0_85/A sky130_fd_sc_hd__nand2_2_7/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_9 la_data_out[118] sky130_fd_sc_hd__clkinv_1_9/A vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_166 sky130_fd_sc_hd__nor2_1_170/B sky130_fd_sc_hd__nor2_1_166/Y
+ sky130_fd_sc_hd__nor2_1_166/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_42 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__clkbuf_1_25/X
+ sky130_fd_sc_hd__nand2_1_78/B sky130_fd_sc_hd__dfxtp_1_132/Q sky130_fd_sc_hd__a22oi_1_42/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_177 sky130_fd_sc_hd__or2_0_61/A sky130_fd_sc_hd__nor2_1_177/Y
+ sky130_fd_sc_hd__or2_0_60/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_53 sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__dfxtp_1_105/Q sky130_fd_sc_hd__dfxtp_1_73/Q sky130_fd_sc_hd__a22oi_1_53/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_64 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__nor2_4_3/Y
+ sky130_fd_sc_hd__nand2_1_67/B sky130_fd_sc_hd__dfxtp_1_143/Q sky130_fd_sc_hd__a22oi_1_64/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_188 sky130_fd_sc_hd__nor2_1_188/B sky130_fd_sc_hd__nor2_1_188/Y
+ sky130_fd_sc_hd__nor2_1_188/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_199 sky130_fd_sc_hd__buf_2_21/X sky130_fd_sc_hd__nor2_1_199/Y
+ sky130_fd_sc_hd__nor2_1_87/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_75 sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__dfxtp_1_116/Q sky130_fd_sc_hd__dfxtp_1_84/Q sky130_fd_sc_hd__a22oi_1_75/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_86 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__nor2_4_3/Y
+ sky130_fd_sc_hd__nand2_1_54/B sky130_fd_sc_hd__dfxtp_1_154/Q sky130_fd_sc_hd__a22oi_1_86/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_97 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_187/Q sky130_fd_sc_hd__dfxtp_1_155/Q sky130_fd_sc_hd__o21ai_1_3/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_340 sky130_fd_sc_hd__buf_12_65/X sky130_fd_sc_hd__buf_12_506/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_351 sky130_fd_sc_hd__buf_12_351/A sky130_fd_sc_hd__buf_12_591/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_210 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__and2b_4_8/X sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__a22oi_1_210/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_362 sky130_fd_sc_hd__buf_12_362/A sky130_fd_sc_hd__buf_12_553/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_221 sky130_fd_sc_hd__buf_2_28/A sky130_fd_sc_hd__buf_2_25/A
+ sky130_fd_sc_hd__and2b_4_12/X sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__a22oi_1_221/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_373 sky130_fd_sc_hd__buf_12_373/A sky130_fd_sc_hd__buf_12_557/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_384 sky130_fd_sc_hd__buf_12_384/A sky130_fd_sc_hd__buf_12_657/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_395 sky130_fd_sc_hd__buf_12_395/A sky130_fd_sc_hd__buf_12_576/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_540 sky130_fd_sc_hd__nand2_1_538/A sky130_fd_sc_hd__nor2_2_24/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_103 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_103/B sky130_fd_sc_hd__inv_2_38/A
+ sky130_fd_sc_hd__xnor2_1_103/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_551 sky130_fd_sc_hd__nand2_1_549/A sky130_fd_sc_hd__nor2_2_23/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_114 vssd1 vccd1 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__nor2_4_12/A
+ sky130_fd_sc_hd__xnor2_1_114/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_562 sky130_fd_sc_hd__a21oi_2_17/B1 sky130_fd_sc_hd__nand2_1_566/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_125 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_423/X sky130_fd_sc_hd__xnor2_1_125/Y
+ sky130_fd_sc_hd__xnor2_1_125/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_573 sky130_fd_sc_hd__nand2_1_581/A sky130_fd_sc_hd__nor2_1_187/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_136 vssd1 vccd1 sky130_fd_sc_hd__o21ai_2_12/Y sky130_fd_sc_hd__inv_2_63/A
+ sky130_fd_sc_hd__xnor2_1_136/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_584 sky130_fd_sc_hd__nand2_1_607/A sky130_fd_sc_hd__nor2_2_30/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_147 vssd1 vccd1 sky130_fd_sc_hd__fa_2_357/A sky130_fd_sc_hd__and3_4_23/C
+ sky130_fd_sc_hd__xnor2_1_147/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_595 sky130_fd_sc_hd__nand2_1_623/A sky130_fd_sc_hd__nor2_1_207/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_158 vssd1 vccd1 sky130_fd_sc_hd__o21ai_2_15/Y sky130_fd_sc_hd__xnor2_1_158/Y
+ sky130_fd_sc_hd__xnor2_1_158/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_4_20 sky130_fd_sc_hd__conb_1_147/HI sky130_fd_sc_hd__clkinv_4_20/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__xnor2_1_169 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_169/B sky130_fd_sc_hd__xnor2_1_169/Y
+ sky130_fd_sc_hd__xnor2_1_169/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_4_31 sky130_fd_sc_hd__nand2_2_2/Y sky130_fd_sc_hd__clkinv_4_31/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_42 sky130_fd_sc_hd__clkinv_8_32/Y sky130_fd_sc_hd__clkinv_8_33/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_53 sky130_fd_sc_hd__clkinv_4_53/A sky130_fd_sc_hd__clkinv_4_53/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_64 sky130_fd_sc_hd__clkinv_4_64/A sky130_fd_sc_hd__clkinv_4_64/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_75 sky130_fd_sc_hd__clkinv_4_75/A sky130_fd_sc_hd__clkinv_4_75/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_1001 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_4_86 wbs_dat_i[17] sky130_fd_sc_hd__clkinv_4_86/Y vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_1012 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_4_97 sky130_fd_sc_hd__clkinv_8_50/Y sky130_fd_sc_hd__clkinv_4_97/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_1023 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1034 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1045 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1056 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1067 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_16_5 sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_5/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__decap_12_1078 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_509 vssd1 vccd1 sky130_fd_sc_hd__nand2_2_12/Y sky130_fd_sc_hd__nand2b_1_13/Y
+ sky130_fd_sc_hd__a22oi_1_205/Y sky130_fd_sc_hd__xor2_1_308/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1089 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__and2b_4_12 sky130_fd_sc_hd__nor2_4_17/A sky130_fd_sc_hd__and2b_4_12/X
+ sky130_fd_sc_hd__and3_4_21/C vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__and2b_4
Xsky130_fd_sc_hd__decap_12_580 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_591 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_303 sky130_fd_sc_hd__fa_2_217/A sky130_fd_sc_hd__xor2_1_303/X
+ sky130_fd_sc_hd__xor2_1_303/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_314 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__xor2_1_314/X
+ sky130_fd_sc_hd__xor2_1_314/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_325 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__fa_2_225/A
+ sky130_fd_sc_hd__xor2_1_325/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_336 sky130_fd_sc_hd__fa_2_239/A sky130_fd_sc_hd__fa_2_232/B
+ sky130_fd_sc_hd__xor2_1_336/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_347 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__xor2_1_347/X
+ sky130_fd_sc_hd__xor2_1_347/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_358 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__fa_2_248/B
+ sky130_fd_sc_hd__xor2_1_358/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_369 sky130_fd_sc_hd__dfxtp_2_5/Q sky130_fd_sc_hd__fa_2_254/A
+ sky130_fd_sc_hd__xor2_1_369/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_307 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2_40/A sky130_fd_sc_hd__buf_8_122/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_318 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_318/X sky130_fd_sc_hd__clkinv_1_882/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_12_1590 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_329 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1_553/D sky130_fd_sc_hd__nor3_1_4/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_11 sky130_fd_sc_hd__buf_8_6/A sky130_fd_sc_hd__dfxtp_1_9/CLK
+ sky130_fd_sc_hd__dfxtp_1_11/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_22 sky130_fd_sc_hd__or4_1_1/C sky130_fd_sc_hd__dfxtp_1_29/CLK
+ sky130_fd_sc_hd__or4_1_3/C vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_33 sky130_fd_sc_hd__nand2_1_83/B sky130_fd_sc_hd__dfxtp_1_46/CLK
+ sky130_fd_sc_hd__dfxtp_1_33/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_44 sky130_fd_sc_hd__nand2_1_70/B sky130_fd_sc_hd__dfxtp_1_46/CLK
+ sky130_fd_sc_hd__dfxtp_1_44/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_55 sky130_fd_sc_hd__nand2_1_58/B sky130_fd_sc_hd__dfxtp_1_57/CLK
+ sky130_fd_sc_hd__dfxtp_1_55/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_66 sky130_fd_sc_hd__dfxtp_1_66/Q sky130_fd_sc_hd__dfxtp_1_78/CLK
+ sky130_fd_sc_hd__dfxtp_1_66/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_77 sky130_fd_sc_hd__dfxtp_1_77/Q sky130_fd_sc_hd__dfxtp_1_78/CLK
+ sky130_fd_sc_hd__dfxtp_1_77/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_88 sky130_fd_sc_hd__dfxtp_1_88/Q sky130_fd_sc_hd__dfxtp_1_89/CLK
+ sky130_fd_sc_hd__dfxtp_1_88/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_99 sky130_fd_sc_hd__dfxtp_1_99/Q sky130_fd_sc_hd__dfxtp_1_99/CLK
+ sky130_fd_sc_hd__dfxtp_1_99/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_305 vccd1 vssd1 sky130_fd_sc_hd__and2_0_305/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_305/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_316 vccd1 vssd1 sky130_fd_sc_hd__and2_0_316/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_316/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_327 vccd1 vssd1 sky130_fd_sc_hd__and2_0_327/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_327/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_338 vccd1 vssd1 sky130_fd_sc_hd__and2_0_395/A sky130_fd_sc_hd__ha_2_45/SUM
+ sky130_fd_sc_hd__and2_0_342/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_349 vccd1 vssd1 sky130_fd_sc_hd__and2_0_349/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__clkbuf_4_8/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__inv_2_105 sky130_fd_sc_hd__inv_2_105/A sky130_fd_sc_hd__inv_2_105/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_116 sky130_fd_sc_hd__inv_2_116/A sky130_fd_sc_hd__buf_8_72/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__or2_0_7 sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__or2_0_7/X sky130_fd_sc_hd__or2_0_7/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__inv_2_127 sky130_fd_sc_hd__buf_8_66/A sky130_fd_sc_hd__inv_2_129/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_138 sky130_fd_sc_hd__inv_2_138/A sky130_fd_sc_hd__buf_12_3/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_149 sky130_fd_sc_hd__buf_8_2/A sky130_fd_sc_hd__inv_2_150/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_sram_1kbyte_1rw1r_32x256_8_1 sky130_fd_sc_hd__clkinv_1_964/Y sky130_fd_sc_hd__clkinv_1_964/Y
+ sky130_fd_sc_hd__buf_12_670/X sky130_fd_sc_hd__buf_12_471/X sky130_fd_sc_hd__buf_12_568/X
+ sky130_fd_sc_hd__buf_12_453/X sky130_fd_sc_hd__buf_12_454/X sky130_fd_sc_hd__buf_12_645/X
+ sky130_fd_sc_hd__buf_12_613/X sky130_fd_sc_hd__clkbuf_1_111/X sky130_fd_sc_hd__buf_12_666/X
+ sky130_fd_sc_hd__buf_12_597/X sky130_fd_sc_hd__buf_12_586/X vccd1 sky130_fd_sc_hd__clkinv_8_38/Y
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[16] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[17]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[18] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[19]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[20] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[21]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[22] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[23]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[24] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[25]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[26] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[27]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[28] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[29]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[30] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[31]
+ sky130_fd_sc_hd__buf_12_528/X sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[1] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[2]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[3] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[4]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[5] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[6]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[7] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[8]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[9] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[10]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[11] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[12]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[13] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[14]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[15] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout1[0]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[10] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[11]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[12] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[13]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[14] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[15]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[16] sky130_fd_sc_hd__buf_12_535/X sky130_fd_sc_hd__buf_12_267/X
+ sky130_fd_sc_hd__buf_12_80/X sky130_fd_sc_hd__buf_12_52/X sky130_fd_sc_hd__buf_12_88/X
+ sky130_fd_sc_hd__clkinv_8_40/Y sky130_fd_sc_hd__buf_2_136/X sky130_fd_sc_hd__buf_2_136/X
+ sky130_fd_sc_hd__buf_2_136/X sky130_fd_sc_hd__buf_2_136/X sky130_fd_sc_hd__buf_2_136/X
+ sky130_fd_sc_hd__buf_2_136/X sky130_fd_sc_hd__buf_2_136/A sky130_fd_sc_hd__buf_2_136/A
+ sky130_fd_sc_hd__buf_2_136/A sky130_fd_sc_hd__buf_2_136/A sky130_fd_sc_hd__buf_2_136/A
+ sky130_fd_sc_hd__buf_2_136/A sky130_fd_sc_hd__buf_2_136/A sky130_fd_sc_hd__buf_12_1/X
+ sky130_fd_sc_hd__buf_12_1/X sky130_fd_sc_hd__buf_12_1/X sky130_fd_sc_hd__buf_12_1/X
+ sky130_fd_sc_hd__buf_12_1/X sky130_fd_sc_hd__buf_12_1/X sky130_fd_sc_hd__buf_12_1/X
+ sky130_fd_sc_hd__buf_12_1/X sky130_fd_sc_hd__buf_12_1/X sky130_fd_sc_hd__buf_12_1/X
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[0] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[1]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[2] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[3]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[4] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[5]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[6] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[7]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[8] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[9]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[25] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[26]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[27] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[28]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[29] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[30]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[31] sky130_fd_sc_hd__buf_12_1/X sky130_fd_sc_hd__buf_12_1/X
+ sky130_fd_sc_hd__buf_12_1/X sky130_fd_sc_hd__buf_12_1/X sky130_fd_sc_hd__buf_12_1/X
+ sky130_fd_sc_hd__buf_12_1/X sky130_fd_sc_hd__buf_12_1/X sky130_fd_sc_hd__buf_12_1/X
+ sky130_fd_sc_hd__buf_12_1/X sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[17] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[18]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[19] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[20]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[21] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[22]
+ sky130_fd_sc_hd__buf_12_668/X sky130_fd_sc_hd__buf_12_548/X sky130_fd_sc_hd__buf_12_496/X
+ sky130_fd_sc_hd__buf_12_539/X sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[23] sky130_sram_1kbyte_1rw1r_32x256_8_1/dout0[24]
+ sky130_sram_1kbyte_1rw1r_32x256_8_1/sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/gnd_uq26
+ vssd1 sky130_sram_1kbyte_1rw1r_32x256_8
Xsky130_fd_sc_hd__buf_12_170 sky130_fd_sc_hd__buf_12_33/X sky130_fd_sc_hd__buf_12_300/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_181 sky130_fd_sc_hd__buf_12_55/X sky130_fd_sc_hd__buf_12_320/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_192 sky130_fd_sc_hd__buf_4_30/X sky130_fd_sc_hd__buf_12_283/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_370 sky130_fd_sc_hd__a21oi_1_54/A1 sky130_fd_sc_hd__a21oi_1_57/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_381 sky130_fd_sc_hd__o21ai_1_356/B1 sky130_fd_sc_hd__nand2_1_272/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_392 sky130_fd_sc_hd__nand2_1_296/A sky130_fd_sc_hd__nor2_1_99/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_2_0 sky130_fd_sc_hd__a21oi_2_0/B1 sky130_fd_sc_hd__or2_0_1/X
+ sky130_fd_sc_hd__o21ai_2_5/Y sky130_fd_sc_hd__xor2_1_21/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_2
Xsky130_fd_sc_hd__a211o_1_6 vssd1 vccd1 sky130_fd_sc_hd__fa_2_277/B sky130_fd_sc_hd__dfxtp_1_69/Q
+ sky130_fd_sc_hd__nor2_1_10/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_6/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__o21ai_1_306 vssd1 vccd1 sky130_fd_sc_hd__buf_2_1/X sky130_fd_sc_hd__nand2b_1_1/Y
+ sky130_fd_sc_hd__o21ai_1_306/B1 sky130_fd_sc_hd__xor2_1_126/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_317 vssd1 vccd1 sky130_fd_sc_hd__inv_2_13/Y sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__o21ai_1_317/B1 sky130_fd_sc_hd__xor2_1_137/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_328 vssd1 vccd1 sky130_fd_sc_hd__buf_2_3/X sky130_fd_sc_hd__nand2b_1_1/Y
+ sky130_fd_sc_hd__o21ai_1_328/B1 sky130_fd_sc_hd__xor2_1_147/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_339 vssd1 vccd1 sky130_fd_sc_hd__buf_2_2/X sky130_fd_sc_hd__nand2b_1_1/Y
+ sky130_fd_sc_hd__o21ai_1_339/B1 sky130_fd_sc_hd__xor2_1_158/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__mux2_2_19 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_19/A1 sky130_fd_sc_hd__buf_2_86/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__fa_2_418/A vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__conb_1_105 sky130_fd_sc_hd__conb_1_105/LO sky130_fd_sc_hd__conb_1_105/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_116 sky130_fd_sc_hd__conb_1_116/LO sky130_fd_sc_hd__conb_1_116/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_127 sky130_fd_sc_hd__conb_1_127/LO sky130_fd_sc_hd__conb_1_127/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_138 sky130_fd_sc_hd__conb_1_138/LO sky130_fd_sc_hd__clkinv_1_4/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_149 sky130_fd_sc_hd__conb_1_149/LO sky130_fd_sc_hd__conb_1_149/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__xor2_1_100 sky130_fd_sc_hd__xor2_1_100/B sky130_fd_sc_hd__xor2_1_100/X
+ sky130_fd_sc_hd__a21oi_2_4/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_111 sky130_fd_sc_hd__fa_2_122/A sky130_fd_sc_hd__fa_2_83/B
+ sky130_fd_sc_hd__xor2_1_111/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_122 sky130_fd_sc_hd__fa_2_110/A sky130_fd_sc_hd__fa_2_91/B
+ sky130_fd_sc_hd__xor2_1_122/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_133 sky130_fd_sc_hd__xor2_1_133/B sky130_fd_sc_hd__xor2_1_133/X
+ sky130_fd_sc_hd__a21oi_2_6/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_144 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__xor2_1_144/X
+ sky130_fd_sc_hd__xor2_1_144/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_155 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__fa_2_114/B
+ sky130_fd_sc_hd__xor2_1_155/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_506 sky130_fd_sc_hd__or4_1_3/A sky130_fd_sc_hd__dfxtp_1_509/CLK
+ sky130_fd_sc_hd__and2_0_397/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_166 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__fa_2_121/B
+ sky130_fd_sc_hd__xor2_1_166/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_517 sky130_fd_sc_hd__ha_2_57/A sky130_fd_sc_hd__dfxtp_1_520/CLK
+ sky130_fd_sc_hd__and2_0_349/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_177 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__xor2_1_177/X
+ sky130_fd_sc_hd__xor2_1_177/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_528 wbs_dat_o[7] sky130_fd_sc_hd__dfxtp_1_532/CLK sky130_fd_sc_hd__nor2b_1_150/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_188 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__xor2_1_188/X
+ sky130_fd_sc_hd__xor2_1_188/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_539 wbs_dat_o[18] sky130_fd_sc_hd__dfxtp_1_544/CLK sky130_fd_sc_hd__nor2b_1_139/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_199 sky130_fd_sc_hd__xor2_1_199/B sky130_fd_sc_hd__xor2_1_199/X
+ sky130_fd_sc_hd__xor2_1_199/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_104 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_49/A1 sky130_fd_sc_hd__clkbuf_1_104/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_115 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_115/X sky130_fd_sc_hd__clkinv_1_990/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_126 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_126/X sky130_fd_sc_hd__clkinv_2_2/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_137 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_137/X sky130_fd_sc_hd__clkinv_1_891/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_208 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__buf_4_6/X
+ sky130_fd_sc_hd__buf_4_1/X sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__nor2_2_5/A
+ sky130_fd_sc_hd__o21ai_1_382/B1 sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_148 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_41/A1 sky130_fd_sc_hd__clkbuf_1_148/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o21ai_1_840 vssd1 vccd1 sky130_fd_sc_hd__inv_2_49/Y sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_840/B1 sky130_fd_sc_hd__xor2_1_613/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_219 vccd1 vssd1 sky130_fd_sc_hd__and3_4_16/X sky130_fd_sc_hd__and2_0_45/A
+ sky130_fd_sc_hd__and2_0_87/A sky130_fd_sc_hd__nor2_2_19/Y sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__o21ai_1_408/B1 sky130_fd_sc_hd__nor2b_2_3/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_159 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_31/A1 sky130_fd_sc_hd__clkbuf_1_159/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_6 sky130_fd_sc_hd__dfxtp_1_6/Q sky130_fd_sc_hd__dfxtp_1_8/CLK
+ la_data_out[63] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_851 vssd1 vccd1 sky130_fd_sc_hd__buf_2_13/X sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_851/B1 sky130_fd_sc_hd__xor2_1_625/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_862 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_640/A sky130_fd_sc_hd__nor2_1_221/Y
+ sky130_fd_sc_hd__nand2_1_665/Y sky130_fd_sc_hd__xnor2_1_188/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_873 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_651/A sky130_fd_sc_hd__nor2_1_232/Y
+ sky130_fd_sc_hd__nand2_1_709/Y sky130_fd_sc_hd__xnor2_1_199/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_884 vssd1 vccd1 sky130_fd_sc_hd__nand2_1_774/Y sky130_fd_sc_hd__a21oi_1_164/Y
+ sky130_fd_sc_hd__a21oi_1_163/Y sky130_fd_sc_hd__o21ai_1_884/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_895 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_678/A sky130_fd_sc_hd__nor2_1_256/Y
+ sky130_fd_sc_hd__nand2_1_801/Y sky130_fd_sc_hd__xnor2_1_292/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__inv_4_16 sky130_fd_sc_hd__inv_4_16/Y wbs_dat_i[18] vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__and2_0_102 vccd1 vssd1 sky130_fd_sc_hd__and2_0_102/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_102/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_10 la_data_out[117] sky130_fd_sc_hd__conb_1_132/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_113 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_65/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_113/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_21 la_data_out[106] sky130_fd_sc_hd__conb_1_121/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_124 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_35/D sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_124/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_32 la_data_out[31] sky130_fd_sc_hd__conb_1_110/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_8_4 sky130_fd_sc_hd__nand2_8_4/A sky130_fd_sc_hd__nand2_8_4/B
+ sky130_fd_sc_hd__buf_2_4/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_8
Xsky130_fd_sc_hd__and2_0_135 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_37/D sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_135/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_43 la_data_out[20] sky130_fd_sc_hd__conb_1_99/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_146 vccd1 vssd1 sky130_fd_sc_hd__and2_0_146/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_146/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_54 la_data_out[9] sky130_fd_sc_hd__conb_1_88/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_157 vccd1 vssd1 sky130_fd_sc_hd__and2_0_157/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_157/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_65 io_out[36] sky130_fd_sc_hd__conb_1_77/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_168 vccd1 vssd1 sky130_fd_sc_hd__and2_0_168/X sky130_fd_sc_hd__o21ai_2_0/B1
+ sky130_fd_sc_hd__and2_0_168/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_76 io_out[25] sky130_fd_sc_hd__conb_1_66/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_179 vccd1 vssd1 sky130_fd_sc_hd__and2_0_179/X sky130_fd_sc_hd__o21ai_2_0/B1
+ sky130_fd_sc_hd__o21ai_1_98/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_87 io_out[14] sky130_fd_sc_hd__conb_1_55/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_98 io_out[3] sky130_fd_sc_hd__conb_1_44/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_1 sky130_fd_sc_hd__nand2_1_7/B sky130_fd_sc_hd__mux2_2_22/X
+ sky130_fd_sc_hd__buf_4_4/A sky130_fd_sc_hd__mux2_2_42/X sky130_fd_sc_hd__nand2_1_8/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_80 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__buf_4_39/X
+ sky130_fd_sc_hd__a22o_1_80/X sky130_fd_sc_hd__a22o_1_80/B2 sky130_fd_sc_hd__nor2_1_269/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__o21ai_1_103 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_105/A2 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_119/Y sky130_fd_sc_hd__and2_0_173/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_114 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_117/A2 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_124/Y sky130_fd_sc_hd__and2_0_160/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_125 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_125/A2 sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__a22oi_1_173/Y sky130_fd_sc_hd__and2_0_146/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_136 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_137/A2 sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__a22oi_1_178/Y sky130_fd_sc_hd__and2_0_133/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_147 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_149/A2 sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__a22oi_1_185/Y sky130_fd_sc_hd__and2_0_118/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_158 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__o21ai_1_160/A1
+ sky130_fd_sc_hd__nand2_1_146/Y sky130_fd_sc_hd__and2_0_104/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_169 vssd1 vccd1 sky130_fd_sc_hd__inv_2_15/Y sky130_fd_sc_hd__nand2b_1_3/Y
+ sky130_fd_sc_hd__a222oi_1_51/Y sky130_fd_sc_hd__xor2_1_3/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nand2_1_507 sky130_fd_sc_hd__or2_0_55/A sky130_fd_sc_hd__nor2_1_165/Y
+ sky130_fd_sc_hd__nor2_1_172/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_518 sky130_fd_sc_hd__nand2_1_518/Y sky130_fd_sc_hd__nor2_1_169/Y
+ sky130_fd_sc_hd__nand2_1_546/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_529 sky130_fd_sc_hd__nand2_1_529/Y sky130_fd_sc_hd__nor2_1_172/Y
+ sky130_fd_sc_hd__nand2_1_546/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_9 sky130_fd_sc_hd__and3_4_13/C sky130_fd_sc_hd__nor2b_1_9/Y
+ sky130_fd_sc_hd__nor2b_1_9/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1109 sky130_fd_sc_hd__clkinv_4_52/A sky130_fd_sc_hd__a22o_1_29/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_70 sky130_fd_sc_hd__nand2_1_70/Y sky130_fd_sc_hd__nand2_1_70/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_81 sky130_fd_sc_hd__nand2_1_81/Y sky130_fd_sc_hd__nand2_1_81/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_92 sky130_fd_sc_hd__nand2_1_92/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__xor2_1_255/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_303 sky130_fd_sc_hd__dfxtp_1_303/Q sky130_fd_sc_hd__clkinv_8_6/Y
+ sky130_fd_sc_hd__and2_0_279/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_314 sky130_fd_sc_hd__nor2_1_239/A sky130_fd_sc_hd__dfxtp_1_319/CLK
+ sky130_fd_sc_hd__and2_0_291/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_325 sky130_fd_sc_hd__dfxtp_1_325/Q sky130_fd_sc_hd__dfxtp_1_343/CLK
+ sky130_fd_sc_hd__and2_0_320/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_336 sky130_fd_sc_hd__a22oi_1_9/B2 sky130_fd_sc_hd__dfxtp_1_339/CLK
+ sky130_fd_sc_hd__and2_0_326/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_347 sky130_fd_sc_hd__dfxtp_1_347/Q sky130_fd_sc_hd__dfxtp_1_356/CLK
+ sky130_fd_sc_hd__and2_0_310/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_358 sky130_fd_sc_hd__dfxtp_1_358/Q sky130_fd_sc_hd__dfxtp_2_7/CLK
+ sky130_fd_sc_hd__ha_2_8/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_369 sky130_fd_sc_hd__dfxtp_1_369/Q sky130_fd_sc_hd__dfxtp_1_371/CLK
+ sky130_fd_sc_hd__nor2b_1_114/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_670 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_767/A2 sky130_fd_sc_hd__nand2b_2_6/Y
+ sky130_fd_sc_hd__o21ai_1_670/B1 sky130_fd_sc_hd__xor2_1_453/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_681 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_681/A2 sky130_fd_sc_hd__nor2_1_173/Y
+ sky130_fd_sc_hd__nand2_1_532/Y sky130_fd_sc_hd__o21ai_1_681/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_208 sky130_fd_sc_hd__or2_0_30/A sky130_fd_sc_hd__nor2_2_12/B
+ sky130_fd_sc_hd__fa_2_208/A sky130_fd_sc_hd__fa_2_208/B sky130_fd_sc_hd__fa_2_208/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o21ai_1_692 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_10/X sky130_fd_sc_hd__nand2_1_529/Y
+ sky130_fd_sc_hd__a21oi_1_112/Y sky130_fd_sc_hd__xnor2_1_139/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_219 sky130_fd_sc_hd__fa_2_215/B sky130_fd_sc_hd__fa_2_222/CIN
+ sky130_fd_sc_hd__fa_2_219/A sky130_fd_sc_hd__fa_2_219/B sky130_fd_sc_hd__fa_2_219/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_11 sky130_fd_sc_hd__fa_2_1/A sky130_fd_sc_hd__fa_2_14/CIN sky130_fd_sc_hd__fa_2_11/A
+ sky130_fd_sc_hd__fa_2_11/B sky130_fd_sc_hd__xor2_1_27/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_22 sky130_fd_sc_hd__fa_2_11/A sky130_fd_sc_hd__fa_2_21/B sky130_fd_sc_hd__fa_2_22/A
+ sky130_fd_sc_hd__fa_2_22/B sky130_fd_sc_hd__xor2_1_36/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_33 sky130_fd_sc_hd__fa_2_18/B sky130_fd_sc_hd__fa_2_35/CIN
+ sky130_fd_sc_hd__fa_2_33/A sky130_fd_sc_hd__fa_2_33/B sky130_fd_sc_hd__fa_2_34/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_44 sky130_fd_sc_hd__fa_2_41/CIN sky130_fd_sc_hd__fa_2_51/A
+ sky130_fd_sc_hd__fa_2_44/A sky130_fd_sc_hd__fa_2_44/B sky130_fd_sc_hd__fa_2_48/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_55 sky130_fd_sc_hd__fa_2_51/B sky130_fd_sc_hd__fa_2_59/CIN
+ sky130_fd_sc_hd__fa_2_55/A sky130_fd_sc_hd__fa_2_55/B sky130_fd_sc_hd__fa_2_55/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_66 sky130_fd_sc_hd__or2_0_3/A sky130_fd_sc_hd__nor2_1_62/B
+ sky130_fd_sc_hd__fa_2_66/A sky130_fd_sc_hd__fa_2_66/B sky130_fd_sc_hd__fa_2_66/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_77 sky130_fd_sc_hd__fa_2_73/B sky130_fd_sc_hd__fa_2_80/CIN
+ sky130_fd_sc_hd__fa_2_77/A sky130_fd_sc_hd__fa_2_77/B sky130_fd_sc_hd__fa_2_77/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_88 sky130_fd_sc_hd__fa_2_84/B sky130_fd_sc_hd__fa_2_89/B sky130_fd_sc_hd__fa_2_88/A
+ sky130_fd_sc_hd__fa_2_88/B sky130_fd_sc_hd__fa_2_88/CIN vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_99 sky130_fd_sc_hd__fa_2_96/CIN sky130_fd_sc_hd__fa_2_99/SUM
+ sky130_fd_sc_hd__fa_2_99/A sky130_fd_sc_hd__fa_2_99/B sky130_fd_sc_hd__fa_2_99/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_203 vccd1 vssd1 sky130_fd_sc_hd__buf_2_203/X sky130_fd_sc_hd__buf_2_203/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_214 vccd1 vssd1 sky130_fd_sc_hd__buf_2_214/X sky130_fd_sc_hd__mux2_4_5/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__a222oi_1_550 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_420/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_452/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_747/A sky130_fd_sc_hd__dfxtp_1_388/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a21oi_1_16 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_45/Y
+ sky130_fd_sc_hd__a21oi_1_16/Y sky130_fd_sc_hd__dfxtp_1_81/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_561 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_409/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_441/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_758/A sky130_fd_sc_hd__dfxtp_1_377/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a21oi_1_27 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_56/Y
+ sky130_fd_sc_hd__a21oi_1_27/Y sky130_fd_sc_hd__dfxtp_1_70/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_572 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_398/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_430/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_769/A sky130_fd_sc_hd__dfxtp_1_366/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a21oi_1_38 sky130_fd_sc_hd__a21oi_1_45/A1 sky130_fd_sc_hd__o21ai_1_188/Y
+ sky130_fd_sc_hd__a21oi_1_38/Y sky130_fd_sc_hd__nor2_1_47/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_583 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_405/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_437/Q sky130_fd_sc_hd__clkbuf_1_32/X
+ sky130_fd_sc_hd__clkinv_1_780/A sky130_fd_sc_hd__dfxtp_1_373/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a21oi_1_49 sky130_fd_sc_hd__nand2_1_250/Y sky130_fd_sc_hd__nand2_1_240/Y
+ sky130_fd_sc_hd__a21oi_1_49/Y sky130_fd_sc_hd__nor2_1_75/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_594 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_399/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_431/Q sky130_fd_sc_hd__clkbuf_1_32/X
+ sky130_fd_sc_hd__clkinv_1_791/A sky130_fd_sc_hd__dfxtp_1_367/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_12 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_23 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_34 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_45 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_150 sky130_fd_sc_hd__clkinv_4_69/Y sky130_fd_sc_hd__nor2b_1_150/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__decap_12_56 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_67 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_78 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_89 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_12 vccd1 vssd1 sky130_fd_sc_hd__buf_6_12/X sky130_fd_sc_hd__buf_6_12/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_23 vccd1 vssd1 sky130_fd_sc_hd__buf_6_23/X sky130_fd_sc_hd__buf_6_23/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_34 vccd1 vssd1 sky130_fd_sc_hd__buf_6_34/X sky130_fd_sc_hd__buf_8_3/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_45 vccd1 vssd1 sky130_fd_sc_hd__buf_6_45/X sky130_fd_sc_hd__buf_8_77/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_56 vccd1 vssd1 sky130_fd_sc_hd__buf_6_56/X sky130_fd_sc_hd__buf_8_12/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_67 vccd1 vssd1 sky130_fd_sc_hd__buf_6_67/X sky130_fd_sc_hd__buf_8_98/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_78 vccd1 vssd1 sky130_fd_sc_hd__buf_6_78/X sky130_fd_sc_hd__buf_8_80/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_89 vccd1 vssd1 sky130_fd_sc_hd__buf_6_89/X sky130_fd_sc_hd__buf_6_89/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_14 sky130_fd_sc_hd__clkinv_4_66/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_25 sky130_fd_sc_hd__clkinv_4_61/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_36 sky130_fd_sc_hd__clkinv_4_53/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_47 sky130_fd_sc_hd__buf_2_189/A vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_58 sky130_fd_sc_hd__buf_2_192/A vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_69 la_data_out[62] vssd1 vccd1 vccd1 vssd1 sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__decap_12_409 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_304 sky130_fd_sc_hd__xnor2_1_57/A sky130_fd_sc_hd__nand2_1_305/Y
+ sky130_fd_sc_hd__or2_0_22/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_903 sky130_fd_sc_hd__clkinv_1_903/Y sky130_fd_sc_hd__clkinv_4_90/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_315 sky130_fd_sc_hd__xnor2_1_4/A sky130_fd_sc_hd__nand2_1_316/Y
+ sky130_fd_sc_hd__or2_0_26/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_914 sky130_fd_sc_hd__clkinv_1_914/Y sky130_fd_sc_hd__inv_2_200/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_326 sky130_fd_sc_hd__nand2_1_326/Y sky130_fd_sc_hd__nor2_1_130/Y
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_925 sky130_fd_sc_hd__clkinv_1_927/A sky130_fd_sc_hd__a21o_2_3/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_337 sky130_fd_sc_hd__nand2_1_337/Y sky130_fd_sc_hd__or2_0_9/A
+ sky130_fd_sc_hd__or2_0_4/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_936 sky130_fd_sc_hd__clkinv_1_937/A sky130_fd_sc_hd__inv_2_126/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_348 sky130_fd_sc_hd__xnor2_1_72/A sky130_fd_sc_hd__nand2_1_349/Y
+ sky130_fd_sc_hd__or2_0_38/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_947 sky130_fd_sc_hd__buf_8_132/A sky130_fd_sc_hd__inv_2_145/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_359 sky130_fd_sc_hd__xnor2_1_76/A sky130_fd_sc_hd__nand2_1_360/Y
+ sky130_fd_sc_hd__nand2_1_359/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_958 sky130_fd_sc_hd__clkinv_2_29/A sky130_fd_sc_hd__buf_2_143/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_969 sky130_fd_sc_hd__buf_2_129/A sky130_fd_sc_hd__clkinv_4_22/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_100 sky130_fd_sc_hd__dfxtp_1_100/Q sky130_fd_sc_hd__dfxtp_1_105/CLK
+ sky130_fd_sc_hd__and2_0_127/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1408 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_111 sky130_fd_sc_hd__dfxtp_1_111/Q sky130_fd_sc_hd__dfxtp_1_97/CLK
+ sky130_fd_sc_hd__and2_0_171/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1419 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_122 sky130_fd_sc_hd__dfxtp_1_122/Q sky130_fd_sc_hd__dfxtp_1_122/CLK
+ sky130_fd_sc_hd__and2_0_238/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_133 sky130_fd_sc_hd__dfxtp_1_133/Q sky130_fd_sc_hd__dfxtp_1_138/CLK
+ sky130_fd_sc_hd__and2_0_136/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_144 sky130_fd_sc_hd__dfxtp_1_144/Q sky130_fd_sc_hd__dfxtp_1_146/CLK
+ sky130_fd_sc_hd__and2_0_191/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_155 sky130_fd_sc_hd__dfxtp_1_155/Q sky130_fd_sc_hd__dfxtp_1_158/CLK
+ sky130_fd_sc_hd__and2_0_246/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_166 sky130_fd_sc_hd__dfxtp_1_166/Q sky130_fd_sc_hd__dfxtp_1_170/CLK
+ sky130_fd_sc_hd__and2_0_138/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_177 sky130_fd_sc_hd__dfxtp_1_177/Q sky130_fd_sc_hd__dfxtp_1_177/CLK
+ sky130_fd_sc_hd__and2_0_193/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_188 sky130_fd_sc_hd__dfxtp_1_188/Q sky130_fd_sc_hd__dfxtp_1_190/CLK
+ sky130_fd_sc_hd__and2_0_8/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_199 sky130_fd_sc_hd__xnor2_1_171/A sky130_fd_sc_hd__dfxtp_2_2/CLK
+ sky130_fd_sc_hd__and2_0_41/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_910 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_921 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_932 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_943 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_954 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_965 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_976 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_860 sky130_fd_sc_hd__o31ai_1_0/A1 sky130_fd_sc_hd__o21ai_1_919/Y
+ sky130_fd_sc_hd__nand2_1_860/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_987 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_998 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o211ai_1_19 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_44/B1
+ sky130_fd_sc_hd__o211ai_1_19/Y sky130_fd_sc_hd__a22oi_1_70/Y sky130_fd_sc_hd__a22oi_1_71/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o21ai_1_60 vssd1 vccd1 sky130_fd_sc_hd__inv_2_60/Y sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_60/B1 sky130_fd_sc_hd__o21ai_1_60/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_71 vssd1 vccd1 sky130_fd_sc_hd__inv_2_57/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__o21ai_1_71/B1 sky130_fd_sc_hd__o21ai_1_71/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_82 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_85/A2 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__o21ai_1_82/B1 sky130_fd_sc_hd__o21ai_1_82/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_93 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_93/A2 sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__o21ai_1_93/B1 sky130_fd_sc_hd__o21ai_1_93/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_380 vccd1 vssd1 sky130_fd_sc_hd__and3_4_23/X sky130_fd_sc_hd__buf_4_7/X
+ sky130_fd_sc_hd__buf_4_0/X sky130_fd_sc_hd__nor2_1_178/Y sky130_fd_sc_hd__buf_2_23/X
+ sky130_fd_sc_hd__o21ai_1_640/B1 sky130_fd_sc_hd__nor2b_1_15/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_391 vccd1 vssd1 sky130_fd_sc_hd__and3_4_24/X sky130_fd_sc_hd__buf_2_23/X
+ sky130_fd_sc_hd__buf_2_31/X sky130_fd_sc_hd__nor2_1_183/Y sky130_fd_sc_hd__buf_2_4/A
+ sky130_fd_sc_hd__o21ai_1_654/B1 sky130_fd_sc_hd__nor2b_1_16/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a21oi_1_107 sky130_fd_sc_hd__o21ai_1_693/Y sky130_fd_sc_hd__o21ai_1_651/Y
+ sky130_fd_sc_hd__o21a_1_4/B1 sky130_fd_sc_hd__nor2_1_165/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_118 sky130_fd_sc_hd__nand2_1_572/Y sky130_fd_sc_hd__nor2_1_181/A
+ sky130_fd_sc_hd__a21oi_1_118/Y sky130_fd_sc_hd__or2_0_63/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_129 sky130_fd_sc_hd__nor2_1_205/Y sky130_fd_sc_hd__o21ai_1_834/Y
+ sky130_fd_sc_hd__xor2_1_602/A sky130_fd_sc_hd__o21ai_1_839/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_500 sky130_fd_sc_hd__buf_12_500/A sky130_fd_sc_hd__buf_12_581/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_511 sky130_fd_sc_hd__buf_12_511/A sky130_fd_sc_hd__buf_12_511/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_522 sky130_fd_sc_hd__buf_12_522/A sky130_fd_sc_hd__buf_12_522/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_533 sky130_fd_sc_hd__buf_12_533/A sky130_fd_sc_hd__buf_12_533/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_544 sky130_fd_sc_hd__buf_12_544/A sky130_fd_sc_hd__buf_12_544/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_555 sky130_fd_sc_hd__buf_12_555/A sky130_fd_sc_hd__buf_12_555/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_566 sky130_fd_sc_hd__buf_12_566/A sky130_fd_sc_hd__buf_12_566/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_8_3 sky130_fd_sc_hd__buf_12_66/A sky130_fd_sc_hd__buf_8_69/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_8
Xsky130_fd_sc_hd__buf_12_577 sky130_fd_sc_hd__buf_12_577/A sky130_fd_sc_hd__buf_12_577/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_206 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_588 sky130_fd_sc_hd__buf_12_588/A sky130_fd_sc_hd__buf_12_588/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_217 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_599 sky130_fd_sc_hd__buf_12_599/A sky130_fd_sc_hd__buf_12_599/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__nand2_1_101 sky130_fd_sc_hd__o21ai_1_67/B1 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__xor2_1_296/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_228 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_700 sky130_fd_sc_hd__nand2_1_789/A sky130_fd_sc_hd__ha_2_9/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_112 sky130_fd_sc_hd__o21ai_1_90/B1 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__xor2_1_346/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_239 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_711 sky130_fd_sc_hd__nor2b_1_90/A sky130_fd_sc_hd__fa_2_462/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_123 sky130_fd_sc_hd__nand2_1_123/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_123/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_722 sky130_fd_sc_hd__nor2b_1_101/A sky130_fd_sc_hd__xnor2_1_294/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_134 sky130_fd_sc_hd__nand2_1_134/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_135/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_733 sky130_fd_sc_hd__nor2b_1_112/A sky130_fd_sc_hd__xor2_1_685/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_145 sky130_fd_sc_hd__nand2_1_145/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__xor2_1_421/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_744 sky130_fd_sc_hd__fa_2_467/A sky130_fd_sc_hd__clkinv_1_744/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_307 vssd1 vccd1 sky130_fd_sc_hd__ha_2_51/SUM sky130_fd_sc_hd__xnor2_1_307/Y
+ la_data_out[46] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_156 sky130_fd_sc_hd__nand2_1_156/Y sky130_fd_sc_hd__nor2_1_72/Y
+ sky130_fd_sc_hd__clkbuf_1_3/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_755 sky130_fd_sc_hd__fa_2_478/A sky130_fd_sc_hd__clkinv_1_755/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_167 sky130_fd_sc_hd__nand2_1_167/Y sky130_fd_sc_hd__nand2_1_168/Y
+ sky130_fd_sc_hd__or2_0_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_766 sky130_fd_sc_hd__fa_2_489/A sky130_fd_sc_hd__clkinv_1_766/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_178 sky130_fd_sc_hd__nand2_1_178/Y sky130_fd_sc_hd__or2_0_58/A
+ sky130_fd_sc_hd__or2_0_9/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_777 sky130_fd_sc_hd__and2_0_330/A sky130_fd_sc_hd__clkinv_1_777/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_189 sky130_fd_sc_hd__nand2_1_189/Y sky130_fd_sc_hd__or2_0_58/B
+ sky130_fd_sc_hd__or2_0_42/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_788 sky130_fd_sc_hd__and2_0_319/A sky130_fd_sc_hd__clkinv_1_788/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_799 sky130_fd_sc_hd__and2_0_308/A sky130_fd_sc_hd__clkinv_1_799/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1205 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_5 sky130_fd_sc_hd__fa_2_75/A sky130_fd_sc_hd__xor3_1_8/C
+ sky130_fd_sc_hd__xor2_1_5/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1216 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1227 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1238 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1249 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_8_3 sky130_fd_sc_hd__clkinv_8_3/Y sky130_fd_sc_hd__clkinv_8_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_12_740 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_751 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_762 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_773 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_784 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_795 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_507 sky130_fd_sc_hd__fa_2_379/A sky130_fd_sc_hd__fa_2_335/B
+ sky130_fd_sc_hd__xor2_1_507/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_690 sky130_fd_sc_hd__xnor2_1_195/A sky130_fd_sc_hd__nand2_1_691/Y
+ sky130_fd_sc_hd__or2_0_79/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_518 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__xor2_1_518/X
+ sky130_fd_sc_hd__xor2_1_518/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_529 sky130_fd_sc_hd__fa_2_357/A sky130_fd_sc_hd__xor2_1_529/X
+ sky130_fd_sc_hd__xor2_1_529/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1750 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1761 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_60 sky130_fd_sc_hd__inv_2_60/A sky130_fd_sc_hd__inv_2_60/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1772 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_71 sky130_fd_sc_hd__inv_2_71/A sky130_fd_sc_hd__inv_2_71/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1783 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_82 la_data_out[45] sky130_fd_sc_hd__inv_4_9/A vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1794 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_93 sky130_fd_sc_hd__inv_2_93/A sky130_fd_sc_hd__inv_2_93/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__ha_2_14 vssd1 vccd1 sky130_fd_sc_hd__ha_2_14/A sky130_fd_sc_hd__or2_0_96/A
+ sky130_fd_sc_hd__ha_2_14/SUM sky130_fd_sc_hd__ha_2_14/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_25 vssd1 vccd1 la_data_out[58] sky130_fd_sc_hd__ha_2_24/B sky130_fd_sc_hd__ha_2_25/SUM
+ la_data_out[57] vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_36 vssd1 vccd1 sky130_fd_sc_hd__ha_2_36/A sky130_fd_sc_hd__ha_2_35/B
+ sky130_fd_sc_hd__ha_2_36/SUM sky130_fd_sc_hd__ha_2_36/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_47 vssd1 vccd1 sky130_fd_sc_hd__ha_2_47/A sky130_fd_sc_hd__ha_2_50/B
+ sky130_fd_sc_hd__ha_2_47/SUM sky130_fd_sc_hd__ha_2_47/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__and2b_4_9 sky130_fd_sc_hd__or2b_2_2/A sky130_fd_sc_hd__and2b_4_9/X
+ sky130_fd_sc_hd__and3_4_19/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__and2b_4
Xsky130_fd_sc_hd__ha_2_58 vssd1 vccd1 sky130_fd_sc_hd__ha_2_58/A sky130_fd_sc_hd__ha_2_58/COUT
+ sky130_fd_sc_hd__ha_2_58/SUM sky130_fd_sc_hd__ha_2_58/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__sdlclkp_4_10 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_4_1/Y
+ sky130_fd_sc_hd__dfxtp_1_99/CLK sky130_fd_sc_hd__clkbuf_1_11/X vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_380 sky130_fd_sc_hd__fa_2_378/CIN sky130_fd_sc_hd__fa_2_381/CIN
+ sky130_fd_sc_hd__fa_2_380/A sky130_fd_sc_hd__fa_2_380/B sky130_fd_sc_hd__xor2_1_560/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_21 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_8_61/Y
+ sky130_fd_sc_hd__dfxtp_2_2/CLK sky130_fd_sc_hd__o21ai_2_2/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_391 sky130_fd_sc_hd__fa_2_386/A sky130_fd_sc_hd__fa_2_390/B
+ sky130_fd_sc_hd__fa_2_391/A sky130_fd_sc_hd__fa_2_391/B sky130_fd_sc_hd__fa_2_391/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_32 sky130_fd_sc_hd__conb_1_145/LO sky130_fd_sc_hd__clkinv_2_11/A
+ sky130_fd_sc_hd__dfxtp_1_339/CLK sky130_fd_sc_hd__nand4_1_1/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_43 sky130_fd_sc_hd__conb_1_145/LO sky130_fd_sc_hd__clkinv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_423/CLK sky130_fd_sc_hd__o21ai_1_891/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_54 sky130_fd_sc_hd__conb_1_149/LO sky130_fd_sc_hd__clkinv_4_117/A
+ sky130_fd_sc_hd__dfxtp_1_552/CLK sky130_fd_sc_hd__or2_0_113/X vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_101 sky130_fd_sc_hd__buf_4_1/X sky130_fd_sc_hd__nor2_1_44/B
+ sky130_fd_sc_hd__buf_4_6/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_112 sky130_fd_sc_hd__nor2_1_113/B sky130_fd_sc_hd__nor2_1_112/Y
+ sky130_fd_sc_hd__nor2_1_112/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_123 sky130_fd_sc_hd__nor2_1_126/A sky130_fd_sc_hd__nor2_1_123/Y
+ sky130_fd_sc_hd__nor2_1_123/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_10 sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__dfxtp_1_286/Q sky130_fd_sc_hd__o211ai_1_10/Y sky130_fd_sc_hd__nand2_1_12/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_134 sky130_fd_sc_hd__nor2_1_134/B sky130_fd_sc_hd__nor2_1_134/Y
+ sky130_fd_sc_hd__nor2_1_137/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_145 sky130_fd_sc_hd__nor2_1_145/B sky130_fd_sc_hd__nor2_1_145/Y
+ sky130_fd_sc_hd__nor2_1_145/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_21 sky130_fd_sc_hd__nor2_4_0/Y sky130_fd_sc_hd__nor2_2_0/Y
+ sky130_fd_sc_hd__dfxtp_1_330/Q sky130_fd_sc_hd__or2_0_91/A sky130_fd_sc_hd__nand2_1_15/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_156 sky130_fd_sc_hd__nor2_1_159/Y sky130_fd_sc_hd__nor2_1_156/Y
+ sky130_fd_sc_hd__nor2_1_157/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_32 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__clkbuf_1_25/X
+ sky130_fd_sc_hd__nand2_1_81/B sky130_fd_sc_hd__dfxtp_1_127/Q sky130_fd_sc_hd__a22oi_1_32/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_43 sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__dfxtp_1_100/Q sky130_fd_sc_hd__dfxtp_1_68/Q sky130_fd_sc_hd__a22oi_1_43/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_167 sky130_fd_sc_hd__nor2_1_167/B sky130_fd_sc_hd__nor2_1_167/Y
+ sky130_fd_sc_hd__nor2_1_167/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_178 sky130_fd_sc_hd__and3_4_23/A sky130_fd_sc_hd__nor2_1_178/Y
+ sky130_fd_sc_hd__and3_4_23/C vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_54 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__nor2_4_3/Y
+ sky130_fd_sc_hd__nand2_1_72/B sky130_fd_sc_hd__dfxtp_1_138/Q sky130_fd_sc_hd__a22oi_1_54/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_65 sky130_fd_sc_hd__clkbuf_1_24/X sky130_fd_sc_hd__clkbuf_1_23/X
+ sky130_fd_sc_hd__dfxtp_1_111/Q sky130_fd_sc_hd__dfxtp_1_79/Q sky130_fd_sc_hd__a22oi_1_65/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_189 sky130_fd_sc_hd__nor2_1_193/Y sky130_fd_sc_hd__nor2_1_189/Y
+ sky130_fd_sc_hd__nor2_1_191/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_76 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__nor2_4_3/Y
+ sky130_fd_sc_hd__nand2_1_61/B sky130_fd_sc_hd__dfxtp_1_149/Q sky130_fd_sc_hd__a22oi_1_76/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_87 sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__dfxtp_1_122/Q sky130_fd_sc_hd__dfxtp_1_90/Q sky130_fd_sc_hd__a22oi_1_87/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_98 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_186/Q sky130_fd_sc_hd__dfxtp_1_154/Q sky130_fd_sc_hd__o21ai_1_4/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_330 sky130_fd_sc_hd__buf_12_330/A sky130_fd_sc_hd__buf_12_537/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_341 sky130_fd_sc_hd__buf_12_341/A sky130_fd_sc_hd__buf_12_663/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_200 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__and2b_4_1/X sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__a22oi_1_200/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_352 sky130_fd_sc_hd__buf_12_352/A sky130_fd_sc_hd__buf_12_562/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_211 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__and2b_4_5/X sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__a22oi_1_211/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_363 sky130_fd_sc_hd__buf_12_363/A sky130_fd_sc_hd__buf_12_648/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_222 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__and2b_4_9/X sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__a22oi_1_222/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_374 sky130_fd_sc_hd__buf_12_374/A sky130_fd_sc_hd__buf_12_560/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_385 sky130_fd_sc_hd__buf_12_60/X sky130_fd_sc_hd__buf_12_497/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_396 sky130_fd_sc_hd__buf_12_81/X sky130_fd_sc_hd__buf_12_600/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_530 sky130_fd_sc_hd__o21ai_1_679/A2 sky130_fd_sc_hd__xnor2_1_137/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_541 sky130_fd_sc_hd__o21ai_1_713/A2 sky130_fd_sc_hd__xnor2_1_143/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_104 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_104/B sky130_fd_sc_hd__xnor2_1_104/Y
+ sky130_fd_sc_hd__xnor2_1_104/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_552 sky130_fd_sc_hd__o21ai_1_733/A2 sky130_fd_sc_hd__xnor2_1_148/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_115 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_115/B sky130_fd_sc_hd__inv_2_34/A
+ sky130_fd_sc_hd__xnor2_1_115/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_563 sky130_fd_sc_hd__o21ai_1_767/A2 sky130_fd_sc_hd__xnor2_1_155/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_126 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_126/B sky130_fd_sc_hd__xnor2_1_126/Y
+ sky130_fd_sc_hd__xnor2_1_126/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_574 sky130_fd_sc_hd__clkinv_1_574/Y sky130_fd_sc_hd__nand2_1_592/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_137 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_137/B sky130_fd_sc_hd__xnor2_1_137/Y
+ sky130_fd_sc_hd__xnor2_1_137/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_585 sky130_fd_sc_hd__clkinv_1_585/Y sky130_fd_sc_hd__nand2_1_616/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_148 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_148/B sky130_fd_sc_hd__xnor2_1_148/Y
+ sky130_fd_sc_hd__xnor2_1_148/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_596 sky130_fd_sc_hd__xor2_1_612/B sky130_fd_sc_hd__o21ai_1_839/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_4_10 sky130_fd_sc_hd__clkinv_8_7/Y sky130_fd_sc_hd__clkinv_4_11/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__xnor2_1_159 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_159/B sky130_fd_sc_hd__xnor2_1_159/Y
+ sky130_fd_sc_hd__xnor2_1_159/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_4_21 sky130_fd_sc_hd__clkinv_4_21/A sky130_fd_sc_hd__clkinv_4_21/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_32 sky130_fd_sc_hd__nand2_1_12/Y sky130_fd_sc_hd__inv_2_156/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_43 sky130_fd_sc_hd__clkinv_4_43/A sky130_fd_sc_hd__buf_12_77/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_54 sky130_fd_sc_hd__clkinv_4_54/A sky130_fd_sc_hd__clkinv_4_54/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_65 sky130_fd_sc_hd__clkinv_4_65/A sky130_fd_sc_hd__clkinv_4_65/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_76 sky130_fd_sc_hd__clkinv_4_76/A sky130_fd_sc_hd__clkinv_4_76/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_1002 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_4_87 wbs_dat_i[16] sky130_fd_sc_hd__clkinv_4_87/Y vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_1013 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_4_98 sky130_fd_sc_hd__clkinv_8_54/Y sky130_fd_sc_hd__clkinv_8_56/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_1024 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1035 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1046 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1057 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1068 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_16_6 sky130_fd_sc_hd__inv_16_6/Y sky130_fd_sc_hd__inv_16_6/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__decap_12_1079 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__and2b_4_13 sky130_fd_sc_hd__nor2_4_19/A sky130_fd_sc_hd__and2b_4_13/X
+ sky130_fd_sc_hd__nor2_4_19/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__and2b_4
Xsky130_fd_sc_hd__decap_12_570 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_581 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_592 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_304 sky130_fd_sc_hd__fa_2_239/A sky130_fd_sc_hd__fa_2_203/A
+ sky130_fd_sc_hd__xor2_1_304/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_315 sky130_fd_sc_hd__fa_2_239/A sky130_fd_sc_hd__fa_2_220/B
+ sky130_fd_sc_hd__xor2_1_315/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_326 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__xor2_1_326/X
+ sky130_fd_sc_hd__xor2_1_326/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_337 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__fa_2_229/A
+ sky130_fd_sc_hd__xor2_1_337/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_348 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__fa_2_241/B
+ sky130_fd_sc_hd__xor2_1_348/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_359 sky130_fd_sc_hd__xor2_1_359/B sky130_fd_sc_hd__xor2_1_359/X
+ sky130_fd_sc_hd__xor2_1_359/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_308 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_308/X sky130_fd_sc_hd__clkinv_1_858/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_12_1580 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_319 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_319/X sky130_fd_sc_hd__clkinv_1_859/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_12_1591 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_12 sky130_fd_sc_hd__dfxtp_1_12/Q sky130_fd_sc_hd__dfxtp_1_8/CLK
+ sky130_fd_sc_hd__dfxtp_1_12/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_23 sky130_fd_sc_hd__ha_2_3/A sky130_fd_sc_hd__dfxtp_1_29/CLK
+ sky130_fd_sc_hd__or4_1_3/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_34 sky130_fd_sc_hd__nand2_1_80/B sky130_fd_sc_hd__dfxtp_1_46/CLK
+ sky130_fd_sc_hd__dfxtp_1_34/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_45 sky130_fd_sc_hd__nand2_1_69/B sky130_fd_sc_hd__dfxtp_1_45/CLK
+ sky130_fd_sc_hd__dfxtp_1_45/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_56 sky130_fd_sc_hd__nand2_1_57/B sky130_fd_sc_hd__dfxtp_1_57/CLK
+ sky130_fd_sc_hd__dfxtp_1_56/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_67 sky130_fd_sc_hd__dfxtp_1_67/Q sky130_fd_sc_hd__dfxtp_1_72/CLK
+ sky130_fd_sc_hd__dfxtp_1_67/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_78 sky130_fd_sc_hd__dfxtp_1_78/Q sky130_fd_sc_hd__dfxtp_1_78/CLK
+ sky130_fd_sc_hd__dfxtp_1_78/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_89 sky130_fd_sc_hd__dfxtp_1_89/Q sky130_fd_sc_hd__dfxtp_1_89/CLK
+ sky130_fd_sc_hd__dfxtp_1_89/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_306 vccd1 vssd1 sky130_fd_sc_hd__and2_0_306/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_306/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_317 vccd1 vssd1 sky130_fd_sc_hd__and2_0_317/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_317/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_328 vccd1 vssd1 sky130_fd_sc_hd__and2_0_328/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_328/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_339 vccd1 vssd1 sky130_fd_sc_hd__and2_0_394/A sky130_fd_sc_hd__xor2_1_692/X
+ sky130_fd_sc_hd__and2_0_342/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__inv_2_106 sky130_fd_sc_hd__inv_2_107/A sky130_fd_sc_hd__inv_2_106/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_117 sky130_fd_sc_hd__inv_6_1/Y sky130_fd_sc_hd__buf_6_17/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__or2_0_8 sky130_fd_sc_hd__or2_0_8/A sky130_fd_sc_hd__or2_0_8/X sky130_fd_sc_hd__or2_0_8/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__inv_2_128 sky130_fd_sc_hd__inv_2_128/A sky130_fd_sc_hd__buf_6_18/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_139 sky130_fd_sc_hd__inv_2_139/A sky130_fd_sc_hd__buf_8_54/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_sram_1kbyte_1rw1r_32x256_8_2 sky130_fd_sc_hd__buf_2_128/X sky130_fd_sc_hd__buf_2_128/X
+ sky130_fd_sc_hd__buf_12_652/X sky130_fd_sc_hd__buf_12_621/X sky130_fd_sc_hd__buf_12_452/X
+ sky130_fd_sc_hd__buf_12_627/X sky130_fd_sc_hd__buf_12_344/X sky130_fd_sc_hd__buf_12_614/X
+ sky130_fd_sc_hd__buf_12_646/X sky130_fd_sc_hd__clkinv_1_967/Y sky130_fd_sc_hd__buf_12_612/X
+ sky130_fd_sc_hd__buf_12_522/X sky130_fd_sc_hd__buf_12_529/X vccd1 sky130_fd_sc_hd__clkinv_8_31/Y
+ sky130_fd_sc_hd__buf_2_112/A sky130_fd_sc_hd__buf_2_111/A sky130_fd_sc_hd__buf_2_110/A
+ sky130_fd_sc_hd__buf_2_109/A sky130_fd_sc_hd__buf_2_108/A sky130_fd_sc_hd__buf_2_107/A
+ sky130_fd_sc_hd__buf_2_106/A sky130_fd_sc_hd__buf_2_105/A sky130_fd_sc_hd__buf_2_104/A
+ sky130_fd_sc_hd__buf_2_103/A sky130_fd_sc_hd__buf_2_102/A sky130_fd_sc_hd__buf_2_101/A
+ sky130_fd_sc_hd__buf_2_100/A sky130_fd_sc_hd__buf_2_99/A sky130_fd_sc_hd__buf_2_98/A
+ sky130_fd_sc_hd__buf_2_97/A sky130_fd_sc_hd__buf_12_220/X sky130_fd_sc_hd__buf_2_126/A
+ sky130_fd_sc_hd__buf_2_125/A sky130_fd_sc_hd__buf_2_124/A sky130_fd_sc_hd__buf_2_123/A
+ sky130_fd_sc_hd__clkbuf_4_17/A sky130_fd_sc_hd__buf_2_122/A sky130_fd_sc_hd__buf_2_121/A
+ sky130_fd_sc_hd__buf_2_120/A sky130_fd_sc_hd__buf_2_119/A sky130_fd_sc_hd__buf_2_118/A
+ sky130_fd_sc_hd__buf_2_117/A sky130_fd_sc_hd__buf_2_116/A sky130_fd_sc_hd__buf_2_115/A
+ sky130_fd_sc_hd__buf_2_114/A sky130_fd_sc_hd__buf_2_113/A sky130_fd_sc_hd__buf_2_127/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[10] sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[11]
+ sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[12] sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[13]
+ sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[14] sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[15]
+ sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[16] sky130_fd_sc_hd__buf_12_542/X sky130_fd_sc_hd__buf_12_141/X
+ sky130_fd_sc_hd__buf_12_171/X sky130_fd_sc_hd__buf_12_303/X sky130_fd_sc_hd__buf_12_121/X
+ sky130_fd_sc_hd__dfxtp_1_9/CLK sky130_fd_sc_hd__clkinv_1_982/Y sky130_fd_sc_hd__buf_2_167/X
+ sky130_fd_sc_hd__clkinv_1_978/Y sky130_fd_sc_hd__clkinv_4_25/Y sky130_fd_sc_hd__clkinv_4_24/Y
+ sky130_fd_sc_hd__clkinv_1_975/Y sky130_fd_sc_hd__clkinv_1_972/Y sky130_fd_sc_hd__clkinv_1_971/Y
+ sky130_fd_sc_hd__inv_2_153/Y sky130_fd_sc_hd__clkinv_1_968/Y sky130_fd_sc_hd__clkinv_1_991/Y
+ sky130_fd_sc_hd__clkbuf_1_315/X sky130_fd_sc_hd__clkinv_1_987/Y sky130_fd_sc_hd__inv_2_154/Y
+ sky130_fd_sc_hd__clkinv_1_985/Y sky130_fd_sc_hd__clkinv_2_34/Y sky130_fd_sc_hd__clkbuf_1_132/X
+ sky130_fd_sc_hd__clkbuf_1_130/X sky130_fd_sc_hd__clkbuf_1_129/X sky130_fd_sc_hd__clkbuf_1_128/X
+ sky130_fd_sc_hd__buf_2_134/X sky130_fd_sc_hd__clkbuf_1_127/X sky130_fd_sc_hd__clkbuf_1_126/X
+ sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[0] sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[1]
+ sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[2] sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[3]
+ sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[4] sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[5]
+ sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[6] sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[7]
+ sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[8] sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[9]
+ sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[25] sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[26]
+ sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[27] sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[28]
+ sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[29] sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[30]
+ sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[31] sky130_fd_sc_hd__clkinv_1_992/Y sky130_fd_sc_hd__clkbuf_1_125/X
+ sky130_fd_sc_hd__clkbuf_1_123/X sky130_fd_sc_hd__clkbuf_1_122/X sky130_fd_sc_hd__clkbuf_1_121/X
+ sky130_fd_sc_hd__clkbuf_1_120/X sky130_fd_sc_hd__clkbuf_1_119/X sky130_fd_sc_hd__clkbuf_1_118/X
+ sky130_fd_sc_hd__clkbuf_1_116/X sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[17] sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[18]
+ sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[19] sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[20]
+ sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[21] sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[22]
+ sky130_fd_sc_hd__buf_12_520/X sky130_fd_sc_hd__buf_12_606/X sky130_fd_sc_hd__buf_12_525/X
+ sky130_fd_sc_hd__buf_12_556/X sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[23] sky130_sram_1kbyte_1rw1r_32x256_8_2/dout0[24]
+ sky130_sram_1kbyte_1rw1r_32x256_8_2/sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/gnd_uq26
+ vssd1 sky130_sram_1kbyte_1rw1r_32x256_8
Xsky130_fd_sc_hd__buf_12_160 sky130_fd_sc_hd__buf_12_31/X sky130_fd_sc_hd__buf_12_377/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_171 sky130_fd_sc_hd__buf_12_34/X sky130_fd_sc_hd__buf_12_171/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_182 sky130_fd_sc_hd__buf_12_54/X sky130_fd_sc_hd__buf_12_318/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_193 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__buf_12_400/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_360 sky130_fd_sc_hd__a21oi_2_5/B1 sky130_fd_sc_hd__nand2_1_233/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_371 sky130_fd_sc_hd__nand2_1_256/A sky130_fd_sc_hd__nor2_1_74/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_382 sky130_fd_sc_hd__o21ai_1_356/A1 sky130_fd_sc_hd__nor2_1_89/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_393 sky130_fd_sc_hd__a21oi_1_63/B1 sky130_fd_sc_hd__nand2_1_303/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_2_1 sky130_fd_sc_hd__a21oi_2_1/B1 sky130_fd_sc_hd__or2_0_2/X
+ sky130_fd_sc_hd__o21ai_2_6/Y sky130_fd_sc_hd__xor2_1_42/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_2
Xsky130_fd_sc_hd__a211o_1_7 vssd1 vccd1 sky130_fd_sc_hd__fa_2_275/A sky130_fd_sc_hd__dfxtp_1_70/Q
+ sky130_fd_sc_hd__nor2_1_11/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_7/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__o21ai_1_307 vssd1 vccd1 sky130_fd_sc_hd__inv_2_19/Y sky130_fd_sc_hd__nand2b_2_0/Y
+ sky130_fd_sc_hd__o21ai_1_307/B1 sky130_fd_sc_hd__xor2_1_127/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_318 vssd1 vccd1 sky130_fd_sc_hd__buf_2_2/X sky130_fd_sc_hd__nand2b_1_7/Y
+ sky130_fd_sc_hd__o21ai_1_318/B1 sky130_fd_sc_hd__xor2_1_138/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_329 vssd1 vccd1 sky130_fd_sc_hd__inv_2_26/Y sky130_fd_sc_hd__nand2b_1_7/Y
+ sky130_fd_sc_hd__nand2_1_157/Y sky130_fd_sc_hd__xor2_1_148/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__conb_1_106 sky130_fd_sc_hd__conb_1_106/LO sky130_fd_sc_hd__conb_1_106/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_117 sky130_fd_sc_hd__conb_1_117/LO sky130_fd_sc_hd__conb_1_117/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_128 sky130_fd_sc_hd__conb_1_128/LO sky130_fd_sc_hd__conb_1_128/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_139 sky130_fd_sc_hd__conb_1_139/LO sky130_fd_sc_hd__clkinv_1_3/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__xor2_1_101 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__fa_2_76/CIN
+ sky130_fd_sc_hd__xor2_1_101/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_112 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__fa_2_83/A
+ sky130_fd_sc_hd__xor2_1_112/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_123 sky130_fd_sc_hd__fa_2_97/A sky130_fd_sc_hd__fa_2_90/B
+ sky130_fd_sc_hd__xor2_1_123/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_134 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__fa_2_99/CIN
+ sky130_fd_sc_hd__xor2_1_134/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_145 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__fa_2_107/B
+ sky130_fd_sc_hd__xor2_1_145/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_156 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__fa_2_114/A
+ sky130_fd_sc_hd__xor2_1_156/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_507 sky130_fd_sc_hd__or4_1_3/C sky130_fd_sc_hd__dfxtp_1_509/CLK
+ sky130_fd_sc_hd__and2_0_393/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_167 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__fa_2_121/A
+ sky130_fd_sc_hd__xor2_1_167/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_518 sky130_fd_sc_hd__ha_2_60/A sky130_fd_sc_hd__dfxtp_1_520/CLK
+ sky130_fd_sc_hd__and2_0_346/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_178 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__fa_2_128/B
+ sky130_fd_sc_hd__xor2_1_178/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_529 wbs_dat_o[8] sky130_fd_sc_hd__dfxtp_1_532/CLK sky130_fd_sc_hd__nor2b_1_149/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_189 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__xor2_1_189/X
+ sky130_fd_sc_hd__xor2_1_189/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_105 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_52/A1 sky130_fd_sc_hd__clkbuf_1_105/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_116 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_116/X sky130_fd_sc_hd__inv_2_4/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_127 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_127/X sky130_fd_sc_hd__clkinv_2_1/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_138 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_138/X sky130_fd_sc_hd__clkinv_1_885/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o21ai_1_830 vssd1 vccd1 sky130_fd_sc_hd__inv_2_46/Y sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__o21ai_1_830/B1 sky130_fd_sc_hd__xor2_1_604/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_209 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__or2_0_52/B
+ sky130_fd_sc_hd__or2_0_53/A sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__buf_2_32/X
+ sky130_fd_sc_hd__o21ai_1_384/B1 sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_149 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_1/A1 sky130_fd_sc_hd__clkbuf_1_149/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o21ai_1_841 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_127/A sky130_fd_sc_hd__nor2_1_212/Y
+ sky130_fd_sc_hd__nand2_1_634/Y sky130_fd_sc_hd__xnor2_1_177/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_7 sky130_fd_sc_hd__buf_8_7/A sky130_fd_sc_hd__dfxtp_1_9/CLK
+ sky130_fd_sc_hd__dfxtp_1_7/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_852 vssd1 vccd1 sky130_fd_sc_hd__inv_2_48/Y sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_852/B1 sky130_fd_sc_hd__xor2_1_626/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_863 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_641/A sky130_fd_sc_hd__nor2_1_222/Y
+ sky130_fd_sc_hd__nand2_1_669/Y sky130_fd_sc_hd__xnor2_1_189/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_874 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_652/A sky130_fd_sc_hd__nor2_1_235/Y
+ sky130_fd_sc_hd__nand2_1_726/Y sky130_fd_sc_hd__xnor2_1_205/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_885 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_243/Y sky130_fd_sc_hd__nand2_1_773/Y
+ sky130_fd_sc_hd__nand2_1_772/Y sky130_fd_sc_hd__o21ai_1_885/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_896 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_679/A sky130_fd_sc_hd__nor2_1_257/Y
+ sky130_fd_sc_hd__nand2_1_805/Y sky130_fd_sc_hd__xnor2_1_293/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__inv_4_17 sky130_fd_sc_hd__inv_4_17/Y wbs_dat_i[15] vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__xor2_1_690 la_data_out[47] sky130_fd_sc_hd__xor2_1_690/X sky130_fd_sc_hd__xor2_1_690/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__and2_0_103 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_31/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_103/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_11 la_data_out[116] sky130_fd_sc_hd__conb_1_131/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_114 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_33/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_114/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_22 la_data_out[105] sky130_fd_sc_hd__conb_1_120/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_125 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_67/D sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_125/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_33 la_data_out[30] sky130_fd_sc_hd__conb_1_109/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_136 vccd1 vssd1 sky130_fd_sc_hd__and2_0_136/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_136/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_44 la_data_out[19] sky130_fd_sc_hd__conb_1_98/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_147 vccd1 vssd1 sky130_fd_sc_hd__and2_0_147/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_147/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_55 la_data_out[8] sky130_fd_sc_hd__conb_1_87/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_158 vccd1 vssd1 sky130_fd_sc_hd__and2_0_158/X sky130_fd_sc_hd__o21ai_2_0/B1
+ sky130_fd_sc_hd__and2_0_158/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_66 io_out[35] sky130_fd_sc_hd__conb_1_76/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_169 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_44/D sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_169/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_77 io_out[24] sky130_fd_sc_hd__conb_1_65/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_88 io_out[13] sky130_fd_sc_hd__conb_1_54/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_99 io_out[2] sky130_fd_sc_hd__conb_1_43/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_0 sky130_fd_sc_hd__buf_8_0/A sky130_fd_sc_hd__buf_8_0/X vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__a22o_1_2 sky130_fd_sc_hd__nand2_1_7/B sky130_fd_sc_hd__or2_0_76/B
+ sky130_fd_sc_hd__buf_4_2/A sky130_fd_sc_hd__or2_0_76/A sky130_fd_sc_hd__nand2_1_8/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_190 sky130_fd_sc_hd__o22ai_1_45/B1 sky130_fd_sc_hd__dfxtp_1_177/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_70 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__buf_2_188/X
+ sky130_fd_sc_hd__a22o_1_70/X sky130_fd_sc_hd__ha_2_39/SUM sky130_fd_sc_hd__a22o_1_71/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__inv_12_0 sky130_fd_sc_hd__inv_12_0/A sky130_fd_sc_hd__inv_12_0/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__inv_12
Xsky130_fd_sc_hd__o21ai_1_104 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_105/A2 sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__a22oi_1_162/Y sky130_fd_sc_hd__and2_0_172/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_115 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_117/A2 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_125/Y sky130_fd_sc_hd__and2_0_159/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_126 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_129/A2 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_130/Y sky130_fd_sc_hd__and2_0_145/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_137 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_137/A2 sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__a22oi_1_179/Y sky130_fd_sc_hd__and2_0_132/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_148 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_149/A2 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_140/Y sky130_fd_sc_hd__and2_0_117/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_159 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_2/B sky130_fd_sc_hd__o21ai_1_160/A1
+ sky130_fd_sc_hd__nand2_1_148/Y sky130_fd_sc_hd__and2_0_103/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__inv_8_0 sky130_fd_sc_hd__inv_8_0/A sky130_fd_sc_hd__inv_8_0/Y vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__inv_8
Xsky130_fd_sc_hd__nand2_1_508 sky130_fd_sc_hd__nor2_1_165/A sky130_fd_sc_hd__or2_0_56/X
+ sky130_fd_sc_hd__or2_0_57/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_519 sky130_fd_sc_hd__nor2_1_169/A sky130_fd_sc_hd__or2_0_58/X
+ sky130_fd_sc_hd__nand2_1_531/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_60 sky130_fd_sc_hd__nand2_1_60/Y sky130_fd_sc_hd__nand2_1_60/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_71 sky130_fd_sc_hd__nand2_1_71/Y sky130_fd_sc_hd__nand2_1_71/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_82 sky130_fd_sc_hd__nand2_1_82/Y sky130_fd_sc_hd__nand2_1_82/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_93 sky130_fd_sc_hd__nand2_1_93/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__xor2_1_255/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_304 sky130_fd_sc_hd__dfxtp_1_304/Q sky130_fd_sc_hd__clkinv_8_6/Y
+ sky130_fd_sc_hd__and2_0_280/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_315 sky130_fd_sc_hd__or2_0_88/A sky130_fd_sc_hd__dfxtp_1_319/CLK
+ sky130_fd_sc_hd__and2_0_292/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_326 sky130_fd_sc_hd__dfxtp_1_326/Q sky130_fd_sc_hd__dfxtp_1_343/CLK
+ sky130_fd_sc_hd__and2_0_317/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_337 sky130_fd_sc_hd__a22oi_1_7/B2 sky130_fd_sc_hd__dfxtp_1_339/CLK
+ sky130_fd_sc_hd__and2_0_324/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_348 sky130_fd_sc_hd__dfxtp_1_348/Q sky130_fd_sc_hd__dfxtp_1_356/CLK
+ sky130_fd_sc_hd__and2_0_309/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_359 sky130_fd_sc_hd__dfxtp_1_359/Q sky130_fd_sc_hd__dfxtp_1_29/CLK
+ sky130_fd_sc_hd__ha_2_7/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_660 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_681/A2 sky130_fd_sc_hd__nor2_1_166/A
+ sky130_fd_sc_hd__a21oi_1_109/Y sky130_fd_sc_hd__o21ai_1_660/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_671 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_671/A2 sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_671/B1 sky130_fd_sc_hd__xor2_1_454/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_682 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_771/A2 sky130_fd_sc_hd__nand2b_2_6/Y
+ sky130_fd_sc_hd__o21ai_1_682/B1 sky130_fd_sc_hd__xor2_1_461/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_209 sky130_fd_sc_hd__fa_2_205/CIN sky130_fd_sc_hd__fa_2_215/A
+ sky130_fd_sc_hd__fa_2_209/A sky130_fd_sc_hd__fa_2_209/B sky130_fd_sc_hd__fa_2_213/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o21ai_1_693 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_176/Y sky130_fd_sc_hd__nor2_1_172/A
+ sky130_fd_sc_hd__nor2_1_171/Y sky130_fd_sc_hd__o21ai_1_693/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_12 sky130_fd_sc_hd__fa_2_6/CIN sky130_fd_sc_hd__fa_2_9/B sky130_fd_sc_hd__fa_2_12/A
+ sky130_fd_sc_hd__fa_2_12/B sky130_fd_sc_hd__xor2_1_23/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_23 sky130_fd_sc_hd__fa_2_14/B sky130_fd_sc_hd__fa_2_24/B sky130_fd_sc_hd__fa_2_23/A
+ sky130_fd_sc_hd__fa_2_23/B sky130_fd_sc_hd__xor2_1_40/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_34 sky130_fd_sc_hd__fa_2_18/A sky130_fd_sc_hd__fa_2_34/SUM
+ sky130_fd_sc_hd__fa_2_34/A sky130_fd_sc_hd__fa_2_34/B sky130_fd_sc_hd__fa_2_34/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_45 sky130_fd_sc_hd__fa_2_37/B sky130_fd_sc_hd__fa_2_49/A sky130_fd_sc_hd__fa_2_45/A
+ sky130_fd_sc_hd__fa_2_45/B sky130_fd_sc_hd__fa_2_45/CIN vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_56 sky130_fd_sc_hd__fa_2_45/CIN sky130_fd_sc_hd__fa_2_58/A
+ sky130_fd_sc_hd__fa_2_56/A sky130_fd_sc_hd__fa_2_56/B sky130_fd_sc_hd__xor2_1_77/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_67 sky130_fd_sc_hd__fa_2_63/CIN sky130_fd_sc_hd__fa_2_73/A
+ sky130_fd_sc_hd__fa_2_67/A sky130_fd_sc_hd__fa_2_67/B sky130_fd_sc_hd__fa_2_71/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_78 sky130_fd_sc_hd__fa_2_71/A sky130_fd_sc_hd__fa_2_76/B sky130_fd_sc_hd__fa_2_78/A
+ sky130_fd_sc_hd__fa_2_78/B sky130_fd_sc_hd__fa_2_78/CIN vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_89 sky130_fd_sc_hd__fa_2_86/B sky130_fd_sc_hd__fa_2_92/CIN
+ sky130_fd_sc_hd__fa_2_89/A sky130_fd_sc_hd__fa_2_89/B sky130_fd_sc_hd__fa_2_89/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_204 vccd1 vssd1 la_data_out[74] sky130_fd_sc_hd__mux2_4_2/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__a222oi_1_540 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__buf_8_0/A
+ sky130_fd_sc_hd__buf_4_6/X sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__buf_4_1/X
+ sky130_fd_sc_hd__o21ai_1_852/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_551 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_419/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_451/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_748/A sky130_fd_sc_hd__dfxtp_1_387/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a21oi_1_17 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_46/Y
+ sky130_fd_sc_hd__a21oi_1_17/Y sky130_fd_sc_hd__dfxtp_1_80/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_562 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_408/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_440/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_759/A sky130_fd_sc_hd__dfxtp_1_376/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a21oi_1_28 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_57/Y
+ sky130_fd_sc_hd__a21oi_1_28/Y sky130_fd_sc_hd__dfxtp_1_69/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_573 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_396/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_428/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_770/A sky130_fd_sc_hd__dfxtp_1_364/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a21oi_1_39 sky130_fd_sc_hd__a21oi_1_39/A1 sky130_fd_sc_hd__nor2_1_45/A
+ sky130_fd_sc_hd__a21oi_1_39/Y sky130_fd_sc_hd__or2_0_10/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_584 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_407/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_439/Q sky130_fd_sc_hd__clkbuf_1_32/X
+ sky130_fd_sc_hd__clkinv_1_781/A sky130_fd_sc_hd__dfxtp_1_375/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_595 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_422/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_454/Q sky130_fd_sc_hd__nor2_4_19/B
+ sky130_fd_sc_hd__clkinv_1_792/A sky130_fd_sc_hd__dfxtp_1_390/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_13 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_24 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_35 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_140 sky130_fd_sc_hd__clkinv_4_59/Y sky130_fd_sc_hd__nor2b_1_140/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__decap_12_46 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_151 sky130_fd_sc_hd__clkinv_4_70/Y sky130_fd_sc_hd__nor2b_1_151/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__decap_12_57 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_68 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_79 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__bufbuf_8_0 sky130_fd_sc_hd__buf_6_17/X sky130_fd_sc_hd__buf_6_38/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__bufbuf_8
Xsky130_fd_sc_hd__buf_6_13 vccd1 vssd1 sky130_fd_sc_hd__buf_6_13/X sky130_fd_sc_hd__buf_6_13/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_24 vccd1 vssd1 sky130_fd_sc_hd__buf_6_24/X sky130_fd_sc_hd__buf_6_24/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_35 vccd1 vssd1 sky130_fd_sc_hd__buf_6_35/X sky130_fd_sc_hd__buf_8_97/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_46 vccd1 vssd1 sky130_fd_sc_hd__buf_6_46/X sky130_fd_sc_hd__buf_8_25/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_57 vccd1 vssd1 sky130_fd_sc_hd__buf_6_57/X sky130_fd_sc_hd__buf_6_57/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_68 vccd1 vssd1 sky130_fd_sc_hd__buf_6_68/X sky130_fd_sc_hd__buf_6_68/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_79 vccd1 vssd1 sky130_fd_sc_hd__buf_6_79/X sky130_fd_sc_hd__buf_6_79/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_15 sky130_fd_sc_hd__clkinv_4_72/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_26 sky130_fd_sc_hd__clkinv_4_61/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_37 sky130_fd_sc_hd__clkinv_4_45/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_48 sky130_fd_sc_hd__buf_2_189/A vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_59 sky130_fd_sc_hd__buf_2_192/A vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__nand2_1_305 sky130_fd_sc_hd__nand2_1_305/Y sky130_fd_sc_hd__or2_0_22/A
+ sky130_fd_sc_hd__or2_0_22/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_904 sky130_fd_sc_hd__clkinv_1_904/Y sky130_fd_sc_hd__clkinv_4_90/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_316 sky130_fd_sc_hd__nand2_1_316/Y sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__inv_6_0/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_915 sky130_fd_sc_hd__clkinv_1_917/A sky130_fd_sc_hd__buf_2_50/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_327 sky130_fd_sc_hd__nand2_1_327/Y sky130_fd_sc_hd__nor2_2_19/Y
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_926 sky130_fd_sc_hd__clkinv_1_926/Y sky130_fd_sc_hd__clkinv_1_927/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__bufinv_8_0 sky130_fd_sc_hd__bufinv_8_0/A sky130_fd_sc_hd__bufinv_8_0/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__bufinv_8
Xsky130_fd_sc_hd__nand2_1_338 sky130_fd_sc_hd__xnor2_2_1/A sky130_fd_sc_hd__nand2_1_339/Y
+ sky130_fd_sc_hd__or2_0_27/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_937 sky130_fd_sc_hd__inv_2_128/A sky130_fd_sc_hd__clkinv_1_937/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_349 sky130_fd_sc_hd__nand2_1_349/Y sky130_fd_sc_hd__or2_0_58/A
+ sky130_fd_sc_hd__or2_0_9/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_948 sky130_fd_sc_hd__clkinv_1_948/Y sky130_fd_sc_hd__inv_2_145/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_959 sky130_fd_sc_hd__clkinv_1_959/Y sky130_fd_sc_hd__clkinv_1_959/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_101 sky130_fd_sc_hd__dfxtp_1_101/Q sky130_fd_sc_hd__dfxtp_1_105/CLK
+ sky130_fd_sc_hd__and2_0_132/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1409 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_112 sky130_fd_sc_hd__dfxtp_1_112/Q sky130_fd_sc_hd__dfxtp_1_97/CLK
+ sky130_fd_sc_hd__and2_0_188/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_123 sky130_fd_sc_hd__dfxtp_1_123/Q sky130_fd_sc_hd__dfxtp_1_126/CLK
+ sky130_fd_sc_hd__and2_0_243/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_134 sky130_fd_sc_hd__dfxtp_1_134/Q sky130_fd_sc_hd__dfxtp_1_138/CLK
+ sky130_fd_sc_hd__and2_0_141/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_145 sky130_fd_sc_hd__dfxtp_1_145/Q sky130_fd_sc_hd__dfxtp_1_154/CLK
+ sky130_fd_sc_hd__and2_0_196/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_156 sky130_fd_sc_hd__dfxtp_1_156/Q sky130_fd_sc_hd__dfxtp_1_158/CLK
+ sky130_fd_sc_hd__and2_0_248/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_167 sky130_fd_sc_hd__dfxtp_1_167/Q sky130_fd_sc_hd__dfxtp_1_170/CLK
+ sky130_fd_sc_hd__and2_0_142/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_178 sky130_fd_sc_hd__dfxtp_1_178/Q sky130_fd_sc_hd__clkinv_4_2/Y
+ sky130_fd_sc_hd__and2_0_198/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_189 sky130_fd_sc_hd__dfxtp_1_189/Q sky130_fd_sc_hd__dfxtp_1_190/CLK
+ sky130_fd_sc_hd__and2_0_12/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_490 vssd1 vccd1 sky130_fd_sc_hd__inv_2_27/Y sky130_fd_sc_hd__nand2b_1_12/Y
+ sky130_fd_sc_hd__nand2_1_324/Y sky130_fd_sc_hd__xor2_1_290/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_900 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_911 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_922 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_933 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_944 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_955 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_966 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_850 sky130_fd_sc_hd__a31oi_1_0/A3 sky130_fd_sc_hd__nor2_1_274/Y
+ sky130_fd_sc_hd__nor2b_1_121/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_977 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_861 sky130_fd_sc_hd__nand2_1_861/Y sky130_fd_sc_hd__nand2_1_861/B
+ la_data_out[52] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_988 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_999 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_50 vssd1 vccd1 sky130_fd_sc_hd__inv_2_59/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_92/Y sky130_fd_sc_hd__o21ai_1_50/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_61 vssd1 vccd1 sky130_fd_sc_hd__inv_2_60/Y sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__o21ai_1_61/B1 sky130_fd_sc_hd__o21ai_1_61/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_72 vssd1 vccd1 sky130_fd_sc_hd__inv_2_57/Y sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__o21ai_1_72/B1 sky130_fd_sc_hd__o21ai_1_72/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_83 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_85/A2 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__o21ai_1_83/B1 sky130_fd_sc_hd__o21ai_1_83/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_94 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_98/A2 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__o21ai_1_94/B1 sky130_fd_sc_hd__o21ai_1_94/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__mux2_8_0 sky130_fd_sc_hd__mux2_8_0/S sky130_fd_sc_hd__mux2_8_0/A1
+ vccd1 vssd1 sky130_fd_sc_hd__buf_8_1/X la_data_out[67] vssd1 vccd1 sky130_fd_sc_hd__mux2_8
Xsky130_fd_sc_hd__a222oi_1_370 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__buf_4_7/X
+ sky130_fd_sc_hd__buf_4_0/X sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__buf_2_23/X
+ sky130_fd_sc_hd__o21ai_1_612/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_381 vccd1 vssd1 sky130_fd_sc_hd__and3_1_2/X sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__buf_8_0/X sky130_fd_sc_hd__nor2_1_174/Y sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__o21ai_1_641/B1 sky130_fd_sc_hd__nor2b_1_14/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_392 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__or2_0_61/A
+ sky130_fd_sc_hd__or2_0_61/B sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__or2_0_58/B
+ sky130_fd_sc_hd__o21ai_1_655/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a21oi_1_108 sky130_fd_sc_hd__clkinv_1_549/Y sky130_fd_sc_hd__o21ai_1_660/Y
+ sky130_fd_sc_hd__a21oi_1_108/Y sky130_fd_sc_hd__nor2_1_166/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_119 sky130_fd_sc_hd__nand2_1_593/Y sky130_fd_sc_hd__nand2_1_583/Y
+ sky130_fd_sc_hd__a21oi_1_119/Y sky130_fd_sc_hd__nor2_1_189/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_501 sky130_fd_sc_hd__buf_12_501/A sky130_fd_sc_hd__buf_12_533/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_512 sky130_fd_sc_hd__buf_12_512/A sky130_fd_sc_hd__buf_12_513/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_523 sky130_fd_sc_hd__buf_12_523/A sky130_fd_sc_hd__buf_12_523/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_534 sky130_fd_sc_hd__buf_12_534/A sky130_fd_sc_hd__buf_12_534/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_545 sky130_fd_sc_hd__buf_12_545/A sky130_fd_sc_hd__buf_12_545/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_556 sky130_fd_sc_hd__buf_12_556/A sky130_fd_sc_hd__buf_12_556/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_567 sky130_fd_sc_hd__buf_12_567/A sky130_fd_sc_hd__buf_12_567/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_578 sky130_fd_sc_hd__buf_12_578/A sky130_fd_sc_hd__buf_12_578/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_207 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_589 sky130_fd_sc_hd__buf_12_589/A sky130_fd_sc_hd__buf_12_589/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_218 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_102 sky130_fd_sc_hd__o21ai_1_70/B1 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__xnor2_1_86/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_229 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_701 sky130_fd_sc_hd__o31ai_2_0/A2 sky130_fd_sc_hd__or4_1_1/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_113 sky130_fd_sc_hd__o21ai_1_91/B1 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__xor2_1_346/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_712 sky130_fd_sc_hd__nor2b_1_91/A sky130_fd_sc_hd__fa_2_464/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_124 sky130_fd_sc_hd__nand2_1_124/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__xor2_1_384/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_723 sky130_fd_sc_hd__nor2b_1_102/A sky130_fd_sc_hd__xor2_1_680/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_135 sky130_fd_sc_hd__nand2_1_135/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_135/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_734 sky130_fd_sc_hd__nor2b_1_113/A sky130_fd_sc_hd__xnor2_1_300/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_146 sky130_fd_sc_hd__nand2_1_146/Y sky130_fd_sc_hd__xnor2_1_125/Y
+ sky130_fd_sc_hd__nor2_1_3/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_745 sky130_fd_sc_hd__fa_2_468/A sky130_fd_sc_hd__clkinv_1_745/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_308 vssd1 vccd1 sky130_fd_sc_hd__ha_2_55/SUM sky130_fd_sc_hd__nand4_1_3/D
+ la_data_out[51] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_157 sky130_fd_sc_hd__nand2_1_157/Y sky130_fd_sc_hd__nor2_2_7/Y
+ sky130_fd_sc_hd__clkbuf_1_3/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_756 sky130_fd_sc_hd__fa_2_479/A sky130_fd_sc_hd__clkinv_1_756/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_168 sky130_fd_sc_hd__nand2_1_168/Y sky130_fd_sc_hd__or2_0_0/A
+ sky130_fd_sc_hd__or2_0_0/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_767 sky130_fd_sc_hd__fa_2_490/A sky130_fd_sc_hd__clkinv_1_767/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_179 sky130_fd_sc_hd__xnor2_1_10/A sky130_fd_sc_hd__nand2_1_180/Y
+ sky130_fd_sc_hd__or2_0_1/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_778 sky130_fd_sc_hd__and2_0_329/A sky130_fd_sc_hd__clkinv_1_778/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_789 sky130_fd_sc_hd__and2_0_318/A sky130_fd_sc_hd__clkinv_1_789/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__or2_0_110 sky130_fd_sc_hd__or2_0_110/A sky130_fd_sc_hd__or2_0_110/X
+ sky130_fd_sc_hd__or2_0_110/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__decap_12_1206 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_6 sky130_fd_sc_hd__xor2_1_6/B sky130_fd_sc_hd__xor3_1_8/B
+ sky130_fd_sc_hd__xor2_1_6/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1217 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1228 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1239 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_8_4 sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__clkinv_8_4/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_12_730 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_741 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_752 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_763 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_774 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_785 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_796 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_680 sky130_fd_sc_hd__xor2_1_644/B sky130_fd_sc_hd__nand2_1_681/Y
+ sky130_fd_sc_hd__nand2_1_680/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_508 sky130_fd_sc_hd__xor2_1_548/B sky130_fd_sc_hd__fa_2_335/A
+ sky130_fd_sc_hd__xor2_1_508/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_691 sky130_fd_sc_hd__nand2_1_691/Y sky130_fd_sc_hd__or2_0_79/A
+ sky130_fd_sc_hd__or2_0_79/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_519 sky130_fd_sc_hd__xor2_1_548/B sky130_fd_sc_hd__xor2_1_519/X
+ sky130_fd_sc_hd__xor2_1_519/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1740 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1751 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_50 sky130_fd_sc_hd__inv_2_50/A sky130_fd_sc_hd__inv_2_50/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1762 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_61 sky130_fd_sc_hd__inv_2_61/A sky130_fd_sc_hd__inv_2_61/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1773 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_72 sky130_fd_sc_hd__inv_2_72/A sky130_fd_sc_hd__inv_2_72/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1784 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_83 sky130_fd_sc_hd__inv_2_83/A sky130_fd_sc_hd__inv_2_83/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1795 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_94 sky130_fd_sc_hd__inv_2_94/A sky130_fd_sc_hd__inv_2_94/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__ha_2_15 vssd1 vccd1 sky130_fd_sc_hd__ha_2_15/A sky130_fd_sc_hd__fa_2_446/B
+ sky130_fd_sc_hd__ha_2_15/SUM sky130_fd_sc_hd__ha_2_15/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_26 vssd1 vccd1 la_data_out[46] sky130_fd_sc_hd__xor2_1_690/A
+ sky130_fd_sc_hd__ha_2_26/SUM sky130_fd_sc_hd__ha_2_26/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_37 vssd1 vccd1 la_data_out[51] sky130_fd_sc_hd__ha_2_36/B sky130_fd_sc_hd__ha_2_37/SUM
+ sky130_fd_sc_hd__ha_2_37/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_48 vssd1 vccd1 sky130_fd_sc_hd__ha_2_48/A sky130_fd_sc_hd__ha_2_49/B
+ sky130_fd_sc_hd__maj3_1_1/A sky130_fd_sc_hd__ha_2_48/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_59 vssd1 vccd1 sky130_fd_sc_hd__ha_2_59/A sky130_fd_sc_hd__ha_2_58/B
+ sky130_fd_sc_hd__ha_2_59/SUM sky130_fd_sc_hd__ha_2_59/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_370 sky130_fd_sc_hd__fa_2_366/B sky130_fd_sc_hd__fa_2_371/B
+ sky130_fd_sc_hd__fa_2_370/A sky130_fd_sc_hd__fa_2_370/B sky130_fd_sc_hd__xor2_1_544/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_11 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_4_3/Y
+ sky130_fd_sc_hd__dfxtp_1_97/CLK sky130_fd_sc_hd__clkbuf_1_11/X vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_381 sky130_fd_sc_hd__fah_1_7/B sky130_fd_sc_hd__fah_1_6/CI
+ sky130_fd_sc_hd__fa_2_381/A sky130_fd_sc_hd__fa_2_381/B sky130_fd_sc_hd__fa_2_381/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_22 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_8_61/Y
+ sky130_fd_sc_hd__dfxtp_2_1/CLK sky130_fd_sc_hd__o21ai_2_2/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_392 sky130_fd_sc_hd__fa_2_390/CIN sky130_fd_sc_hd__fa_2_395/A
+ sky130_fd_sc_hd__fa_2_392/A sky130_fd_sc_hd__fa_2_392/B sky130_fd_sc_hd__xor2_1_583/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_33 sky130_fd_sc_hd__conb_1_145/LO sky130_fd_sc_hd__clkinv_2_11/A
+ sky130_fd_sc_hd__dfxtp_1_354/CLK sky130_fd_sc_hd__nand4_1_1/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_44 sky130_fd_sc_hd__conb_1_145/LO sky130_fd_sc_hd__clkinv_4_11/Y
+ sky130_fd_sc_hd__dfxtp_1_446/CLK sky130_fd_sc_hd__o31ai_2_0/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_55 sky130_fd_sc_hd__conb_1_149/LO sky130_fd_sc_hd__clkinv_4_119/A
+ sky130_fd_sc_hd__dfxtp_1_532/CLK sky130_fd_sc_hd__or2_0_113/X vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_102 sky130_fd_sc_hd__buf_8_0/X sky130_fd_sc_hd__nor2_1_102/Y
+ sky130_fd_sc_hd__buf_4_6/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_113 sky130_fd_sc_hd__nor2_1_113/B sky130_fd_sc_hd__nor2_1_113/Y
+ sky130_fd_sc_hd__nor2_1_116/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_124 sky130_fd_sc_hd__nor2_1_124/B sky130_fd_sc_hd__nor2_1_124/Y
+ sky130_fd_sc_hd__nor2_1_124/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_135 sky130_fd_sc_hd__buf_6_4/X sky130_fd_sc_hd__nor2_1_135/Y
+ sky130_fd_sc_hd__buf_6_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_11 sky130_fd_sc_hd__nor2_4_0/Y sky130_fd_sc_hd__nor2_2_0/Y
+ sky130_fd_sc_hd__dfxtp_1_335/Q sky130_fd_sc_hd__nor2_1_238/A sky130_fd_sc_hd__nand2_1_12/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_22 sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__dfxtp_1_280/Q sky130_fd_sc_hd__o211ai_1_4/Y sky130_fd_sc_hd__nand2_1_16/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_146 sky130_fd_sc_hd__buf_6_1/X sky130_fd_sc_hd__nor2_1_146/Y
+ sky130_fd_sc_hd__nor2_1_87/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_157 sky130_fd_sc_hd__buf_4_7/X sky130_fd_sc_hd__nor2_1_157/Y
+ sky130_fd_sc_hd__buf_4_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_33 sky130_fd_sc_hd__clkbuf_1_24/X sky130_fd_sc_hd__clkbuf_1_23/X
+ sky130_fd_sc_hd__dfxtp_1_95/Q sky130_fd_sc_hd__dfxtp_1_63/Q sky130_fd_sc_hd__a22oi_1_33/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_168 sky130_fd_sc_hd__nor2_1_168/B sky130_fd_sc_hd__nor2_1_168/Y
+ sky130_fd_sc_hd__nor2_1_168/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_44 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__clkbuf_1_25/X
+ sky130_fd_sc_hd__nand2_1_77/B sky130_fd_sc_hd__dfxtp_1_133/Q sky130_fd_sc_hd__a22oi_1_44/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_179 sky130_fd_sc_hd__nor2_1_179/B sky130_fd_sc_hd__nor2_1_179/Y
+ sky130_fd_sc_hd__nor2_1_179/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_55 sky130_fd_sc_hd__clkbuf_1_24/X sky130_fd_sc_hd__clkbuf_1_23/X
+ sky130_fd_sc_hd__dfxtp_1_106/Q sky130_fd_sc_hd__dfxtp_1_74/Q sky130_fd_sc_hd__a22oi_1_55/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_66 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__nor2_4_3/Y
+ sky130_fd_sc_hd__nand2_1_66/B sky130_fd_sc_hd__dfxtp_1_144/Q sky130_fd_sc_hd__a22oi_1_66/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_77 sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__dfxtp_1_117/Q sky130_fd_sc_hd__dfxtp_1_85/Q sky130_fd_sc_hd__a22oi_1_77/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_88 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__nor2_4_3/Y
+ sky130_fd_sc_hd__nand2_1_53/B sky130_fd_sc_hd__dfxtp_1_155/Q sky130_fd_sc_hd__a22oi_1_88/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_99 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_189/Q sky130_fd_sc_hd__dfxtp_1_157/Q sky130_fd_sc_hd__o21ai_1_5/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_320 sky130_fd_sc_hd__buf_12_320/A sky130_fd_sc_hd__buf_12_638/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_331 sky130_fd_sc_hd__buf_12_331/A sky130_fd_sc_hd__buf_12_588/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_342 sky130_fd_sc_hd__buf_12_84/X sky130_fd_sc_hd__buf_12_498/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_201 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__and2b_4_2/X sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__a22oi_1_201/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_353 sky130_fd_sc_hd__buf_12_353/A sky130_fd_sc_hd__buf_12_535/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_212 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__and2b_4_6/X sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__a22oi_1_212/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_364 sky130_fd_sc_hd__buf_12_364/A sky130_fd_sc_hd__buf_12_474/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_223 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__buf_2_25/A
+ sky130_fd_sc_hd__and2b_4_10/X sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__a22oi_1_223/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_375 sky130_fd_sc_hd__buf_12_375/A sky130_fd_sc_hd__buf_12_578/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_386 sky130_fd_sc_hd__buf_12_386/A sky130_fd_sc_hd__buf_12_656/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_397 sky130_fd_sc_hd__buf_12_58/X sky130_fd_sc_hd__buf_12_575/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_520 sky130_fd_sc_hd__nor2_1_164/B sky130_fd_sc_hd__nand2_1_516/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_531 sky130_fd_sc_hd__o21ai_1_681/A2 sky130_fd_sc_hd__o21ai_1_693/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_542 sky130_fd_sc_hd__clkinv_1_542/Y sky130_fd_sc_hd__nor2_1_176/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_105 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_105/B sky130_fd_sc_hd__inv_2_33/A
+ sky130_fd_sc_hd__xnor2_1_105/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_553 sky130_fd_sc_hd__nor2_1_179/B sky130_fd_sc_hd__nand2_1_559/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_116 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_118/A sky130_fd_sc_hd__and3_4_11/C
+ sky130_fd_sc_hd__xor2_1_409/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_564 sky130_fd_sc_hd__nor2_1_181/A sky130_fd_sc_hd__nand2_1_574/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_127 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_127/B sky130_fd_sc_hd__buf_2_12/A
+ sky130_fd_sc_hd__xnor2_1_127/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_575 sky130_fd_sc_hd__o21ai_1_799/A2 sky130_fd_sc_hd__nand2_1_593/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_138 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_140/B sky130_fd_sc_hd__and3_1_2/A
+ sky130_fd_sc_hd__xor2_1_475/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_586 sky130_fd_sc_hd__nand2_1_610/A sky130_fd_sc_hd__nor2_1_199/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_149 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_149/B sky130_fd_sc_hd__inv_2_57/A
+ sky130_fd_sc_hd__xnor2_1_149/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_597 sky130_fd_sc_hd__nand2_1_627/A sky130_fd_sc_hd__nor2_1_209/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_4_11 sky130_fd_sc_hd__clkinv_4_11/A sky130_fd_sc_hd__clkinv_4_11/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_22 sky130_fd_sc_hd__nand2_2_3/Y sky130_fd_sc_hd__clkinv_4_22/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_33 sky130_fd_sc_hd__clkinv_4_33/A sky130_fd_sc_hd__inv_2_157/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_44 sky130_fd_sc_hd__clkinv_4_44/A sky130_fd_sc_hd__buf_8_116/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_55 sky130_fd_sc_hd__clkinv_4_55/A sky130_fd_sc_hd__clkinv_4_55/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_66 sky130_fd_sc_hd__clkinv_4_66/A sky130_fd_sc_hd__clkinv_4_66/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_77 sky130_fd_sc_hd__clkinv_8_75/A sky130_fd_sc_hd__clkinv_4_77/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_1003 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_4_88 wbs_dat_i[11] sky130_fd_sc_hd__clkinv_4_88/Y vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_1014 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_4_99 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkinv_4_99/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_1025 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1036 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1047 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1058 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1069 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__and2b_4_14 sky130_fd_sc_hd__dfxtp_1_30/Q sky130_fd_sc_hd__o31ai_2_0/B1
+ sky130_fd_sc_hd__clkinv_1_703/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__and2b_4
Xsky130_fd_sc_hd__decap_12_560 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_571 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_582 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_593 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_305 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__xor2_1_305/X
+ sky130_fd_sc_hd__xor2_1_305/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_316 sky130_fd_sc_hd__fa_2_217/A sky130_fd_sc_hd__xor2_1_316/X
+ sky130_fd_sc_hd__xor2_1_316/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_327 sky130_fd_sc_hd__fa_2_239/A sky130_fd_sc_hd__xor2_1_327/X
+ sky130_fd_sc_hd__xor2_1_327/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_338 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__xor2_1_338/X
+ sky130_fd_sc_hd__xor2_1_338/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_349 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__fa_2_241/A
+ sky130_fd_sc_hd__xor2_1_349/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nor2b_1_90 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_90/Y
+ sky130_fd_sc_hd__nor2b_1_90/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1090 sky130_fd_sc_hd__nor2_2_0/B sky130_fd_sc_hd__nor2_4_0/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1570 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_309 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_309/X sky130_fd_sc_hd__clkbuf_1_309/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_12_1581 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1592 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_13 sky130_fd_sc_hd__buf_8_26/A sky130_fd_sc_hd__dfxtp_1_9/CLK
+ sky130_fd_sc_hd__buf_2_192/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_24 sky130_fd_sc_hd__ha_2_4/A sky130_fd_sc_hd__clkinv_8_68/Y
+ sky130_fd_sc_hd__ha_2_42/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_35 sky130_fd_sc_hd__nand2_1_79/B sky130_fd_sc_hd__dfxtp_1_45/CLK
+ sky130_fd_sc_hd__dfxtp_1_35/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_46 sky130_fd_sc_hd__nand2_1_68/B sky130_fd_sc_hd__dfxtp_1_46/CLK
+ sky130_fd_sc_hd__dfxtp_1_46/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_57 sky130_fd_sc_hd__nand2_1_56/B sky130_fd_sc_hd__dfxtp_1_57/CLK
+ sky130_fd_sc_hd__dfxtp_1_57/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_68 sky130_fd_sc_hd__dfxtp_1_68/Q sky130_fd_sc_hd__dfxtp_1_72/CLK
+ sky130_fd_sc_hd__dfxtp_1_68/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_79 sky130_fd_sc_hd__dfxtp_1_79/Q sky130_fd_sc_hd__dfxtp_1_85/CLK
+ sky130_fd_sc_hd__dfxtp_1_79/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_307 vccd1 vssd1 sky130_fd_sc_hd__and2_0_307/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_307/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_318 vccd1 vssd1 sky130_fd_sc_hd__and2_0_318/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_318/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_329 vccd1 vssd1 sky130_fd_sc_hd__and2_0_329/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_329/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__inv_2_107 sky130_fd_sc_hd__inv_2_107/A sky130_fd_sc_hd__inv_2_107/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_118 sky130_fd_sc_hd__inv_2_118/A sky130_fd_sc_hd__buf_8_27/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__or2_0_9 sky130_fd_sc_hd__or2_0_9/A sky130_fd_sc_hd__or2_0_9/X sky130_fd_sc_hd__or2_0_9/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__inv_2_129 sky130_fd_sc_hd__inv_2_129/A sky130_fd_sc_hd__buf_8_15/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_sram_1kbyte_1rw1r_32x256_8_3 sky130_fd_sc_hd__clkinv_1_965/Y sky130_fd_sc_hd__clkinv_1_965/Y
+ sky130_fd_sc_hd__buf_12_287/X sky130_fd_sc_hd__buf_12_622/X sky130_fd_sc_hd__buf_12_602/X
+ sky130_fd_sc_hd__buf_12_504/X sky130_fd_sc_hd__buf_12_605/X sky130_fd_sc_hd__buf_12_640/X
+ sky130_fd_sc_hd__buf_12_578/X sky130_fd_sc_hd__clkbuf_1_225/A sky130_fd_sc_hd__buf_12_559/X
+ sky130_fd_sc_hd__buf_12_580/X sky130_fd_sc_hd__buf_12_540/X vccd1 sky130_fd_sc_hd__clkinv_2_46/Y
+ sky130_fd_sc_hd__a22o_1_37/B2 sky130_fd_sc_hd__a22o_1_36/B2 sky130_fd_sc_hd__clkbuf_1_169/A
+ sky130_fd_sc_hd__clkbuf_1_183/A sky130_fd_sc_hd__clkbuf_1_170/A sky130_fd_sc_hd__clkbuf_1_171/A
+ sky130_fd_sc_hd__clkbuf_1_309/A sky130_fd_sc_hd__clkbuf_1_173/A sky130_fd_sc_hd__clkbuf_1_174/A
+ sky130_fd_sc_hd__clkbuf_1_176/A sky130_fd_sc_hd__clkbuf_1_177/A sky130_fd_sc_hd__clkbuf_1_175/A
+ sky130_fd_sc_hd__clkbuf_1_178/A sky130_fd_sc_hd__clkbuf_1_179/A sky130_fd_sc_hd__clkbuf_1_181/A
+ sky130_fd_sc_hd__clkbuf_1_182/A sky130_fd_sc_hd__buf_12_526/X sky130_fd_sc_hd__a22o_1_52/B2
+ sky130_fd_sc_hd__a22o_1_51/B2 sky130_fd_sc_hd__a22o_1_50/B2 sky130_fd_sc_hd__a22o_1_49/B2
+ sky130_fd_sc_hd__a22o_1_48/B2 sky130_fd_sc_hd__a22o_1_47/B2 sky130_fd_sc_hd__a22o_1_46/B2
+ sky130_fd_sc_hd__a22o_1_45/B2 sky130_fd_sc_hd__a22o_1_44/B2 sky130_fd_sc_hd__a22o_1_43/B2
+ sky130_fd_sc_hd__a22o_1_42/B2 sky130_fd_sc_hd__a22o_1_41/B2 sky130_fd_sc_hd__a22o_1_40/B2
+ sky130_fd_sc_hd__a22o_1_39/B2 sky130_fd_sc_hd__a22o_1_38/B2 sky130_fd_sc_hd__a22o_1_53/B2
+ sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[10] sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[11]
+ sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[12] sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[13]
+ sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[14] sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[15]
+ sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[16] sky130_fd_sc_hd__buf_12_555/X sky130_fd_sc_hd__buf_12_270/X
+ sky130_fd_sc_hd__buf_12_62/X sky130_fd_sc_hd__buf_12_82/X sky130_fd_sc_hd__buf_12_119/X
+ sky130_fd_sc_hd__clkinv_8_43/Y sky130_fd_sc_hd__clkinv_1_983/Y sky130_fd_sc_hd__clkbuf_1_324/X
+ sky130_fd_sc_hd__clkinv_1_979/Y sky130_fd_sc_hd__clkbuf_1_114/X sky130_fd_sc_hd__clkbuf_1_113/X
+ sky130_fd_sc_hd__buf_2_131/X sky130_fd_sc_hd__clkinv_1_973/Y sky130_fd_sc_hd__buf_2_130/X
+ sky130_fd_sc_hd__clkbuf_1_112/X sky130_fd_sc_hd__buf_2_129/X sky130_fd_sc_hd__inv_2_156/Y
+ sky130_fd_sc_hd__clkbuf_1_115/X sky130_fd_sc_hd__clkinv_1_988/Y sky130_fd_sc_hd__inv_2_155/Y
+ sky130_fd_sc_hd__clkinv_1_986/Y sky130_fd_sc_hd__clkinv_1_984/Y sky130_fd_sc_hd__clkinv_1_1015/Y
+ sky130_fd_sc_hd__clkbuf_1_131/X sky130_fd_sc_hd__clkinv_1_1013/Y sky130_fd_sc_hd__clkinv_1_1011/Y
+ sky130_fd_sc_hd__clkinv_1_1009/Y sky130_fd_sc_hd__clkinv_1_1007/Y sky130_fd_sc_hd__clkinv_1_1005/Y
+ sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[0] sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[1]
+ sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[2] sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[3]
+ sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[4] sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[5]
+ sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[6] sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[7]
+ sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[8] sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[9]
+ sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[25] sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[26]
+ sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[27] sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[28]
+ sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[29] sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[30]
+ sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[31] sky130_fd_sc_hd__inv_2_157/Y sky130_fd_sc_hd__clkinv_1_1003/Y
+ sky130_fd_sc_hd__clkbuf_1_124/X sky130_fd_sc_hd__clkinv_2_36/Y sky130_fd_sc_hd__clkinv_1_1000/Y
+ sky130_fd_sc_hd__clkinv_1_998/Y sky130_fd_sc_hd__clkinv_1_996/Y sky130_fd_sc_hd__clkinv_1_994/Y
+ sky130_fd_sc_hd__clkbuf_1_117/X sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[17] sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[18]
+ sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[19] sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[20]
+ sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[21] sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[22]
+ sky130_fd_sc_hd__buf_12_650/X sky130_fd_sc_hd__buf_12_544/X sky130_fd_sc_hd__buf_12_534/X
+ sky130_fd_sc_hd__buf_12_547/X sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[23] sky130_sram_1kbyte_1rw1r_32x256_8_3/dout0[24]
+ sky130_sram_1kbyte_1rw1r_32x256_8_3/sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/gnd_uq26
+ vssd1 sky130_sram_1kbyte_1rw1r_32x256_8
Xsky130_fd_sc_hd__buf_12_150 sky130_fd_sc_hd__buf_8_38/X sky130_fd_sc_hd__buf_12_374/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_161 sky130_fd_sc_hd__buf_8_49/X sky130_fd_sc_hd__buf_12_161/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_172 sky130_fd_sc_hd__buf_8_121/X sky130_fd_sc_hd__buf_12_447/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_183 sky130_fd_sc_hd__buf_12_57/X sky130_fd_sc_hd__buf_12_383/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_194 sky130_fd_sc_hd__buf_8_164/X sky130_fd_sc_hd__buf_12_458/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_350 sky130_fd_sc_hd__nand2_1_217/A sky130_fd_sc_hd__nor2_1_65/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_361 sky130_fd_sc_hd__nand2_1_234/A sky130_fd_sc_hd__nor2_1_71/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_372 sky130_fd_sc_hd__nand2_1_257/A sky130_fd_sc_hd__nor2_1_81/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_383 sky130_fd_sc_hd__nand2_1_273/A sky130_fd_sc_hd__nor2_1_90/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_394 sky130_fd_sc_hd__a21oi_1_64/B1 sky130_fd_sc_hd__nand2_1_300/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_2_2 sky130_fd_sc_hd__a21oi_2_2/B1 sky130_fd_sc_hd__or2_0_3/X
+ sky130_fd_sc_hd__xnor2_1_19/B sky130_fd_sc_hd__xor2_1_63/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_2
Xsky130_fd_sc_hd__a211o_1_8 vssd1 vccd1 sky130_fd_sc_hd__fa_2_273/A sky130_fd_sc_hd__dfxtp_1_71/Q
+ sky130_fd_sc_hd__nor2_1_12/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_8/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__o21ai_1_308 vssd1 vccd1 sky130_fd_sc_hd__inv_2_24/Y sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__o21ai_1_308/B1 sky130_fd_sc_hd__xor2_1_128/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_319 vssd1 vccd1 sky130_fd_sc_hd__inv_2_16/Y sky130_fd_sc_hd__nand2b_1_1/Y
+ sky130_fd_sc_hd__o21ai_1_319/B1 sky130_fd_sc_hd__xor2_1_139/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__conb_1_107 sky130_fd_sc_hd__conb_1_107/LO sky130_fd_sc_hd__conb_1_107/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_118 sky130_fd_sc_hd__conb_1_118/LO sky130_fd_sc_hd__conb_1_118/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_129 sky130_fd_sc_hd__conb_1_129/LO sky130_fd_sc_hd__conb_1_129/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_390 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_102 sky130_fd_sc_hd__fa_2_97/A sky130_fd_sc_hd__fa_2_78/B
+ sky130_fd_sc_hd__xor2_1_102/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_113 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__fa_2_85/CIN
+ sky130_fd_sc_hd__xor2_1_113/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_124 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__fa_2_87/A
+ sky130_fd_sc_hd__xor2_1_124/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_135 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__fa_2_99/B
+ sky130_fd_sc_hd__xor2_1_135/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_146 sky130_fd_sc_hd__xor2_1_146/B sky130_fd_sc_hd__xor2_1_146/X
+ sky130_fd_sc_hd__xor2_1_146/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_157 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__fah_1_1/CI
+ sky130_fd_sc_hd__xor2_1_157/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_508 sky130_fd_sc_hd__or4_1_3/B sky130_fd_sc_hd__dfxtp_1_509/CLK
+ sky130_fd_sc_hd__and2_0_394/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_168 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__fa_2_120/B
+ sky130_fd_sc_hd__xor2_1_168/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_519 sky130_fd_sc_hd__ha_2_59/A sky130_fd_sc_hd__dfxtp_1_520/CLK
+ sky130_fd_sc_hd__and2_0_345/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_179 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__fa_2_127/B
+ sky130_fd_sc_hd__xor2_1_179/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_106 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_50/A1 sky130_fd_sc_hd__clkbuf_1_106/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_117 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_117/X sky130_fd_sc_hd__buf_2_132/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_128 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_128/X sky130_fd_sc_hd__inv_4_1/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o21ai_1_820 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_3/Y sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_820/B1 sky130_fd_sc_hd__xor2_1_593/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_1_139 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_139/X sky130_fd_sc_hd__clkbuf_4_7/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o21ai_1_831 vssd1 vccd1 sky130_fd_sc_hd__nand2_2_13/Y sky130_fd_sc_hd__nand2b_2_6/Y
+ sky130_fd_sc_hd__a22oi_1_219/Y sky130_fd_sc_hd__xor2_1_605/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_842 vssd1 vccd1 sky130_fd_sc_hd__buf_2_13/X sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__o21ai_1_842/B1 sky130_fd_sc_hd__xor2_1_614/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_8 sky130_fd_sc_hd__dfxtp_1_8/Q sky130_fd_sc_hd__dfxtp_1_8/CLK
+ la_data_out[62] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_853 vssd1 vccd1 sky130_fd_sc_hd__inv_2_46/Y sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_853/B1 sky130_fd_sc_hd__xor2_1_627/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_864 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_642/A sky130_fd_sc_hd__nor2_1_223/Y
+ sky130_fd_sc_hd__nand2_1_673/Y sky130_fd_sc_hd__xnor2_1_190/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_875 vssd1 vccd1 sky130_fd_sc_hd__a21oi_1_153/Y sky130_fd_sc_hd__nand2_1_727/Y
+ sky130_fd_sc_hd__a21oi_1_151/Y sky130_fd_sc_hd__o21ai_1_875/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_886 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_246/Y sky130_fd_sc_hd__nand2_1_776/Y
+ sky130_fd_sc_hd__nand2_1_775/Y sky130_fd_sc_hd__o21ai_1_886/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_897 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_680/A sky130_fd_sc_hd__nor2_1_258/Y
+ sky130_fd_sc_hd__nand2_1_809/Y sky130_fd_sc_hd__xnor2_1_294/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__inv_4_18 sky130_fd_sc_hd__inv_4_18/Y wbs_dat_i[14] vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__xor2_1_680 sky130_fd_sc_hd__xor2_1_680/B sky130_fd_sc_hd__xor2_1_680/X
+ sky130_fd_sc_hd__xor2_1_680/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_691 la_data_out[56] sky130_fd_sc_hd__xor2_1_691/X sky130_fd_sc_hd__xor2_1_691/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__and2_0_104 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_63/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_104/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_12 la_data_out[115] sky130_fd_sc_hd__conb_1_130/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_115 vccd1 vssd1 sky130_fd_sc_hd__and2_0_115/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_115/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_23 la_data_out[104] sky130_fd_sc_hd__conb_1_119/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_126 vccd1 vssd1 sky130_fd_sc_hd__and2_0_126/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_126/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_34 la_data_out[29] sky130_fd_sc_hd__conb_1_108/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_137 vccd1 vssd1 sky130_fd_sc_hd__and2_0_137/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_137/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_45 la_data_out[18] sky130_fd_sc_hd__conb_1_97/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_148 vccd1 vssd1 sky130_fd_sc_hd__and2_0_148/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_148/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_56 la_data_out[7] sky130_fd_sc_hd__conb_1_86/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_159 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_42/D sky130_fd_sc_hd__o21ai_2_0/B1
+ sky130_fd_sc_hd__and2_0_159/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_67 io_out[34] sky130_fd_sc_hd__conb_1_75/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_78 io_out[23] sky130_fd_sc_hd__conb_1_64/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_89 io_out[12] sky130_fd_sc_hd__conb_1_53/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_1 sky130_fd_sc_hd__buf_8_1/A sky130_fd_sc_hd__buf_8_1/X vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__a22o_1_3 sky130_fd_sc_hd__nand2_1_7/B sky130_fd_sc_hd__mux2_2_8/X
+ sky130_fd_sc_hd__buf_4_3/A sky130_fd_sc_hd__mux2_2_39/X sky130_fd_sc_hd__nand2_1_8/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_180 sky130_fd_sc_hd__o22ai_1_22/B1 sky130_fd_sc_hd__dfxtp_1_117/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_191 sky130_fd_sc_hd__nor2_1_22/A sky130_fd_sc_hd__dfxtp_1_145/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_60 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__and2_0_354/A
+ sky130_fd_sc_hd__a22o_1_60/X sky130_fd_sc_hd__ha_2_31/SUM sky130_fd_sc_hd__a22o_1_71/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_71 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__and2_0_352/A
+ sky130_fd_sc_hd__a22o_1_71/X sky130_fd_sc_hd__a22o_1_71/B2 sky130_fd_sc_hd__a22o_1_71/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__inv_12_1 sky130_fd_sc_hd__inv_4_11/Y sky130_fd_sc_hd__inv_12_1/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__inv_12
Xsky130_fd_sc_hd__o21ai_1_105 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_105/A2 sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__a22oi_1_163/Y sky130_fd_sc_hd__and2_0_171/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_116 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_117/A2 sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__a22oi_1_168/Y sky130_fd_sc_hd__and2_0_158/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_127 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_129/A2 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_131/Y sky130_fd_sc_hd__and2_0_144/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_138 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_141/A2 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_136/Y sky130_fd_sc_hd__and2_0_130/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_149 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_149/A2 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_141/Y sky130_fd_sc_hd__and2_0_116/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__inv_8_1 sky130_fd_sc_hd__inv_8_1/A sky130_fd_sc_hd__inv_8_1/Y vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__inv_8
Xsky130_fd_sc_hd__nand2_1_509 sky130_fd_sc_hd__xnor2_1_131/A sky130_fd_sc_hd__nand2_1_510/Y
+ sky130_fd_sc_hd__or2_0_54/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_50 sky130_fd_sc_hd__o21ai_2_1/A2 sky130_fd_sc_hd__nor2_1_0/Y
+ sky130_fd_sc_hd__nand2_1_8/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_61 sky130_fd_sc_hd__nand2_1_61/Y sky130_fd_sc_hd__nand2_1_61/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_72 sky130_fd_sc_hd__nand2_1_72/Y sky130_fd_sc_hd__nand2_1_72/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_83 sky130_fd_sc_hd__nand2_1_83/Y sky130_fd_sc_hd__nand2_1_83/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_94 sky130_fd_sc_hd__nand2_1_94/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__xnor2_1_78/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_305 sky130_fd_sc_hd__dfxtp_1_305/Q sky130_fd_sc_hd__clkinv_8_6/Y
+ sky130_fd_sc_hd__and2_0_281/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_316 sky130_fd_sc_hd__or2_0_89/A sky130_fd_sc_hd__dfxtp_1_319/CLK
+ sky130_fd_sc_hd__and2_0_293/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_327 sky130_fd_sc_hd__dfxtp_1_327/Q sky130_fd_sc_hd__dfxtp_1_339/CLK
+ sky130_fd_sc_hd__and2_0_321/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_338 sky130_fd_sc_hd__a22oi_1_5/B2 sky130_fd_sc_hd__dfxtp_1_339/CLK
+ sky130_fd_sc_hd__and2_0_332/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_349 sky130_fd_sc_hd__dfxtp_1_349/Q sky130_fd_sc_hd__dfxtp_1_356/CLK
+ sky130_fd_sc_hd__and2_0_308/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_650 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_10/X sky130_fd_sc_hd__or2_0_55/X
+ sky130_fd_sc_hd__o21a_1_4/X sky130_fd_sc_hd__xnor2_1_131/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_661 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_751/A2 sky130_fd_sc_hd__nand2b_2_6/Y
+ sky130_fd_sc_hd__o21ai_1_661/B1 sky130_fd_sc_hd__xor2_1_444/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_672 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_10/X sky130_fd_sc_hd__nand2_1_518/Y
+ sky130_fd_sc_hd__a21oi_1_110/Y sky130_fd_sc_hd__xnor2_1_135/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_683 vssd1 vccd1 sky130_fd_sc_hd__buf_2_12/X sky130_fd_sc_hd__nand2b_1_20/Y
+ sky130_fd_sc_hd__o21ai_1_683/B1 sky130_fd_sc_hd__xor2_1_462/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_694 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_780/A2 sky130_fd_sc_hd__nand2b_2_6/Y
+ sky130_fd_sc_hd__o21ai_1_694/B1 sky130_fd_sc_hd__xor2_1_472/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_13 sky130_fd_sc_hd__fa_2_4/A sky130_fd_sc_hd__fa_2_14/A sky130_fd_sc_hd__fa_2_13/A
+ sky130_fd_sc_hd__fa_2_13/B sky130_fd_sc_hd__xor2_1_29/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_24 sky130_fd_sc_hd__fa_2_15/A sky130_fd_sc_hd__fa_2_25/B sky130_fd_sc_hd__fa_2_24/A
+ sky130_fd_sc_hd__fa_2_24/B sky130_fd_sc_hd__fa_2_24/CIN vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_35 sky130_fd_sc_hd__or2_0_1/A sky130_fd_sc_hd__nor2_1_52/B
+ sky130_fd_sc_hd__fa_2_35/A sky130_fd_sc_hd__fa_2_35/B sky130_fd_sc_hd__fa_2_35/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_46 sky130_fd_sc_hd__fa_2_41/A sky130_fd_sc_hd__fa_2_47/B sky130_fd_sc_hd__fa_2_46/A
+ sky130_fd_sc_hd__fa_2_46/B sky130_fd_sc_hd__fa_2_46/CIN vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_57 sky130_fd_sc_hd__fa_2_44/B sky130_fd_sc_hd__fa_2_57/SUM
+ sky130_fd_sc_hd__fa_2_57/A sky130_fd_sc_hd__fa_2_57/B sky130_fd_sc_hd__xor2_1_75/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_68 sky130_fd_sc_hd__fa_2_63/B sky130_fd_sc_hd__fa_2_70/B sky130_fd_sc_hd__fa_2_68/A
+ sky130_fd_sc_hd__fa_2_68/B sky130_fd_sc_hd__xor2_1_92/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_79 sky130_fd_sc_hd__fa_2_67/B sky130_fd_sc_hd__fa_2_79/SUM
+ sky130_fd_sc_hd__fa_2_79/A sky130_fd_sc_hd__fa_2_79/B sky130_fd_sc_hd__fa_2_79/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_205 vccd1 vssd1 la_data_out[66] sky130_fd_sc_hd__or2_0_84/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__a222oi_1_530 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__buf_6_2/A
+ sky130_fd_sc_hd__buf_4_1/X sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__buf_4_0/A
+ sky130_fd_sc_hd__o21ai_1_837/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_541 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__buf_8_0/A sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__buf_4_6/X
+ sky130_fd_sc_hd__o21ai_1_853/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_552 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_418/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_450/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_749/A sky130_fd_sc_hd__dfxtp_1_386/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a21oi_1_18 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_47/Y
+ sky130_fd_sc_hd__a21oi_1_18/Y sky130_fd_sc_hd__dfxtp_1_79/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_563 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_407/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_439/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_760/A sky130_fd_sc_hd__dfxtp_1_375/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a21oi_1_29 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_58/Y
+ sky130_fd_sc_hd__a21oi_1_29/Y sky130_fd_sc_hd__dfxtp_1_68/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_574 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_397/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_429/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_771/A sky130_fd_sc_hd__dfxtp_1_365/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_585 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_402/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_434/Q sky130_fd_sc_hd__clkbuf_1_32/X
+ sky130_fd_sc_hd__clkinv_1_782/A sky130_fd_sc_hd__dfxtp_1_370/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_596 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_423/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_455/Q sky130_fd_sc_hd__nor2_4_19/B
+ sky130_fd_sc_hd__clkinv_1_793/A sky130_fd_sc_hd__dfxtp_1_391/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_14 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_25 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_130 sky130_fd_sc_hd__clkinv_4_49/Y sky130_fd_sc_hd__nor2b_1_130/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__decap_12_36 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_141 sky130_fd_sc_hd__clkinv_4_60/Y sky130_fd_sc_hd__nor2b_1_141/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__decap_12_47 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_152 sky130_fd_sc_hd__clkinv_4_71/Y sky130_fd_sc_hd__nor2b_1_152/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__decap_12_58 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_69 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__fah_1_10 sky130_fd_sc_hd__nor2_2_30/A sky130_fd_sc_hd__fah_1_10/B
+ sky130_fd_sc_hd__fah_1_10/A sky130_fd_sc_hd__nor2_1_200/B sky130_fd_sc_hd__fah_1_10/CI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__fah_1
Xsky130_fd_sc_hd__bufbuf_8_1 sky130_fd_sc_hd__buf_2_162/X sky130_fd_sc_hd__buf_12_81/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__bufbuf_8
Xsky130_fd_sc_hd__buf_6_14 vccd1 vssd1 sky130_fd_sc_hd__buf_6_14/X sky130_fd_sc_hd__buf_6_14/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_25 vccd1 vssd1 sky130_fd_sc_hd__buf_6_25/X sky130_fd_sc_hd__buf_6_25/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_36 vccd1 vssd1 sky130_fd_sc_hd__buf_6_36/X sky130_fd_sc_hd__buf_8_84/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_47 vccd1 vssd1 sky130_fd_sc_hd__buf_6_47/X sky130_fd_sc_hd__buf_8_26/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_58 vccd1 vssd1 sky130_fd_sc_hd__buf_6_58/X sky130_fd_sc_hd__buf_8_88/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_69 vccd1 vssd1 sky130_fd_sc_hd__buf_6_69/X sky130_fd_sc_hd__buf_8_11/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_16 sky130_fd_sc_hd__clkinv_4_60/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_27 sky130_fd_sc_hd__clkinv_4_61/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_38 sky130_fd_sc_hd__clkinv_4_48/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_49 sky130_fd_sc_hd__buf_2_189/A vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__nand2_1_306 sky130_fd_sc_hd__xnor2_1_58/A sky130_fd_sc_hd__nand2_1_307/Y
+ sky130_fd_sc_hd__nand2_1_306/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_905 sky130_fd_sc_hd__clkinv_1_905/Y sky130_fd_sc_hd__inv_4_21/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_317 sky130_fd_sc_hd__xor2_1_209/A sky130_fd_sc_hd__o21a_1_1/B1
+ sky130_fd_sc_hd__nand2_1_317/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_916 sky130_fd_sc_hd__clkinv_1_916/Y sky130_fd_sc_hd__inv_2_108/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_328 sky130_fd_sc_hd__nand2_1_328/Y sky130_fd_sc_hd__nor2_2_20/Y
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_927 sky130_fd_sc_hd__inv_6_1/A sky130_fd_sc_hd__clkinv_1_927/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__bufinv_8_1 sky130_fd_sc_hd__bufinv_8_1/A sky130_fd_sc_hd__bufinv_8_1/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__bufinv_8
Xsky130_fd_sc_hd__nand2_1_339 sky130_fd_sc_hd__nand2_1_339/Y sky130_fd_sc_hd__or2_0_27/A
+ sky130_fd_sc_hd__or2_0_27/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_938 sky130_fd_sc_hd__inv_2_130/A sky130_fd_sc_hd__buf_8_15/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_949 sky130_fd_sc_hd__clkbuf_1_49/A sky130_fd_sc_hd__clkinv_4_20/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_102 sky130_fd_sc_hd__dfxtp_1_102/Q sky130_fd_sc_hd__dfxtp_1_105/CLK
+ sky130_fd_sc_hd__and2_0_137/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_113 sky130_fd_sc_hd__dfxtp_1_113/Q sky130_fd_sc_hd__dfxtp_1_122/CLK
+ sky130_fd_sc_hd__and2_0_192/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_124 sky130_fd_sc_hd__dfxtp_1_124/Q sky130_fd_sc_hd__dfxtp_1_126/CLK
+ sky130_fd_sc_hd__and2_0_247/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_135 sky130_fd_sc_hd__dfxtp_1_135/Q sky130_fd_sc_hd__dfxtp_1_138/CLK
+ sky130_fd_sc_hd__and2_0_148/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_146 sky130_fd_sc_hd__dfxtp_1_146/Q sky130_fd_sc_hd__dfxtp_1_146/CLK
+ sky130_fd_sc_hd__and2_0_201/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_157 sky130_fd_sc_hd__dfxtp_1_157/Q sky130_fd_sc_hd__dfxtp_1_158/CLK
+ sky130_fd_sc_hd__and2_0_249/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_168 sky130_fd_sc_hd__dfxtp_1_168/Q sky130_fd_sc_hd__dfxtp_1_170/CLK
+ sky130_fd_sc_hd__and2_0_146/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_179 sky130_fd_sc_hd__dfxtp_1_179/Q sky130_fd_sc_hd__clkinv_4_2/Y
+ sky130_fd_sc_hd__and2_0_202/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_480 vssd1 vccd1 sky130_fd_sc_hd__inv_2_28/Y sky130_fd_sc_hd__nand2b_1_13/Y
+ sky130_fd_sc_hd__o21ai_1_480/B1 sky130_fd_sc_hd__xor2_1_281/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_491 vssd1 vccd1 sky130_fd_sc_hd__inv_2_32/Y sky130_fd_sc_hd__nand2b_1_9/Y
+ sky130_fd_sc_hd__o21ai_1_491/B1 sky130_fd_sc_hd__xor2_1_292/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_901 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_912 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_923 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_934 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_945 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_956 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_840 sky130_fd_sc_hd__xor2_1_688/A sky130_fd_sc_hd__nand2_1_841/Y
+ sky130_fd_sc_hd__nand2_1_840/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_967 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_851 sky130_fd_sc_hd__o31ai_1_1/B1 sky130_fd_sc_hd__o31ai_1_1/A1
+ sky130_fd_sc_hd__nor2_1_273/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_978 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_862 sky130_fd_sc_hd__nor4_1_1/D wbs_stb_i wbs_cyc_i vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_989 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_40 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_41/A2 sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__o21ai_1_40/B1 sky130_fd_sc_hd__and2_0_12/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_51 vssd1 vccd1 sky130_fd_sc_hd__inv_2_59/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_93/Y sky130_fd_sc_hd__o21ai_1_51/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_62 vssd1 vccd1 sky130_fd_sc_hd__inv_2_55/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_98/Y sky130_fd_sc_hd__o21ai_1_62/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_73 vssd1 vccd1 sky130_fd_sc_hd__inv_2_57/Y sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_73/B1 sky130_fd_sc_hd__o21ai_1_73/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_84 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_85/A2 sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__o21ai_1_84/B1 sky130_fd_sc_hd__o21ai_1_84/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_95 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_98/A2 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__o21ai_1_95/B1 sky130_fd_sc_hd__o21ai_1_95/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nand2_4_0 sky130_fd_sc_hd__buf_2_25/A sky130_fd_sc_hd__nand2_4_0/A
+ sky130_fd_sc_hd__nand2_4_0/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_4
Xsky130_fd_sc_hd__mux2_8_1 sky130_fd_sc_hd__mux2_8_1/S sky130_fd_sc_hd__mux2_8_1/A1
+ vccd1 vssd1 sky130_fd_sc_hd__buf_4_10/X la_data_out[71] vssd1 vccd1 sky130_fd_sc_hd__mux2_8
Xsky130_fd_sc_hd__a222oi_1_360 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__buf_4_0/X
+ sky130_fd_sc_hd__buf_2_23/X sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__buf_2_31/X
+ sky130_fd_sc_hd__o21ai_1_594/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_371 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__buf_8_0/X sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__o21ai_1_613/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_382 vccd1 vssd1 sky130_fd_sc_hd__and3_4_25/X sky130_fd_sc_hd__buf_2_21/X
+ sky130_fd_sc_hd__nor2_1_87/A sky130_fd_sc_hd__nor2_1_186/Y sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__o21ai_1_643/B1 sky130_fd_sc_hd__nor2b_1_17/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_393 vccd1 vssd1 sky130_fd_sc_hd__and3_4_21/X sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__or2_0_60/B sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__or2_0_60/A
+ sky130_fd_sc_hd__o21ai_1_656/B1 sky130_fd_sc_hd__and2b_4_12/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a21oi_1_109 sky130_fd_sc_hd__clkinv_1_523/Y sky130_fd_sc_hd__nor2_1_164/A
+ sky130_fd_sc_hd__a21oi_1_109/Y sky130_fd_sc_hd__or2_0_57/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_502 sky130_fd_sc_hd__buf_12_502/A sky130_fd_sc_hd__buf_12_502/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_513 sky130_fd_sc_hd__buf_12_513/A sky130_fd_sc_hd__buf_12_546/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_524 sky130_fd_sc_hd__buf_12_524/A sky130_fd_sc_hd__buf_12_524/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_535 sky130_fd_sc_hd__buf_12_535/A sky130_fd_sc_hd__buf_12_535/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_546 sky130_fd_sc_hd__buf_12_546/A sky130_fd_sc_hd__buf_12_546/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_557 sky130_fd_sc_hd__buf_12_557/A sky130_fd_sc_hd__buf_12_557/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_568 sky130_fd_sc_hd__buf_12_568/A sky130_fd_sc_hd__buf_12_568/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_579 sky130_fd_sc_hd__buf_12_579/A sky130_fd_sc_hd__buf_12_579/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_208 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_219 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_103 sky130_fd_sc_hd__o21ai_1_71/B1 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__xnor2_1_86/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_702 sky130_fd_sc_hd__nand4_1_0/B sky130_fd_sc_hd__ha_2_8/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_114 sky130_fd_sc_hd__o21ai_1_94/B1 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__xor2_1_359/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_713 sky130_fd_sc_hd__nor2b_1_92/A sky130_fd_sc_hd__fa_2_466/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_125 sky130_fd_sc_hd__nand2_1_125/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__xor2_1_384/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_724 sky130_fd_sc_hd__nor2b_1_103/A sky130_fd_sc_hd__xnor2_1_295/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_136 sky130_fd_sc_hd__nand2_1_136/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__xor2_1_411/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_735 sky130_fd_sc_hd__nor2b_1_114/A sky130_fd_sc_hd__xor2_1_686/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_147 sky130_fd_sc_hd__nor2_1_36/A sky130_fd_sc_hd__nor2_1_40/A
+ sky130_fd_sc_hd__nand2_1_147/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_746 sky130_fd_sc_hd__fa_2_469/A sky130_fd_sc_hd__clkinv_1_746/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_309 vssd1 vccd1 la_data_out[48] sky130_fd_sc_hd__nand4_1_3/C
+ sky130_fd_sc_hd__xnor2_1_309/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_158 sky130_fd_sc_hd__nand2_1_158/Y sky130_fd_sc_hd__nor2_2_8/Y
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_757 sky130_fd_sc_hd__fa_2_480/A sky130_fd_sc_hd__clkinv_1_757/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_169 sky130_fd_sc_hd__nand2_1_169/Y sky130_fd_sc_hd__nor2_1_47/Y
+ sky130_fd_sc_hd__nand2_1_203/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_768 sky130_fd_sc_hd__fa_2_491/A sky130_fd_sc_hd__clkinv_1_768/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_779 sky130_fd_sc_hd__and2_0_328/A sky130_fd_sc_hd__clkinv_1_779/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__or2_0_100 sky130_fd_sc_hd__or2_0_100/A sky130_fd_sc_hd__or2_0_100/X
+ sky130_fd_sc_hd__or2_0_100/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_111 sky130_fd_sc_hd__or2_0_111/A sky130_fd_sc_hd__or2_0_111/X
+ sky130_fd_sc_hd__or2_0_111/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__decap_12_1207 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_7 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__xor3_1_7/A
+ sky130_fd_sc_hd__xor2_1_7/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1218 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1229 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_8_5 sky130_fd_sc_hd__clkinv_8_5/Y sky130_fd_sc_hd__clkinv_8_5/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_12_720 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_731 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_742 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_753 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_764 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_775 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_786 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_670 sky130_fd_sc_hd__xnor2_1_190/A sky130_fd_sc_hd__nand2_1_671/Y
+ sky130_fd_sc_hd__or2_0_75/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_797 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_681 sky130_fd_sc_hd__nand2_1_681/Y sky130_fd_sc_hd__mux2_2_18/X
+ sky130_fd_sc_hd__mux2_2_37/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_509 sky130_fd_sc_hd__xor2_1_509/B sky130_fd_sc_hd__inv_2_56/A
+ sky130_fd_sc_hd__xor2_1_509/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_692 sky130_fd_sc_hd__xor2_1_647/B sky130_fd_sc_hd__nand2_1_693/Y
+ sky130_fd_sc_hd__nand2_1_692/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_1730 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1741 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_40 sky130_fd_sc_hd__inv_2_40/A sky130_fd_sc_hd__inv_2_40/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1752 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_51 sky130_fd_sc_hd__inv_2_51/A sky130_fd_sc_hd__inv_2_51/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1763 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_62 sky130_fd_sc_hd__buf_6_3/X sky130_fd_sc_hd__inv_2_62/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1774 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_73 sky130_fd_sc_hd__inv_2_73/A sky130_fd_sc_hd__inv_2_73/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1785 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_84 sky130_fd_sc_hd__inv_2_84/A sky130_fd_sc_hd__inv_2_84/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1796 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_95 sky130_fd_sc_hd__inv_2_95/A sky130_fd_sc_hd__inv_2_95/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__ha_2_16 vssd1 vccd1 sky130_fd_sc_hd__ha_2_16/A sky130_fd_sc_hd__ha_2_16/COUT
+ sky130_fd_sc_hd__fa_2_423/A sky130_fd_sc_hd__ha_2_16/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_27 vssd1 vccd1 la_data_out[45] sky130_fd_sc_hd__ha_2_26/B sky130_fd_sc_hd__ha_2_27/SUM
+ sky130_fd_sc_hd__ha_2_27/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_38 vssd1 vccd1 la_data_out[50] sky130_fd_sc_hd__ha_2_37/B sky130_fd_sc_hd__ha_2_38/SUM
+ sky130_fd_sc_hd__ha_2_38/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__a222oi_1_190 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__nor2_2_5/B
+ sky130_fd_sc_hd__nor2_2_4/B sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__buf_2_4/A
+ sky130_fd_sc_hd__o21ai_1_352/B1 sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__ha_2_49 vssd1 vccd1 sky130_fd_sc_hd__ha_2_49/A sky130_fd_sc_hd__ha_2_47/B
+ sky130_fd_sc_hd__ha_2_49/SUM sky130_fd_sc_hd__ha_2_49/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_360 sky130_fd_sc_hd__fa_2_353/A sky130_fd_sc_hd__fa_2_358/B
+ sky130_fd_sc_hd__fa_2_360/A sky130_fd_sc_hd__fa_2_360/B sky130_fd_sc_hd__fa_2_360/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_371 sky130_fd_sc_hd__fa_2_368/B sky130_fd_sc_hd__fa_2_374/CIN
+ sky130_fd_sc_hd__fa_2_371/A sky130_fd_sc_hd__fa_2_371/B sky130_fd_sc_hd__fa_2_371/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_12 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_8_3/Y
+ sky130_fd_sc_hd__dfxtp_1_122/CLK sky130_fd_sc_hd__clkbuf_1_11/X vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_382 sky130_fd_sc_hd__fa_2_376/CIN sky130_fd_sc_hd__fah_1_11/B
+ sky130_fd_sc_hd__fa_2_382/A sky130_fd_sc_hd__fa_2_382/B sky130_fd_sc_hd__xor2_1_564/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_23 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_2_60/A
+ sky130_fd_sc_hd__dfxtp_1_230/CLK sky130_fd_sc_hd__o21ai_2_3/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_393 sky130_fd_sc_hd__fa_2_391/CIN sky130_fd_sc_hd__fa_2_392/B
+ sky130_fd_sc_hd__fa_2_393/A sky130_fd_sc_hd__fa_2_393/B sky130_fd_sc_hd__xor2_1_584/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_34 sky130_fd_sc_hd__conb_1_145/LO sky130_fd_sc_hd__clkinv_2_12/Y
+ sky130_fd_sc_hd__dfxtp_1_356/CLK sky130_fd_sc_hd__nand4_1_1/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_45 sky130_fd_sc_hd__conb_1_145/LO sky130_fd_sc_hd__clkinv_4_11/Y
+ sky130_fd_sc_hd__dfxtp_1_439/CLK sky130_fd_sc_hd__o31ai_2_0/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_103 sky130_fd_sc_hd__xor2_1_208/X sky130_fd_sc_hd__nor2_1_103/Y
+ sky130_fd_sc_hd__o21ai_1_33/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_114 sky130_fd_sc_hd__nor2_1_114/B sky130_fd_sc_hd__nor2_1_114/Y
+ sky130_fd_sc_hd__nor2_1_114/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_125 sky130_fd_sc_hd__nor2_1_125/B sky130_fd_sc_hd__nor2_1_125/Y
+ sky130_fd_sc_hd__nor2_1_125/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_136 sky130_fd_sc_hd__nor2_1_140/Y sky130_fd_sc_hd__nor2_1_136/Y
+ sky130_fd_sc_hd__nor2_1_144/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_12 sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__dfxtp_1_285/Q sky130_fd_sc_hd__o211ai_1_9/Y sky130_fd_sc_hd__nand2_2_3/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_147 sky130_fd_sc_hd__nor2_1_147/B sky130_fd_sc_hd__nor2_1_147/Y
+ sky130_fd_sc_hd__nor2_1_147/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_23 sky130_fd_sc_hd__nor2_4_0/Y sky130_fd_sc_hd__nor2_2_0/Y
+ sky130_fd_sc_hd__dfxtp_1_329/Q sky130_fd_sc_hd__nor2_1_240/A sky130_fd_sc_hd__nand2_1_16/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_34 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__clkbuf_1_25/X
+ sky130_fd_sc_hd__nand2_1_82/B sky130_fd_sc_hd__dfxtp_1_128/Q sky130_fd_sc_hd__a22oi_1_34/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_158 sky130_fd_sc_hd__nor2_1_161/Y sky130_fd_sc_hd__nor2_1_158/Y
+ sky130_fd_sc_hd__nor2_1_160/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_169 sky130_fd_sc_hd__nor2_1_170/B sky130_fd_sc_hd__nor2_1_169/Y
+ sky130_fd_sc_hd__nor2_1_169/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_45 sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__dfxtp_1_101/Q sky130_fd_sc_hd__dfxtp_1_69/Q sky130_fd_sc_hd__a22oi_1_45/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_56 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__nor2_4_3/Y
+ sky130_fd_sc_hd__nand2_1_71/B sky130_fd_sc_hd__dfxtp_1_139/Q sky130_fd_sc_hd__a22oi_1_56/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_67 sky130_fd_sc_hd__clkbuf_1_24/X sky130_fd_sc_hd__clkbuf_1_23/X
+ sky130_fd_sc_hd__dfxtp_1_112/Q sky130_fd_sc_hd__dfxtp_1_80/Q sky130_fd_sc_hd__a22oi_1_67/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_78 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__nor2_4_3/Y
+ sky130_fd_sc_hd__nand2_1_60/B sky130_fd_sc_hd__dfxtp_1_150/Q sky130_fd_sc_hd__a22oi_1_78/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_89 sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__dfxtp_1_123/Q sky130_fd_sc_hd__dfxtp_1_91/Q sky130_fd_sc_hd__a22oi_1_89/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_310 sky130_fd_sc_hd__buf_12_310/A sky130_fd_sc_hd__buf_12_463/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_321 sky130_fd_sc_hd__buf_12_321/A sky130_fd_sc_hd__buf_12_567/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_332 sky130_fd_sc_hd__buf_12_332/A sky130_fd_sc_hd__buf_12_597/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_343 sky130_fd_sc_hd__buf_12_343/A sky130_fd_sc_hd__buf_12_532/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_202 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__nor2b_1_7/Y sky130_fd_sc_hd__nor2_1_109/Y sky130_fd_sc_hd__a22oi_1_202/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_354 sky130_fd_sc_hd__buf_12_354/A sky130_fd_sc_hd__buf_12_550/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_213 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__buf_2_25/A
+ sky130_fd_sc_hd__nor2b_1_13/Y sky130_fd_sc_hd__nor2_1_167/Y sky130_fd_sc_hd__a22oi_1_213/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_365 sky130_fd_sc_hd__buf_12_78/X sky130_fd_sc_hd__buf_12_528/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_376 sky130_fd_sc_hd__buf_12_376/A sky130_fd_sc_hd__buf_12_468/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_387 sky130_fd_sc_hd__buf_12_387/A sky130_fd_sc_hd__buf_12_559/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_398 sky130_fd_sc_hd__buf_12_398/A sky130_fd_sc_hd__buf_12_470/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_510 sky130_fd_sc_hd__and3_4_9/A sky130_fd_sc_hd__xor2_1_424/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_521 sky130_fd_sc_hd__o21ai_1_658/A2 sky130_fd_sc_hd__xnor2_1_133/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_532 sky130_fd_sc_hd__nor2_1_170/B sky130_fd_sc_hd__nor2_1_172/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_543 sky130_fd_sc_hd__nor2_1_176/B sky130_fd_sc_hd__nand2_1_548/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_106 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_383/A sky130_fd_sc_hd__nor2b_2_4/A
+ sky130_fd_sc_hd__xnor2_1_109/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_554 sky130_fd_sc_hd__a21oi_2_13/B1 sky130_fd_sc_hd__nand2_1_556/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_117 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_117/B sky130_fd_sc_hd__xnor2_1_117/Y
+ sky130_fd_sc_hd__xnor2_1_117/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_565 sky130_fd_sc_hd__nand2_1_570/A sky130_fd_sc_hd__nor2_2_25/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_128 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_128/B sky130_fd_sc_hd__clkbuf_1_9/A
+ sky130_fd_sc_hd__xnor2_1_128/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_576 sky130_fd_sc_hd__nor2_1_190/B sky130_fd_sc_hd__nor2_1_192/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_139 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_139/B sky130_fd_sc_hd__xnor2_1_139/Y
+ sky130_fd_sc_hd__xnor2_1_139/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_587 sky130_fd_sc_hd__nand2_1_612/A sky130_fd_sc_hd__nor2_1_200/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_598 sky130_fd_sc_hd__nand2_1_629/A sky130_fd_sc_hd__nor2_1_210/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_4_12 sky130_fd_sc_hd__ha_2_39/A sky130_fd_sc_hd__inv_2_77/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_23 sky130_fd_sc_hd__nand2_2_4/Y sky130_fd_sc_hd__clkinv_4_23/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_34 sky130_fd_sc_hd__clkinv_4_34/A sky130_fd_sc_hd__buf_8_151/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_90 sky130_fd_sc_hd__buf_6_1/X sky130_fd_sc_hd__nor2_1_90/Y
+ sky130_fd_sc_hd__buf_6_5/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_45 sky130_fd_sc_hd__clkinv_4_45/A sky130_fd_sc_hd__clkinv_4_45/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_56 sky130_fd_sc_hd__clkinv_4_56/A sky130_fd_sc_hd__clkinv_4_56/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_67 sky130_fd_sc_hd__clkinv_4_67/A sky130_fd_sc_hd__clkinv_4_67/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_78 wbs_dat_i[28] sky130_fd_sc_hd__inv_2_195/A vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_1004 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_4_89 wbs_dat_i[8] sky130_fd_sc_hd__clkinv_4_89/Y vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_1015 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1026 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1037 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1048 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1059 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21a_1_0 sky130_fd_sc_hd__o21a_1_0/X sky130_fd_sc_hd__or2_0_5/A
+ sky130_fd_sc_hd__o21a_1_0/B1 sky130_fd_sc_hd__o21a_1_0/A2 vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__decap_12_550 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_561 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_572 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_583 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_594 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_306 sky130_fd_sc_hd__fa_2_250/A sky130_fd_sc_hd__xor2_1_306/X
+ sky130_fd_sc_hd__xor2_1_306/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_317 sky130_fd_sc_hd__fa_2_217/A sky130_fd_sc_hd__and3_4_14/A
+ sky130_fd_sc_hd__xor2_1_317/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_328 sky130_fd_sc_hd__fa_2_250/A sky130_fd_sc_hd__fa_2_227/A
+ sky130_fd_sc_hd__xor2_1_328/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_339 sky130_fd_sc_hd__fa_2_262/A sky130_fd_sc_hd__fa_2_237/B
+ sky130_fd_sc_hd__xor2_1_339/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nor2b_1_80 sky130_fd_sc_hd__or2_0_82/A sky130_fd_sc_hd__fa_2_491/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_91 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_91/Y
+ sky130_fd_sc_hd__nor2b_1_91/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1080 sky130_fd_sc_hd__maj3_1_0/C sky130_fd_sc_hd__ha_2_51/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1091 sky130_fd_sc_hd__a22o_1_71/B1 sky130_fd_sc_hd__and2_4_0/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1560 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1571 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1582 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1593 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_14 sky130_fd_sc_hd__buf_2_192/A sky130_fd_sc_hd__dfxtp_1_8/CLK
+ sky130_fd_sc_hd__dfxtp_1_14/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_25 sky130_fd_sc_hd__ha_2_6/A sky130_fd_sc_hd__dfxtp_1_29/CLK
+ sky130_fd_sc_hd__ha_2_43/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_36 sky130_fd_sc_hd__nand2_1_78/B sky130_fd_sc_hd__dfxtp_1_45/CLK
+ sky130_fd_sc_hd__dfxtp_1_36/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_190 sky130_fd_sc_hd__fa_2_184/CIN sky130_fd_sc_hd__fa_2_190/SUM
+ sky130_fd_sc_hd__fa_2_190/A sky130_fd_sc_hd__fa_2_190/B sky130_fd_sc_hd__xor2_1_279/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_47 sky130_fd_sc_hd__nand2_1_67/B sky130_fd_sc_hd__dfxtp_1_51/CLK
+ sky130_fd_sc_hd__dfxtp_1_47/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_58 sky130_fd_sc_hd__nand2_1_54/B sky130_fd_sc_hd__dfxtp_1_62/CLK
+ sky130_fd_sc_hd__dfxtp_1_58/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_69 sky130_fd_sc_hd__dfxtp_1_69/Q sky130_fd_sc_hd__dfxtp_1_72/CLK
+ sky130_fd_sc_hd__dfxtp_1_69/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_308 vccd1 vssd1 sky130_fd_sc_hd__and2_0_308/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_308/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_319 vccd1 vssd1 sky130_fd_sc_hd__and2_0_319/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_319/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__inv_2_108 sky130_fd_sc_hd__inv_2_108/A sky130_fd_sc_hd__inv_2_108/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_119 sky130_fd_sc_hd__inv_2_120/A sky130_fd_sc_hd__buf_8_67/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_sram_1kbyte_1rw1r_32x256_8_4 sky130_fd_sc_hd__inv_8_1/Y sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__buf_12_584/X sky130_fd_sc_hd__buf_12_179/X sky130_fd_sc_hd__buf_12_603/X
+ sky130_fd_sc_hd__buf_12_664/X sky130_fd_sc_hd__buf_12_598/X sky130_fd_sc_hd__buf_12_659/X
+ sky130_fd_sc_hd__buf_12_595/X sky130_fd_sc_hd__clkinv_4_21/Y sky130_fd_sc_hd__buf_12_609/X
+ sky130_fd_sc_hd__buf_12_587/X sky130_fd_sc_hd__buf_12_588/X vccd1 sky130_fd_sc_hd__clkinv_4_37/Y
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[16] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[17]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[18] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[19]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[20] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[21]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[22] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[23]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[24] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[25]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[26] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[27]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[28] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[29]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[30] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[31]
+ sky130_fd_sc_hd__buf_12_560/X sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[1] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[2]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[3] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[4]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[5] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[6]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[7] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[8]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[9] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[10]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[11] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[12]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[13] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[14]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[15] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout1[0]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[10] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[11]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[12] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[13]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[14] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[15]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[16] sky130_fd_sc_hd__buf_12_550/X sky130_fd_sc_hd__buf_12_124/X
+ sky130_fd_sc_hd__buf_12_101/X sky130_fd_sc_hd__buf_12_167/X sky130_fd_sc_hd__buf_12_293/X
+ sky130_fd_sc_hd__clkinv_4_38/Y sky130_fd_sc_hd__buf_6_8/X sky130_fd_sc_hd__buf_6_8/X
+ sky130_fd_sc_hd__buf_6_8/X sky130_fd_sc_hd__buf_6_8/X sky130_fd_sc_hd__buf_6_8/X
+ sky130_fd_sc_hd__buf_6_8/X sky130_fd_sc_hd__buf_6_8/X sky130_fd_sc_hd__buf_6_8/X
+ sky130_fd_sc_hd__buf_6_8/X sky130_fd_sc_hd__buf_6_8/X sky130_fd_sc_hd__buf_6_8/X
+ sky130_fd_sc_hd__buf_6_8/X sky130_fd_sc_hd__clkbuf_4_18/X sky130_fd_sc_hd__clkbuf_4_18/X
+ sky130_fd_sc_hd__clkbuf_4_18/X sky130_fd_sc_hd__clkbuf_4_18/X sky130_fd_sc_hd__clkbuf_4_18/X
+ sky130_fd_sc_hd__clkbuf_4_18/X sky130_fd_sc_hd__clkbuf_4_18/X sky130_fd_sc_hd__buf_2_137/A
+ sky130_fd_sc_hd__buf_2_137/A sky130_fd_sc_hd__buf_2_137/A sky130_fd_sc_hd__buf_2_137/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[0] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[1]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[2] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[3]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[4] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[5]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[6] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[7]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[8] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[9]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[25] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[26]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[27] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[28]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[29] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[30]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[31] sky130_fd_sc_hd__buf_2_137/X sky130_fd_sc_hd__buf_2_137/A
+ sky130_fd_sc_hd__buf_2_137/A sky130_fd_sc_hd__buf_2_137/A sky130_fd_sc_hd__buf_2_137/X
+ sky130_fd_sc_hd__buf_2_137/X sky130_fd_sc_hd__buf_2_137/X sky130_fd_sc_hd__buf_2_137/X
+ sky130_fd_sc_hd__buf_2_137/X sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[17] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[18]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[19] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[20]
+ sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[21] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[22]
+ sky130_fd_sc_hd__buf_12_581/X sky130_fd_sc_hd__buf_12_511/X sky130_fd_sc_hd__buf_12_476/X
+ sky130_fd_sc_hd__buf_12_575/X sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[23] sky130_sram_1kbyte_1rw1r_32x256_8_4/dout0[24]
+ vssd1 vssd1 sky130_sram_1kbyte_1rw1r_32x256_8
Xsky130_fd_sc_hd__buf_12_140 sky130_fd_sc_hd__buf_8_8/X sky130_fd_sc_hd__buf_12_358/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_151 sky130_fd_sc_hd__buf_12_49/X sky130_fd_sc_hd__buf_12_309/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_162 sky130_fd_sc_hd__buf_8_32/X sky130_fd_sc_hd__buf_12_162/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_173 sky130_fd_sc_hd__buf_8_55/X sky130_fd_sc_hd__buf_12_422/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_184 sky130_fd_sc_hd__buf_8_14/X sky130_fd_sc_hd__buf_12_431/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_195 sky130_fd_sc_hd__buf_4_27/X sky130_fd_sc_hd__buf_12_438/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_340 sky130_fd_sc_hd__a21oi_2_2/B1 sky130_fd_sc_hd__nand2_1_202/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_351 sky130_fd_sc_hd__o21ai_1_280/B1 sky130_fd_sc_hd__o21ai_1_281/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_362 sky130_fd_sc_hd__nand2_1_236/A sky130_fd_sc_hd__nor2_2_3/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_373 sky130_fd_sc_hd__a21oi_1_55/B1 sky130_fd_sc_hd__nand2_1_260/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_384 sky130_fd_sc_hd__xor2_1_171/A sky130_fd_sc_hd__o21ai_1_360/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_395 sky130_fd_sc_hd__xnor2_1_56/B sky130_fd_sc_hd__a21oi_1_65/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_2_3 sky130_fd_sc_hd__a21oi_2_3/B1 sky130_fd_sc_hd__or2_0_6/X
+ sky130_fd_sc_hd__xnor2_1_23/B sky130_fd_sc_hd__xor2_1_83/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_2
Xsky130_fd_sc_hd__a211o_1_9 vssd1 vccd1 sky130_fd_sc_hd__fa_2_270/B sky130_fd_sc_hd__dfxtp_1_72/Q
+ sky130_fd_sc_hd__nor2_1_13/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_9/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__o21ai_1_309 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_0/A sky130_fd_sc_hd__nor2_1_73/Y
+ sky130_fd_sc_hd__nand2_1_239/Y sky130_fd_sc_hd__xnor2_1_33/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__conb_1_108 sky130_fd_sc_hd__conb_1_108/LO sky130_fd_sc_hd__conb_1_108/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_119 sky130_fd_sc_hd__conb_1_119/LO sky130_fd_sc_hd__conb_1_119/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_380 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_391 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_103 sky130_fd_sc_hd__fa_2_75/A sky130_fd_sc_hd__fa_2_75/CIN
+ sky130_fd_sc_hd__xor2_1_103/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_114 sky130_fd_sc_hd__fa_2_97/A sky130_fd_sc_hd__fa_2_82/CIN
+ sky130_fd_sc_hd__xor2_1_114/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_125 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__fa_2_95/CIN
+ sky130_fd_sc_hd__xor2_1_125/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_136 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__fa_2_99/A
+ sky130_fd_sc_hd__xor2_1_136/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_147 sky130_fd_sc_hd__fa_2_122/A sky130_fd_sc_hd__fa_2_112/B
+ sky130_fd_sc_hd__xor2_1_147/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_158 sky130_fd_sc_hd__fa_2_122/A sky130_fd_sc_hd__xor2_1_158/X
+ sky130_fd_sc_hd__xor2_1_158/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_509 sky130_fd_sc_hd__ha_2_46/B sky130_fd_sc_hd__dfxtp_1_509/CLK
+ sky130_fd_sc_hd__and2_0_391/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_169 sky130_fd_sc_hd__fa_2_122/A sky130_fd_sc_hd__xor2_1_169/X
+ sky130_fd_sc_hd__xor2_1_169/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_107 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_53/A1 sky130_fd_sc_hd__clkbuf_1_107/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_118 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_118/X sky130_fd_sc_hd__inv_2_3/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o21ai_1_810 vssd1 vccd1 sky130_fd_sc_hd__inv_2_48/Y sky130_fd_sc_hd__nand2b_2_6/Y
+ sky130_fd_sc_hd__o21ai_1_810/B1 sky130_fd_sc_hd__xor2_1_585/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1390 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_129 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_129/X sky130_fd_sc_hd__inv_4_0/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o21ai_1_821 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_2/Y sky130_fd_sc_hd__nand2b_2_6/Y
+ sky130_fd_sc_hd__o21ai_1_821/B1 sky130_fd_sc_hd__xor2_1_594/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_832 vssd1 vccd1 sky130_fd_sc_hd__inv_2_44/Y sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_832/B1 sky130_fd_sc_hd__xor2_1_606/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_843 vssd1 vccd1 sky130_fd_sc_hd__inv_2_48/Y sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_843/B1 sky130_fd_sc_hd__xor2_1_615/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_9 sky130_fd_sc_hd__buf_8_5/A sky130_fd_sc_hd__dfxtp_1_9/CLK
+ sky130_fd_sc_hd__dfxtp_1_9/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_854 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_2/A sky130_fd_sc_hd__nor2_1_218/Y
+ sky130_fd_sc_hd__nand2_1_653/Y sky130_fd_sc_hd__xnor2_1_183/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_865 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_643/A sky130_fd_sc_hd__nor2_1_224/Y
+ sky130_fd_sc_hd__nand2_1_677/Y sky130_fd_sc_hd__xnor2_1_191/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_876 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_237/Y sky130_fd_sc_hd__nand2_1_735/Y
+ sky130_fd_sc_hd__nand2_1_733/Y sky130_fd_sc_hd__o21ai_1_876/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_887 vssd1 vccd1 sky130_fd_sc_hd__nand2_1_779/Y sky130_fd_sc_hd__a21oi_1_166/Y
+ sky130_fd_sc_hd__a21oi_1_165/Y sky130_fd_sc_hd__o21ai_1_887/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_898 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_681/A sky130_fd_sc_hd__nor2_1_259/Y
+ sky130_fd_sc_hd__nand2_1_813/Y sky130_fd_sc_hd__xnor2_1_295/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nand2b_2_0 sky130_fd_sc_hd__nor2_2_9/B sky130_fd_sc_hd__nand2b_2_0/Y
+ sky130_fd_sc_hd__nor2_2_9/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_2
Xsky130_fd_sc_hd__inv_4_19 sky130_fd_sc_hd__inv_4_19/Y wbs_dat_i[13] vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__xor2_1_670 la_data_out[84] sky130_fd_sc_hd__xor2_1_670/X la_data_out[85]
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_681 sky130_fd_sc_hd__xor2_1_681/B sky130_fd_sc_hd__xor2_1_681/X
+ sky130_fd_sc_hd__xor2_1_681/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_692 sky130_fd_sc_hd__or4_1_3/B sky130_fd_sc_hd__xor2_1_692/X
+ sky130_fd_sc_hd__xor2_1_692/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__and2_0_105 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_95/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_105/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_13 la_data_out[114] sky130_fd_sc_hd__conb_1_129/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_116 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_66/D sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_116/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_24 la_data_out[103] sky130_fd_sc_hd__conb_1_118/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_127 vccd1 vssd1 sky130_fd_sc_hd__and2_0_127/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_127/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_35 la_data_out[28] sky130_fd_sc_hd__conb_1_107/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_138 vccd1 vssd1 sky130_fd_sc_hd__and2_0_138/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_138/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_46 la_data_out[17] sky130_fd_sc_hd__conb_1_96/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_149 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_72/D sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_149/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_57 la_data_out[6] sky130_fd_sc_hd__conb_1_85/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__fa_2_0 sky130_fd_sc_hd__xor2_1_0/B sky130_fd_sc_hd__or2_0_0/B sky130_fd_sc_hd__fa_2_0/A
+ sky130_fd_sc_hd__fa_2_0/B sky130_fd_sc_hd__fa_2_5/SUM vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_1_68 io_out[33] sky130_fd_sc_hd__conb_1_74/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_79 io_out[22] sky130_fd_sc_hd__conb_1_63/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_170 sky130_fd_sc_hd__nor2_1_28/A sky130_fd_sc_hd__dfxtp_1_151/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_2 sky130_fd_sc_hd__buf_8_2/A sky130_fd_sc_hd__buf_8_2/X vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__a22o_1_4 sky130_fd_sc_hd__nand2_1_7/B sky130_fd_sc_hd__mux2_2_18/X
+ sky130_fd_sc_hd__buf_6_0/A sky130_fd_sc_hd__mux2_2_37/X sky130_fd_sc_hd__nand2_1_8/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_181 sky130_fd_sc_hd__o22ai_1_42/B1 sky130_fd_sc_hd__dfxtp_1_180/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_192 sky130_fd_sc_hd__o22ai_1_18/B1 sky130_fd_sc_hd__dfxtp_1_113/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_50 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__buf_2_124/X
+ sky130_fd_sc_hd__a22o_1_50/X sky130_fd_sc_hd__a22o_1_50/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_61 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__and2_0_361/A
+ sky130_fd_sc_hd__a22o_1_61/X sky130_fd_sc_hd__ha_2_32/SUM sky130_fd_sc_hd__a22o_1_71/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_72 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__buf_2_180/X
+ sky130_fd_sc_hd__a22o_1_72/X sky130_fd_sc_hd__xor2_1_689/X sky130_fd_sc_hd__nor2_1_269/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__nand4_1_0 sky130_fd_sc_hd__nand4_1_0/C sky130_fd_sc_hd__nand4_1_0/B
+ sky130_fd_sc_hd__nand4_1_0/Y sky130_fd_sc_hd__nand4_1_0/D sky130_fd_sc_hd__nor4_1_0/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__o21ai_1_106 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_109/A2 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_120/Y sky130_fd_sc_hd__and2_0_170/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_117 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_117/A2 sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__a22oi_1_169/Y sky130_fd_sc_hd__and2_0_157/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_128 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_129/A2 sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__a22oi_1_174/Y sky130_fd_sc_hd__and2_0_143/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_139 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_141/A2 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_137/Y sky130_fd_sc_hd__and2_0_129/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__inv_8_2 sky130_fd_sc_hd__inv_8_2/A sky130_fd_sc_hd__inv_8_2/Y vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__inv_8
Xsky130_fd_sc_hd__nand2_1_40 sky130_fd_sc_hd__buf_6_2/A sky130_fd_sc_hd__nand2_1_41/Y
+ sky130_fd_sc_hd__nand2_1_42/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_51 sky130_fd_sc_hd__o21ai_2_3/A2 sky130_fd_sc_hd__ha_2_9/B
+ sky130_fd_sc_hd__nor2b_1_1/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_62 sky130_fd_sc_hd__nand2_1_62/Y sky130_fd_sc_hd__nand2_1_62/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_73 sky130_fd_sc_hd__nand2_1_73/Y sky130_fd_sc_hd__nand2_1_73/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_84 sky130_fd_sc_hd__nand2_1_84/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__xor2_2_1/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_95 sky130_fd_sc_hd__nand2_1_95/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__xnor2_1_78/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_306 sky130_fd_sc_hd__dfxtp_1_306/Q sky130_fd_sc_hd__clkinv_8_6/Y
+ sky130_fd_sc_hd__and2_0_282/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_317 sky130_fd_sc_hd__or2_0_90/A sky130_fd_sc_hd__dfxtp_1_319/CLK
+ sky130_fd_sc_hd__and2_0_294/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_328 sky130_fd_sc_hd__dfxtp_1_328/Q sky130_fd_sc_hd__dfxtp_1_343/CLK
+ sky130_fd_sc_hd__and2_0_316/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_339 sky130_fd_sc_hd__a22oi_1_3/B2 sky130_fd_sc_hd__dfxtp_1_339/CLK
+ sky130_fd_sc_hd__and2_0_322/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_640 vssd1 vccd1 sky130_fd_sc_hd__buf_2_12/X sky130_fd_sc_hd__nand2b_1_19/Y
+ sky130_fd_sc_hd__o21ai_1_640/B1 sky130_fd_sc_hd__xor2_1_428/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_651 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_168/Y sky130_fd_sc_hd__nor2_1_165/A
+ sky130_fd_sc_hd__nor2_1_164/Y sky130_fd_sc_hd__o21ai_1_651/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_662 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_2/Y sky130_fd_sc_hd__nand2b_1_18/Y
+ sky130_fd_sc_hd__o21ai_1_662/B1 sky130_fd_sc_hd__xor2_1_445/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_673 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_681/A2 sky130_fd_sc_hd__nor2_1_169/A
+ sky130_fd_sc_hd__nor2_1_168/Y sky130_fd_sc_hd__o21ai_1_673/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_684 vssd1 vccd1 sky130_fd_sc_hd__inv_2_46/Y sky130_fd_sc_hd__nand2b_1_19/Y
+ sky130_fd_sc_hd__o21ai_1_684/B1 sky130_fd_sc_hd__xor2_1_463/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_695 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_2/Y sky130_fd_sc_hd__nand2b_1_19/Y
+ sky130_fd_sc_hd__o21ai_1_695/B1 sky130_fd_sc_hd__xor2_1_473/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_14 sky130_fd_sc_hd__fa_2_5/A sky130_fd_sc_hd__fa_2_15/B sky130_fd_sc_hd__fa_2_14/A
+ sky130_fd_sc_hd__fa_2_14/B sky130_fd_sc_hd__fa_2_14/CIN vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_25 sky130_fd_sc_hd__fa_2_17/B sky130_fd_sc_hd__fa_2_25/SUM
+ sky130_fd_sc_hd__fa_2_25/A sky130_fd_sc_hd__fa_2_25/B sky130_fd_sc_hd__fa_2_26/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_36 sky130_fd_sc_hd__fa_2_34/CIN sky130_fd_sc_hd__fa_2_42/B
+ sky130_fd_sc_hd__fa_2_36/A sky130_fd_sc_hd__fa_2_36/B sky130_fd_sc_hd__xor2_1_61/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_47 sky130_fd_sc_hd__fa_2_43/B sky130_fd_sc_hd__fa_2_51/CIN
+ sky130_fd_sc_hd__fa_2_47/A sky130_fd_sc_hd__fa_2_47/B sky130_fd_sc_hd__fa_2_47/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_58 sky130_fd_sc_hd__fa_2_50/A sky130_fd_sc_hd__fa_2_57/B sky130_fd_sc_hd__fa_2_58/A
+ sky130_fd_sc_hd__fa_2_58/B sky130_fd_sc_hd__fa_2_58/CIN vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_69 sky130_fd_sc_hd__fa_2_62/A sky130_fd_sc_hd__fa_2_68/B sky130_fd_sc_hd__fa_2_69/A
+ sky130_fd_sc_hd__fa_2_69/B sky130_fd_sc_hd__xor2_1_93/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_206 vccd1 vssd1 sky130_fd_sc_hd__xnor2_2_5/A sky130_fd_sc_hd__mux2_2_49/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__a222oi_1_520 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__buf_2_27/X
+ sky130_fd_sc_hd__buf_2_15/X sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__buf_2_4/A
+ sky130_fd_sc_hd__o21ai_1_820/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_531 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__buf_2_27/X
+ sky130_fd_sc_hd__buf_2_15/X sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__buf_2_4/A
+ sky130_fd_sc_hd__o21ai_1_838/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_542 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__inv_6_0/Y sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__o21ai_1_856/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_553 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_417/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_449/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_750/A sky130_fd_sc_hd__dfxtp_1_385/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a21oi_1_19 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_48/Y
+ sky130_fd_sc_hd__a21oi_1_19/Y sky130_fd_sc_hd__dfxtp_1_78/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_564 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_406/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_438/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_761/A sky130_fd_sc_hd__dfxtp_1_374/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_575 vccd1 vssd1 sky130_fd_sc_hd__inv_2_68/Y sky130_fd_sc_hd__dfxtp_1_427/Q
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__ha_2_9/A sky130_fd_sc_hd__dfxtp_1_459/Q
+ sky130_fd_sc_hd__clkinv_1_772/A sky130_fd_sc_hd__dfxtp_1_395/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_586 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_408/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_440/Q sky130_fd_sc_hd__clkbuf_1_32/X
+ sky130_fd_sc_hd__clkinv_1_783/A sky130_fd_sc_hd__dfxtp_1_376/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_597 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_415/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_447/Q sky130_fd_sc_hd__nor2_4_19/B
+ sky130_fd_sc_hd__clkinv_1_794/A sky130_fd_sc_hd__dfxtp_1_383/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_15 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_120 sky130_fd_sc_hd__and2_0_342/A sky130_fd_sc_hd__and2_0_391/A
+ sky130_fd_sc_hd__ha_2_46/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__decap_12_26 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_131 sky130_fd_sc_hd__clkinv_4_50/Y sky130_fd_sc_hd__nor2b_1_131/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__decap_12_37 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_142 sky130_fd_sc_hd__clkinv_4_61/Y sky130_fd_sc_hd__nor2b_1_142/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__decap_12_48 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_153 sky130_fd_sc_hd__clkinv_4_72/Y sky130_fd_sc_hd__nor2b_1_153/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__decap_12_59 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__fah_1_11 sky130_fd_sc_hd__fa_2_378/A sky130_fd_sc_hd__fah_1_11/B
+ sky130_fd_sc_hd__fah_1_11/A sky130_fd_sc_hd__fa_2_381/B sky130_fd_sc_hd__fah_1_11/CI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__fah_1
Xsky130_fd_sc_hd__buf_6_15 vccd1 vssd1 sky130_fd_sc_hd__buf_6_15/X sky130_fd_sc_hd__buf_6_15/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_26 vccd1 vssd1 sky130_fd_sc_hd__buf_6_26/X sky130_fd_sc_hd__buf_6_26/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_37 vccd1 vssd1 sky130_fd_sc_hd__buf_6_37/X sky130_fd_sc_hd__buf_8_83/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_48 vccd1 vssd1 sky130_fd_sc_hd__buf_6_48/X sky130_fd_sc_hd__buf_8_7/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_59 vccd1 vssd1 sky130_fd_sc_hd__buf_6_59/X sky130_fd_sc_hd__buf_6_59/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_17 sky130_fd_sc_hd__clkinv_4_68/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_28 sky130_fd_sc_hd__clkinv_4_70/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_39 sky130_fd_sc_hd__buf_2_193/A vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__nand2_1_307 sky130_fd_sc_hd__nand2_1_307/Y sky130_fd_sc_hd__buf_4_6/X
+ sky130_fd_sc_hd__buf_8_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_906 sky130_fd_sc_hd__clkinv_1_907/A sky130_fd_sc_hd__buf_2_48/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_0 sky130_fd_sc_hd__nor2_2_1/B sky130_fd_sc_hd__nor2_1_0/Y
+ sky130_fd_sc_hd__nor2_1_0/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nand2_1_318 sky130_fd_sc_hd__o21a_1_1/B1 sky130_fd_sc_hd__o21ai_1_32/Y
+ sky130_fd_sc_hd__xor2_1_210/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_917 sky130_fd_sc_hd__clkinv_1_917/Y sky130_fd_sc_hd__clkinv_1_917/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_329 sky130_fd_sc_hd__nand2_1_329/Y sky130_fd_sc_hd__nor2_4_12/Y
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_928 sky130_fd_sc_hd__buf_2_159/A sky130_fd_sc_hd__inv_6_1/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__bufinv_8_2 sky130_fd_sc_hd__bufinv_8_2/A sky130_fd_sc_hd__bufinv_8_2/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__bufinv_8
Xsky130_fd_sc_hd__clkinv_1_939 sky130_fd_sc_hd__buf_8_93/A sky130_fd_sc_hd__inv_1_0/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_103 sky130_fd_sc_hd__dfxtp_1_103/Q sky130_fd_sc_hd__dfxtp_1_105/CLK
+ sky130_fd_sc_hd__and2_0_143/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_114 sky130_fd_sc_hd__dfxtp_1_114/Q sky130_fd_sc_hd__dfxtp_1_97/CLK
+ sky130_fd_sc_hd__and2_0_197/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_125 sky130_fd_sc_hd__dfxtp_1_125/Q sky130_fd_sc_hd__dfxtp_1_126/CLK
+ sky130_fd_sc_hd__and2_0_5/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_136 sky130_fd_sc_hd__dfxtp_1_136/Q sky130_fd_sc_hd__dfxtp_1_138/CLK
+ sky130_fd_sc_hd__and2_0_151/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_147 sky130_fd_sc_hd__dfxtp_1_147/Q sky130_fd_sc_hd__dfxtp_1_152/CLK
+ sky130_fd_sc_hd__and2_0_206/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_158 sky130_fd_sc_hd__dfxtp_1_158/Q sky130_fd_sc_hd__dfxtp_1_158/CLK
+ sky130_fd_sc_hd__and2_0_251/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_169 sky130_fd_sc_hd__dfxtp_1_169/Q sky130_fd_sc_hd__dfxtp_1_170/CLK
+ sky130_fd_sc_hd__and2_0_152/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_470 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_496/A2 sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_470/B1 sky130_fd_sc_hd__xor2_1_273/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_481 vssd1 vccd1 sky130_fd_sc_hd__nand2_2_12/Y sky130_fd_sc_hd__nand2b_1_12/Y
+ sky130_fd_sc_hd__a22oi_1_204/Y sky130_fd_sc_hd__xor2_1_282/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_492 vssd1 vccd1 sky130_fd_sc_hd__inv_2_35/Y sky130_fd_sc_hd__nand2b_2_3/Y
+ sky130_fd_sc_hd__o21ai_1_492/B1 sky130_fd_sc_hd__xor2_1_293/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_902 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_913 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_924 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_935 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_946 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_830 sky130_fd_sc_hd__xnor2_1_300/A sky130_fd_sc_hd__nand2_1_831/Y
+ sky130_fd_sc_hd__or2_0_109/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_957 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_841 sky130_fd_sc_hd__nand2_1_841/Y sky130_fd_sc_hd__nor2b_1_86/Y
+ sky130_fd_sc_hd__ha_2_18/SUM vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_968 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_852 sky130_fd_sc_hd__o21ai_2_18/A2 sky130_fd_sc_hd__nand3_1_5/B
+ la_data_out[36] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_979 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_863 sky130_fd_sc_hd__nor3_1_5/C wbs_adr_i[28] wbs_adr_i[29]
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o21ai_1_30 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_3/B1 sky130_fd_sc_hd__inv_2_53/A
+ sky130_fd_sc_hd__o21ai_1_30/B1 sky130_fd_sc_hd__fa_2_141/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_41 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_41/A2 sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_41/B1 sky130_fd_sc_hd__and2_0_5/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_52 vssd1 vccd1 sky130_fd_sc_hd__inv_2_59/Y sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_52/B1 sky130_fd_sc_hd__o21ai_1_52/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_63 vssd1 vccd1 sky130_fd_sc_hd__inv_2_55/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_99/Y sky130_fd_sc_hd__o21ai_1_63/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_74 vssd1 vccd1 sky130_fd_sc_hd__inv_2_61/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__o21ai_1_74/B1 sky130_fd_sc_hd__o21ai_1_74/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_85 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_85/A2 sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_85/B1 sky130_fd_sc_hd__o21ai_1_85/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_96 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_99/A2 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__o21ai_1_96/B1 sky130_fd_sc_hd__o21ai_1_96/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nand2_4_1 sky130_fd_sc_hd__buf_4_0/A sky130_fd_sc_hd__nand2_4_1/A
+ sky130_fd_sc_hd__nand2_4_1/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_4
Xsky130_fd_sc_hd__a222oi_1_350 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__and2_0_38/A sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__and2_0_49/A
+ sky130_fd_sc_hd__o21ai_1_578/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_290 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_290/X sky130_fd_sc_hd__clkbuf_1_290/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_361 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__buf_4_7/X
+ sky130_fd_sc_hd__buf_4_0/X sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__buf_2_23/X
+ sky130_fd_sc_hd__o21ai_1_596/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_372 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__inv_6_0/Y sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__o21ai_1_615/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_383 vccd1 vssd1 sky130_fd_sc_hd__and3_4_24/X sky130_fd_sc_hd__buf_2_31/X
+ sky130_fd_sc_hd__buf_2_4/A sky130_fd_sc_hd__nor2_1_183/Y sky130_fd_sc_hd__buf_2_20/X
+ sky130_fd_sc_hd__o21ai_1_644/B1 sky130_fd_sc_hd__nor2b_1_16/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_394 vccd1 vssd1 sky130_fd_sc_hd__and3_4_18/X sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__nor2_1_73/B sky130_fd_sc_hd__nor2_2_32/Y sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__o21ai_1_657/B1 sky130_fd_sc_hd__nor2b_2_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__buf_12_503 sky130_fd_sc_hd__buf_12_503/A sky130_fd_sc_hd__buf_12_654/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_514 sky130_fd_sc_hd__buf_12_514/A sky130_fd_sc_hd__buf_12_675/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_525 sky130_fd_sc_hd__buf_12_525/A sky130_fd_sc_hd__buf_12_525/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_536 sky130_fd_sc_hd__buf_12_536/A sky130_fd_sc_hd__buf_12_677/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_547 sky130_fd_sc_hd__buf_12_547/A sky130_fd_sc_hd__buf_12_547/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_558 sky130_fd_sc_hd__buf_12_558/A sky130_fd_sc_hd__buf_12_558/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_569 sky130_fd_sc_hd__buf_12_569/A sky130_fd_sc_hd__buf_12_569/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_209 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_104 sky130_fd_sc_hd__o21ai_1_74/B1 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__xor2_1_313/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_703 sky130_fd_sc_hd__clkinv_1_703/Y sky130_fd_sc_hd__buf_2_16/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_115 sky130_fd_sc_hd__o21ai_1_95/B1 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__xor2_1_359/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_714 sky130_fd_sc_hd__nor2b_1_93/A sky130_fd_sc_hd__xnor2_1_290/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_126 sky130_fd_sc_hd__nand2_1_126/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_127/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_725 sky130_fd_sc_hd__nor2b_1_104/A sky130_fd_sc_hd__xor2_1_681/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_137 sky130_fd_sc_hd__nand2_1_137/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__xor2_1_411/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_736 sky130_fd_sc_hd__nor2b_1_115/A sky130_fd_sc_hd__xnor2_1_301/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_148 sky130_fd_sc_hd__nand2_1_148/Y sky130_fd_sc_hd__xnor2_1_125/Y
+ sky130_fd_sc_hd__nor2_1_2/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_747 sky130_fd_sc_hd__fa_2_470/A sky130_fd_sc_hd__clkinv_1_747/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_159 sky130_fd_sc_hd__nand2_1_159/Y sky130_fd_sc_hd__nor2_2_9/Y
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_758 sky130_fd_sc_hd__fa_2_481/A sky130_fd_sc_hd__clkinv_1_758/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_769 sky130_fd_sc_hd__fa_2_492/A sky130_fd_sc_hd__clkinv_1_769/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__or2_0_101 sky130_fd_sc_hd__or2_0_101/A sky130_fd_sc_hd__or2_0_101/X
+ sky130_fd_sc_hd__or2_0_101/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_112 sky130_fd_sc_hd__or2_0_112/A sky130_fd_sc_hd__or2_0_112/X
+ sky130_fd_sc_hd__or2_0_112/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__decap_12_1208 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_8 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__xor3_1_9/C
+ sky130_fd_sc_hd__xor2_1_8/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1219 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_8_6 sky130_fd_sc_hd__clkinv_8_6/Y sky130_fd_sc_hd__clkinv_8_6/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_12_710 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_721 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_732 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_743 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_754 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_765 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_776 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_660 sky130_fd_sc_hd__xnor2_1_187/A sky130_fd_sc_hd__nand2_1_661/Y
+ sky130_fd_sc_hd__or2_0_70/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_787 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_671 sky130_fd_sc_hd__nand2_1_671/Y sky130_fd_sc_hd__or2_0_75/A
+ sky130_fd_sc_hd__or2_0_75/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_798 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_682 sky130_fd_sc_hd__xnor2_1_193/A sky130_fd_sc_hd__nand2_1_683/Y
+ sky130_fd_sc_hd__or2_0_77/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_693 sky130_fd_sc_hd__nand2_1_693/Y sky130_fd_sc_hd__mux2_2_31/X
+ sky130_fd_sc_hd__mux2_2_46/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_1720 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1731 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_30 sky130_fd_sc_hd__inv_2_30/A sky130_fd_sc_hd__inv_2_30/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1742 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_41 sky130_fd_sc_hd__inv_2_41/A sky130_fd_sc_hd__inv_2_41/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1753 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_52 sky130_fd_sc_hd__inv_2_52/A sky130_fd_sc_hd__inv_2_52/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1764 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_63 sky130_fd_sc_hd__inv_2_63/A sky130_fd_sc_hd__inv_2_63/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1775 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_74 sky130_fd_sc_hd__inv_2_74/A sky130_fd_sc_hd__inv_2_74/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1786 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_85 la_data_out[43] sky130_fd_sc_hd__inv_2_86/A vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1797 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_96 sky130_fd_sc_hd__inv_4_15/Y sky130_fd_sc_hd__inv_2_96/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__ha_2_17 vssd1 vccd1 sky130_fd_sc_hd__ha_2_17/A sky130_fd_sc_hd__ha_2_17/COUT
+ sky130_fd_sc_hd__fa_2_452/B sky130_fd_sc_hd__ha_2_17/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_28 vssd1 vccd1 la_data_out[44] sky130_fd_sc_hd__ha_2_27/B sky130_fd_sc_hd__ha_2_28/SUM
+ sky130_fd_sc_hd__ha_2_28/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__a222oi_1_180 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__buf_2_4/A
+ sky130_fd_sc_hd__buf_6_5/X sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__o21ai_1_337/B1 sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__ha_2_39 vssd1 vccd1 sky130_fd_sc_hd__ha_2_39/A sky130_fd_sc_hd__ha_2_38/B
+ sky130_fd_sc_hd__ha_2_39/SUM la_data_out[48] vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__a222oi_1_191 vccd1 vssd1 sky130_fd_sc_hd__and3_4_1/X sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__buf_2_32/X sky130_fd_sc_hd__nor2_2_9/Y sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__o21ai_1_353/B1 sky130_fd_sc_hd__and2b_4_3/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_350 sky130_fd_sc_hd__fa_2_345/B sky130_fd_sc_hd__fa_2_352/B
+ sky130_fd_sc_hd__fa_2_350/A sky130_fd_sc_hd__fa_2_350/B sky130_fd_sc_hd__xor2_1_518/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_361 sky130_fd_sc_hd__fa_2_349/B sky130_fd_sc_hd__fa_2_361/SUM
+ sky130_fd_sc_hd__fa_2_361/A sky130_fd_sc_hd__fa_2_361/B sky130_fd_sc_hd__xor2_1_532/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_372 sky130_fd_sc_hd__fa_2_364/B sky130_fd_sc_hd__fa_2_373/A
+ sky130_fd_sc_hd__fa_2_372/A sky130_fd_sc_hd__fa_2_372/B sky130_fd_sc_hd__fa_2_372/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_13 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_4_1/Y
+ sky130_fd_sc_hd__dfxtp_1_138/CLK sky130_fd_sc_hd__o21ai_1_1/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_383 sky130_fd_sc_hd__fa_2_382/B sky130_fd_sc_hd__fa_2_384/A
+ sky130_fd_sc_hd__fa_2_383/A sky130_fd_sc_hd__fa_2_383/B sky130_fd_sc_hd__fa_2_383/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_24 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_2_60/A
+ sky130_fd_sc_hd__dfxtp_1_234/CLK sky130_fd_sc_hd__o21ai_2_3/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_394 sky130_fd_sc_hd__fah_1_16/B sky130_fd_sc_hd__fa_2_395/CIN
+ sky130_fd_sc_hd__fa_2_394/A sky130_fd_sc_hd__fa_2_394/B sky130_fd_sc_hd__fa_2_394/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_35 sky130_fd_sc_hd__conb_1_145/LO sky130_fd_sc_hd__clkinv_2_11/A
+ sky130_fd_sc_hd__dfxtp_1_343/CLK sky130_fd_sc_hd__nand4_1_1/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_46 sky130_fd_sc_hd__conb_1_145/LO sky130_fd_sc_hd__clkinv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_459/CLK sky130_fd_sc_hd__o31ai_2_0/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_104 sky130_fd_sc_hd__xor2_1_210/X sky130_fd_sc_hd__o21a_1_1/A2
+ sky130_fd_sc_hd__o21ai_1_32/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_115 sky130_fd_sc_hd__nor2_1_118/B sky130_fd_sc_hd__nor2_1_115/Y
+ sky130_fd_sc_hd__nor2_1_115/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_126 sky130_fd_sc_hd__nor2_1_126/B sky130_fd_sc_hd__nor2_1_126/Y
+ sky130_fd_sc_hd__nor2_1_126/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_13 sky130_fd_sc_hd__nor2_4_0/Y sky130_fd_sc_hd__nor2_2_0/Y
+ sky130_fd_sc_hd__dfxtp_1_334/Q sky130_fd_sc_hd__or2_0_90/A sky130_fd_sc_hd__nand2_2_3/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_137 sky130_fd_sc_hd__nor2_2_10/B sky130_fd_sc_hd__nor2_1_137/Y
+ sky130_fd_sc_hd__buf_6_4/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_148 sky130_fd_sc_hd__buf_6_1/X sky130_fd_sc_hd__nor2_1_148/Y
+ sky130_fd_sc_hd__buf_6_5/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_24 sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__dfxtp_1_279/Q sky130_fd_sc_hd__o211ai_1_3/Y sky130_fd_sc_hd__nand2_1_17/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_35 sky130_fd_sc_hd__clkbuf_1_24/X sky130_fd_sc_hd__clkbuf_1_23/X
+ sky130_fd_sc_hd__dfxtp_1_96/Q sky130_fd_sc_hd__dfxtp_1_64/Q sky130_fd_sc_hd__a22oi_1_35/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_159 sky130_fd_sc_hd__buf_4_7/X sky130_fd_sc_hd__nor2_1_159/Y
+ sky130_fd_sc_hd__buf_6_2/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_46 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__clkbuf_1_25/X
+ sky130_fd_sc_hd__nand2_1_76/B sky130_fd_sc_hd__dfxtp_1_134/Q sky130_fd_sc_hd__a22oi_1_46/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_57 sky130_fd_sc_hd__clkbuf_1_24/X sky130_fd_sc_hd__clkbuf_1_23/X
+ sky130_fd_sc_hd__dfxtp_1_107/Q sky130_fd_sc_hd__dfxtp_1_75/Q sky130_fd_sc_hd__a22oi_1_57/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_68 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__nor2_4_3/Y
+ sky130_fd_sc_hd__nand2_1_65/B sky130_fd_sc_hd__dfxtp_1_145/Q sky130_fd_sc_hd__a22oi_1_68/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_79 sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__dfxtp_1_118/Q sky130_fd_sc_hd__dfxtp_1_86/Q sky130_fd_sc_hd__a22oi_1_79/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_300 sky130_fd_sc_hd__buf_12_300/A sky130_fd_sc_hd__buf_12_300/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_311 sky130_fd_sc_hd__bufinv_8_2/Y sky130_fd_sc_hd__buf_12_526/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_322 sky130_fd_sc_hd__buf_12_322/A sky130_fd_sc_hd__buf_12_610/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_333 sky130_fd_sc_hd__buf_12_7/X sky130_fd_sc_hd__buf_12_623/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_344 sky130_fd_sc_hd__buf_12_344/A sky130_fd_sc_hd__buf_12_344/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_203 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__nor2b_1_8/Y sky130_fd_sc_hd__nor2_1_117/Y sky130_fd_sc_hd__a22oi_1_203/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_355 sky130_fd_sc_hd__buf_12_355/A sky130_fd_sc_hd__buf_12_658/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_214 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__buf_2_25/A
+ sky130_fd_sc_hd__nor2b_1_14/Y sky130_fd_sc_hd__nor2_1_174/Y sky130_fd_sc_hd__a22oi_1_214/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_366 sky130_fd_sc_hd__buf_12_73/X sky130_fd_sc_hd__buf_12_501/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_377 sky130_fd_sc_hd__buf_12_377/A sky130_fd_sc_hd__buf_12_489/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_388 sky130_fd_sc_hd__buf_12_388/A sky130_fd_sc_hd__buf_12_673/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_399 sky130_fd_sc_hd__buf_12_399/A sky130_fd_sc_hd__buf_12_502/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_500 sky130_fd_sc_hd__nand2_1_473/A sky130_fd_sc_hd__nor2_1_159/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_511 sky130_fd_sc_hd__or2b_2_1/A sky130_fd_sc_hd__dfxtp_1_218/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_522 sky130_fd_sc_hd__nor2_1_164/A sky130_fd_sc_hd__nand2_1_521/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_533 sky130_fd_sc_hd__nand2_1_527/A sky130_fd_sc_hd__nor2_2_21/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_544 sky130_fd_sc_hd__nand2_1_540/B sky130_fd_sc_hd__nor2_1_175/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_107 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_107/B sky130_fd_sc_hd__xnor2_1_107/Y
+ sky130_fd_sc_hd__xnor2_1_107/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_555 sky130_fd_sc_hd__o21ai_1_742/A2 sky130_fd_sc_hd__xnor2_1_150/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_118 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_2_5/Q sky130_fd_sc_hd__nor2_4_13/A
+ sky130_fd_sc_hd__xnor2_1_118/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_566 sky130_fd_sc_hd__o21ai_1_771/A2 sky130_fd_sc_hd__xnor2_1_156/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_129 vssd1 vccd1 sky130_fd_sc_hd__nand2_2_13/B sky130_fd_sc_hd__buf_2_13/A
+ sky130_fd_sc_hd__xnor2_1_129/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_577 sky130_fd_sc_hd__nand2_1_589/A sky130_fd_sc_hd__nor2_1_191/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_588 sky130_fd_sc_hd__o21ai_1_824/B1 sky130_fd_sc_hd__nand2_1_614/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_599 sky130_fd_sc_hd__clkinv_1_599/Y sky130_fd_sc_hd__nand2_1_637/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_4_13 sky130_fd_sc_hd__and2_4_0/B sky130_fd_sc_hd__clkinv_4_13/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_24 sky130_fd_sc_hd__clkinv_4_94/Y sky130_fd_sc_hd__clkinv_4_24/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_80 sky130_fd_sc_hd__nor2_1_80/B sky130_fd_sc_hd__nor2_1_80/Y
+ sky130_fd_sc_hd__nor2_1_80/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_35 sky130_fd_sc_hd__clkinv_8_69/A sky130_fd_sc_hd__clkinv_8_10/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_91 sky130_fd_sc_hd__nor2_1_91/B sky130_fd_sc_hd__nor2_1_91/Y
+ sky130_fd_sc_hd__nor2_1_91/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_46 sky130_fd_sc_hd__clkinv_4_46/A sky130_fd_sc_hd__clkinv_4_46/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_57 sky130_fd_sc_hd__clkinv_4_57/A sky130_fd_sc_hd__clkinv_4_57/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_68 sky130_fd_sc_hd__clkinv_4_68/A sky130_fd_sc_hd__clkinv_4_68/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_79 wbs_dat_i[27] sky130_fd_sc_hd__inv_2_196/A vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_1005 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1016 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1027 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1038 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1049 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21a_1_1 sky130_fd_sc_hd__o21a_1_1/X sky130_fd_sc_hd__o21a_1_1/A1
+ sky130_fd_sc_hd__o21a_1_1/B1 sky130_fd_sc_hd__o21a_1_1/A2 vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__decap_12_540 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_551 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_562 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_573 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_584 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_595 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_307 sky130_fd_sc_hd__fa_2_239/A sky130_fd_sc_hd__fa_2_211/B
+ sky130_fd_sc_hd__xor2_1_307/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_490 sky130_fd_sc_hd__xnor2_1_125/A sky130_fd_sc_hd__nand2_1_491/Y
+ sky130_fd_sc_hd__or2_0_51/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_318 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__fa_2_218/A
+ sky130_fd_sc_hd__xor2_1_318/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_329 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__fa_2_223/B
+ sky130_fd_sc_hd__xor2_1_329/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nor2b_1_70 sky130_fd_sc_hd__mux2_2_48/X sky130_fd_sc_hd__fa_2_486/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_81 sky130_fd_sc_hd__or2_0_82/B sky130_fd_sc_hd__nor2b_1_81/Y
+ sky130_fd_sc_hd__mux2_4_5/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_92 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_92/Y
+ sky130_fd_sc_hd__nor2b_1_92/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__xnor2_1_0 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_0/B sky130_fd_sc_hd__xnor2_1_0/Y
+ sky130_fd_sc_hd__xnor2_1_0/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_1070 sky130_fd_sc_hd__o21ai_1_912/B1 sky130_fd_sc_hd__o31ai_1_1/A1
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1081 sky130_fd_sc_hd__nand2_1_859/B sky130_fd_sc_hd__ha_2_47/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1092 sky130_fd_sc_hd__inv_2_71/A la_data_out[54] vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1550 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1561 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1572 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1583 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1594 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_15 sky130_fd_sc_hd__buf_8_98/A sky130_fd_sc_hd__dfxtp_1_9/CLK
+ sky130_fd_sc_hd__buf_2_193/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_26 sky130_fd_sc_hd__ha_2_7/A sky130_fd_sc_hd__dfxtp_1_29/CLK
+ sky130_fd_sc_hd__or4_1_3/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_180 sky130_fd_sc_hd__fa_2_174/CIN sky130_fd_sc_hd__fa_2_182/CIN
+ sky130_fd_sc_hd__fa_2_180/A sky130_fd_sc_hd__fa_2_180/B sky130_fd_sc_hd__xor2_1_267/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_37 sky130_fd_sc_hd__nand2_1_77/B sky130_fd_sc_hd__dfxtp_1_45/CLK
+ sky130_fd_sc_hd__dfxtp_1_37/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_191 sky130_fd_sc_hd__fa_2_178/A sky130_fd_sc_hd__fa_2_190/B
+ sky130_fd_sc_hd__fa_2_191/A sky130_fd_sc_hd__fa_2_191/B sky130_fd_sc_hd__xor2_1_280/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_48 sky130_fd_sc_hd__nand2_1_66/B sky130_fd_sc_hd__dfxtp_1_51/CLK
+ sky130_fd_sc_hd__dfxtp_1_48/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_59 sky130_fd_sc_hd__nand2_1_53/B sky130_fd_sc_hd__dfxtp_1_62/CLK
+ sky130_fd_sc_hd__dfxtp_1_59/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o22ai_1_90 sky130_fd_sc_hd__xnor2_1_247/Y sky130_fd_sc_hd__xnor2_1_238/Y
+ sky130_fd_sc_hd__fa_2_443/B sky130_fd_sc_hd__inv_2_65/Y sky130_fd_sc_hd__o22ai_1_99/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_309 vccd1 vssd1 sky130_fd_sc_hd__and2_0_309/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_309/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__inv_2_109 sky130_fd_sc_hd__inv_2_109/A sky130_fd_sc_hd__inv_2_160/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_sram_1kbyte_1rw1r_32x256_8_5 sky130_fd_sc_hd__clkinv_2_29/Y sky130_fd_sc_hd__clkinv_2_29/Y
+ sky130_fd_sc_hd__buf_12_660/X sky130_fd_sc_hd__buf_12_442/X sky130_fd_sc_hd__buf_12_604/X
+ sky130_fd_sc_hd__buf_12_502/X sky130_fd_sc_hd__buf_12_282/X sky130_fd_sc_hd__buf_12_643/X
+ sky130_fd_sc_hd__buf_12_635/X sky130_fd_sc_hd__nand2b_2_9/Y sky130_fd_sc_hd__buf_12_212/X
+ sky130_fd_sc_hd__buf_12_596/X sky130_fd_sc_hd__buf_12_611/X vccd1 sky130_fd_sc_hd__dfxtp_2_7/CLK
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[16] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[17]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[18] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[19]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[20] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[21]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[22] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[23]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[24] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[25]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[26] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[27]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[28] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[29]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[30] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[31]
+ sky130_fd_sc_hd__buf_12_541/X sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[1] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[2]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[3] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[4]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[5] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[6]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[7] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[8]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[9] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[10]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[11] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[12]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[13] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[14]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[15] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout1[0]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[10] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[11]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[12] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[13]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[14] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[15]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[16] sky130_fd_sc_hd__buf_12_518/X sky130_fd_sc_hd__buf_12_266/X
+ sky130_fd_sc_hd__buf_12_253/X sky130_fd_sc_hd__buf_12_292/X sky130_fd_sc_hd__buf_12_99/X
+ sky130_fd_sc_hd__clkinv_8_26/Y sky130_fd_sc_hd__buf_2_138/X sky130_fd_sc_hd__buf_2_138/X
+ sky130_fd_sc_hd__buf_2_138/X sky130_fd_sc_hd__buf_2_138/X sky130_fd_sc_hd__buf_2_138/X
+ sky130_fd_sc_hd__buf_2_138/X sky130_fd_sc_hd__buf_2_138/A sky130_fd_sc_hd__buf_2_138/A
+ sky130_fd_sc_hd__buf_2_138/A sky130_fd_sc_hd__buf_2_138/A sky130_fd_sc_hd__buf_2_138/A
+ sky130_fd_sc_hd__buf_2_138/A sky130_fd_sc_hd__buf_2_138/A sky130_fd_sc_hd__buf_2_139/X
+ sky130_fd_sc_hd__buf_2_139/X sky130_fd_sc_hd__buf_2_139/X sky130_fd_sc_hd__buf_2_139/X
+ sky130_fd_sc_hd__buf_2_139/X sky130_fd_sc_hd__buf_2_65/X sky130_fd_sc_hd__buf_2_65/X
+ sky130_fd_sc_hd__buf_2_65/X sky130_fd_sc_hd__buf_6_7/X sky130_fd_sc_hd__buf_6_7/X
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[0] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[1]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[2] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[3]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[4] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[5]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[6] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[7]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[8] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[9]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[25] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[26]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[27] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[28]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[29] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[30]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[31] sky130_fd_sc_hd__buf_6_7/X sky130_fd_sc_hd__buf_6_7/X
+ sky130_fd_sc_hd__buf_6_7/X sky130_fd_sc_hd__buf_6_7/X sky130_fd_sc_hd__buf_6_7/X
+ sky130_fd_sc_hd__buf_6_7/X sky130_fd_sc_hd__buf_6_7/X sky130_fd_sc_hd__buf_6_7/X
+ sky130_fd_sc_hd__buf_6_7/X sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[17] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[18]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[19] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[20]
+ sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[21] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[22]
+ sky130_fd_sc_hd__buf_12_551/X sky130_fd_sc_hd__buf_12_632/X sky130_fd_sc_hd__buf_12_654/X
+ sky130_fd_sc_hd__buf_12_495/X sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[23] sky130_sram_1kbyte_1rw1r_32x256_8_5/dout0[24]
+ vssd1 vssd1 sky130_sram_1kbyte_1rw1r_32x256_8
Xsky130_fd_sc_hd__buf_12_130 sky130_fd_sc_hd__buf_8_54/X sky130_fd_sc_hd__buf_12_408/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_141 sky130_fd_sc_hd__buf_12_11/X sky130_fd_sc_hd__buf_12_141/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_152 sky130_fd_sc_hd__buf_12_45/X sky130_fd_sc_hd__buf_12_423/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_163 sky130_fd_sc_hd__buf_12_38/X sky130_fd_sc_hd__buf_12_302/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_4_0 sky130_fd_sc_hd__and2_0_9/B sky130_fd_sc_hd__buf_2_16/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_12_174 sky130_fd_sc_hd__buf_8_96/X sky130_fd_sc_hd__buf_12_263/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_185 sky130_fd_sc_hd__buf_2_165/X sky130_fd_sc_hd__buf_12_347/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_196 sky130_fd_sc_hd__buf_4_35/X sky130_fd_sc_hd__buf_12_420/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_330 sky130_fd_sc_hd__nor2_1_53/A sky130_fd_sc_hd__nand2_1_200/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_341 sky130_fd_sc_hd__o21ai_1_251/A2 sky130_fd_sc_hd__xnor2_1_20/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_352 sky130_fd_sc_hd__nor2_1_66/B sky130_fd_sc_hd__nand2_1_226/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_363 sky130_fd_sc_hd__nand2_1_238/A sky130_fd_sc_hd__nor2_1_73/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_374 sky130_fd_sc_hd__xnor2_1_41/B sky130_fd_sc_hd__o21ai_2_7/A2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_385 sky130_fd_sc_hd__nand2_1_275/A sky130_fd_sc_hd__nor2_1_91/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_396 sky130_fd_sc_hd__nand2_1_302/A sky130_fd_sc_hd__nor2_1_44/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_2_4 sky130_fd_sc_hd__a21oi_2_4/B1 sky130_fd_sc_hd__or2_0_7/X
+ sky130_fd_sc_hd__o21ai_2_8/Y sky130_fd_sc_hd__a21oi_2_4/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_2
Xsky130_fd_sc_hd__clkinv_4_0 sky130_fd_sc_hd__clkinv_8_1/A sky130_fd_sc_hd__clkinv_4_0/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__conb_1_109 sky130_fd_sc_hd__conb_1_109/LO sky130_fd_sc_hd__conb_1_109/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_370 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_381 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_392 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_104 sky130_fd_sc_hd__fa_2_75/A sky130_fd_sc_hd__and3_4_5/A
+ sky130_fd_sc_hd__xor2_1_104/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_115 sky130_fd_sc_hd__fa_2_110/A sky130_fd_sc_hd__fa_2_85/A
+ sky130_fd_sc_hd__xor2_1_115/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_126 sky130_fd_sc_hd__fa_2_122/A sky130_fd_sc_hd__fa_2_95/B
+ sky130_fd_sc_hd__xor2_1_126/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_137 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__xor2_1_137/X
+ sky130_fd_sc_hd__xor2_1_137/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_148 sky130_fd_sc_hd__xor2_1_6/B sky130_fd_sc_hd__xor2_1_148/X
+ sky130_fd_sc_hd__xor2_1_148/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_159 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__fah_1_1/A
+ sky130_fd_sc_hd__xor2_1_159/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_108 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_3/A1 sky130_fd_sc_hd__clkbuf_1_108/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o21ai_1_800 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_2/Y sky130_fd_sc_hd__nand2b_1_16/Y
+ sky130_fd_sc_hd__o21ai_1_800/B1 sky130_fd_sc_hd__xor2_1_573/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1380 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_119 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_119/X sky130_fd_sc_hd__inv_4_6/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o21ai_1_811 vssd1 vccd1 sky130_fd_sc_hd__nor2_2_30/Y sky130_fd_sc_hd__nand2_1_613/Y
+ sky130_fd_sc_hd__nand2_1_608/Y sky130_fd_sc_hd__o21ai_1_811/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1391 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_822 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_861/A2 sky130_fd_sc_hd__nand2b_1_16/Y
+ sky130_fd_sc_hd__nand2_1_499/Y sky130_fd_sc_hd__xor2_1_595/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_833 vssd1 vccd1 sky130_fd_sc_hd__inv_2_52/Y sky130_fd_sc_hd__nor2_1_207/Y
+ sky130_fd_sc_hd__nand2_1_624/Y sky130_fd_sc_hd__xnor2_1_174/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_844 vssd1 vccd1 sky130_fd_sc_hd__buf_2_12/X sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_844/B1 sky130_fd_sc_hd__xor2_1_617/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_855 vssd1 vccd1 sky130_fd_sc_hd__nand2_2_13/Y sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__a22oi_1_223/Y sky130_fd_sc_hd__xor2_1_628/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_866 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_644/A sky130_fd_sc_hd__nor2_1_225/Y
+ sky130_fd_sc_hd__nand2_1_681/Y sky130_fd_sc_hd__xnor2_1_192/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_877 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_654/A sky130_fd_sc_hd__nor2_1_238/Y
+ sky130_fd_sc_hd__nand2_1_735/Y sky130_fd_sc_hd__xnor2_1_207/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_888 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_251/Y sky130_fd_sc_hd__nand2_1_781/Y
+ sky130_fd_sc_hd__nand2_1_780/Y sky130_fd_sc_hd__o21ai_1_888/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_899 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_682/A sky130_fd_sc_hd__nor2_1_260/Y
+ sky130_fd_sc_hd__nand2_1_817/Y sky130_fd_sc_hd__xnor2_1_296/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nand2b_2_1 sky130_fd_sc_hd__nor2_4_9/B sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__nor2_4_9/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_2
Xsky130_fd_sc_hd__xor2_1_660 sky130_fd_sc_hd__xor2_1_660/B sky130_fd_sc_hd__xor2_1_660/X
+ sky130_fd_sc_hd__xor2_1_660/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_671 sky130_fd_sc_hd__mux2_2_46/X sky130_fd_sc_hd__xor2_1_671/X
+ sky130_fd_sc_hd__or2_0_79/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_682 sky130_fd_sc_hd__xor2_1_682/B sky130_fd_sc_hd__xor2_1_682/X
+ sky130_fd_sc_hd__xor2_1_682/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_693 sky130_fd_sc_hd__ha_2_32/A sky130_fd_sc_hd__nand4_1_2/A
+ sky130_fd_sc_hd__ha_2_48/B vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__and2_0_106 vccd1 vssd1 sky130_fd_sc_hd__and2_0_106/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_106/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_14 la_data_out[113] sky130_fd_sc_hd__conb_1_128/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_117 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_34/D sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_117/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_25 la_data_out[102] sky130_fd_sc_hd__conb_1_117/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_128 vccd1 vssd1 sky130_fd_sc_hd__and2_0_128/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_128/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_36 la_data_out[27] sky130_fd_sc_hd__conb_1_106/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_139 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_70/D sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_139/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_47 la_data_out[16] sky130_fd_sc_hd__conb_1_95/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_58 la_data_out[5] sky130_fd_sc_hd__conb_1_84/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__fa_2_1 sky130_fd_sc_hd__xor3_1_1/C sky130_fd_sc_hd__fa_2_5/CIN sky130_fd_sc_hd__fa_2_1/A
+ sky130_fd_sc_hd__fa_2_1/B sky130_fd_sc_hd__fa_2_8/SUM vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_1_69 io_out[32] sky130_fd_sc_hd__conb_1_73/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_160 sky130_fd_sc_hd__o22ai_1_35/B1 sky130_fd_sc_hd__dfxtp_1_189/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_171 sky130_fd_sc_hd__o21ai_1_8/A2 sky130_fd_sc_hd__dfxtp_1_119/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_3 sky130_fd_sc_hd__buf_8_3/A sky130_fd_sc_hd__buf_8_3/X vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__a22o_1_5 sky130_fd_sc_hd__nand2_1_7/B sky130_fd_sc_hd__or2_0_77/B
+ sky130_fd_sc_hd__buf_6_4/A sky130_fd_sc_hd__or2_0_77/A sky130_fd_sc_hd__nand2_1_8/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_182 sky130_fd_sc_hd__nor2_1_25/A sky130_fd_sc_hd__dfxtp_1_148/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_193 sky130_fd_sc_hd__o22ai_1_46/B1 sky130_fd_sc_hd__dfxtp_1_176/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_40 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__buf_2_115/X
+ sky130_fd_sc_hd__a22o_1_40/X sky130_fd_sc_hd__a22o_1_40/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_51 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__buf_2_125/X
+ sky130_fd_sc_hd__a22o_1_51/X sky130_fd_sc_hd__a22o_1_51/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_62 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__buf_6_6/A
+ sky130_fd_sc_hd__a22o_1_62/X sky130_fd_sc_hd__a22o_1_62/B2 sky130_fd_sc_hd__a22o_1_71/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_73 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__buf_2_181/X
+ sky130_fd_sc_hd__a22o_1_73/X sky130_fd_sc_hd__ha_2_19/SUM sky130_fd_sc_hd__nor2_1_269/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__nand4_1_1 sky130_fd_sc_hd__nand4_1_1/C sky130_fd_sc_hd__nand4_1_1/B
+ sky130_fd_sc_hd__nand4_1_1/Y sky130_fd_sc_hd__nor3b_1_0/Y sky130_fd_sc_hd__nand4_1_1/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__o21ai_1_107 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_109/A2 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_121/Y sky130_fd_sc_hd__and2_0_169/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_118 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_121/A2 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_126/Y sky130_fd_sc_hd__and2_0_155/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_129 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_129/A2 sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__a22oi_1_175/Y sky130_fd_sc_hd__and2_0_142/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__inv_8_3 sky130_fd_sc_hd__inv_8_3/A la_data_out[93] vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__inv_8
Xsky130_fd_sc_hd__nand2_1_30 sky130_fd_sc_hd__nand2_2_8/A sky130_fd_sc_hd__nand2_1_7/B
+ sky130_fd_sc_hd__mux2_2_31/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_41 sky130_fd_sc_hd__nand2_1_41/Y sky130_fd_sc_hd__nand2_1_8/B
+ sky130_fd_sc_hd__xnor2_2_4/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_52 sky130_fd_sc_hd__nand2_1_52/Y sky130_fd_sc_hd__nand2_1_52/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_63 sky130_fd_sc_hd__nand2_1_63/Y sky130_fd_sc_hd__nand2_1_63/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_74 sky130_fd_sc_hd__nand2_1_74/Y sky130_fd_sc_hd__nand2_1_74/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_85 sky130_fd_sc_hd__nand2_1_85/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__xor2_2_1/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_290 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_290/B sky130_fd_sc_hd__xnor2_1_290/Y
+ sky130_fd_sc_hd__xnor2_1_290/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_96 sky130_fd_sc_hd__nand2_1_96/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__xor2_1_276/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_307 sky130_fd_sc_hd__dfxtp_1_307/Q sky130_fd_sc_hd__clkinv_8_6/Y
+ sky130_fd_sc_hd__and2_0_283/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_318 sky130_fd_sc_hd__nor2_1_238/A sky130_fd_sc_hd__dfxtp_1_323/CLK
+ sky130_fd_sc_hd__and2_0_295/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_329 sky130_fd_sc_hd__dfxtp_1_329/Q sky130_fd_sc_hd__dfxtp_1_343/CLK
+ sky130_fd_sc_hd__and2_0_318/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_630 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_447/A sky130_fd_sc_hd__nor2_2_22/Y
+ sky130_fd_sc_hd__nand2_1_517/B sky130_fd_sc_hd__xnor2_1_132/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_641 vssd1 vccd1 sky130_fd_sc_hd__inv_2_46/Y sky130_fd_sc_hd__nand2b_1_18/Y
+ sky130_fd_sc_hd__o21ai_1_641/B1 sky130_fd_sc_hd__xor2_1_429/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_652 vssd1 vccd1 sky130_fd_sc_hd__inv_2_51/Y sky130_fd_sc_hd__nand2b_1_15/Y
+ sky130_fd_sc_hd__o21ai_1_652/B1 sky130_fd_sc_hd__xor2_1_437/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_663 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_861/A2 sky130_fd_sc_hd__nand2b_1_17/Y
+ sky130_fd_sc_hd__nand2_1_492/Y sky130_fd_sc_hd__ha_2_2/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_674 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_126/Y sky130_fd_sc_hd__nand2b_1_16/Y
+ sky130_fd_sc_hd__o21ai_1_674/B1 sky130_fd_sc_hd__xor2_1_455/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_685 vssd1 vccd1 sky130_fd_sc_hd__nand2_2_13/Y sky130_fd_sc_hd__nand2b_1_18/Y
+ sky130_fd_sc_hd__a22oi_1_214/Y sky130_fd_sc_hd__xor2_1_464/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_696 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_861/A2 sky130_fd_sc_hd__nand2b_1_18/Y
+ sky130_fd_sc_hd__nand2_1_493/Y sky130_fd_sc_hd__xor2_1_474/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_15 sky130_fd_sc_hd__fa_2_0/B sky130_fd_sc_hd__fa_2_17/CIN sky130_fd_sc_hd__fa_2_15/A
+ sky130_fd_sc_hd__fa_2_15/B sky130_fd_sc_hd__fa_2_16/SUM vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_26 sky130_fd_sc_hd__fa_2_17/A sky130_fd_sc_hd__fa_2_26/SUM
+ sky130_fd_sc_hd__fa_2_26/A sky130_fd_sc_hd__fa_2_26/B sky130_fd_sc_hd__fa_2_26/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_37 sky130_fd_sc_hd__fa_2_30/CIN sky130_fd_sc_hd__fa_2_39/B
+ sky130_fd_sc_hd__fa_2_37/A sky130_fd_sc_hd__fa_2_37/B sky130_fd_sc_hd__xor2_1_58/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_48 sky130_fd_sc_hd__fa_2_42/CIN sky130_fd_sc_hd__fa_2_48/SUM
+ sky130_fd_sc_hd__fa_2_48/A sky130_fd_sc_hd__fa_2_48/B sky130_fd_sc_hd__xor2_1_66/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_59 sky130_fd_sc_hd__nor2_1_58/A sky130_fd_sc_hd__or2_0_3/B
+ sky130_fd_sc_hd__fa_2_59/A sky130_fd_sc_hd__fa_2_59/B sky130_fd_sc_hd__fa_2_59/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_207 vccd1 vssd1 sky130_fd_sc_hd__buf_2_207/X sky130_fd_sc_hd__or2_1_10/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__xor2_1_490 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__fa_2_328/B
+ sky130_fd_sc_hd__xor2_1_490/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a222oi_1_510 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__buf_2_4/A
+ sky130_fd_sc_hd__buf_2_20/X sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__buf_2_21/X
+ sky130_fd_sc_hd__o21ai_1_807/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_521 vccd1 vssd1 sky130_fd_sc_hd__and3_4_20/X sky130_fd_sc_hd__or2_0_72/A
+ sky130_fd_sc_hd__or2_0_71/B sky130_fd_sc_hd__nor2_4_16/Y sky130_fd_sc_hd__buf_2_29/X
+ sky130_fd_sc_hd__o21ai_1_821/B1 sky130_fd_sc_hd__and2b_4_11/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_532 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__buf_4_0/A
+ sky130_fd_sc_hd__buf_2_27/A sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__buf_2_31/X
+ sky130_fd_sc_hd__o21ai_1_840/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_543 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__or2_0_52/B
+ sky130_fd_sc_hd__or2_0_53/A sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__o21ai_1_859/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_554 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_416/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_448/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_751/A sky130_fd_sc_hd__dfxtp_1_384/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_565 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_405/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_437/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_762/A sky130_fd_sc_hd__dfxtp_1_373/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_576 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_404/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_436/Q sky130_fd_sc_hd__clkbuf_1_32/X
+ sky130_fd_sc_hd__clkinv_1_773/A sky130_fd_sc_hd__dfxtp_1_372/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_587 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_413/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_445/Q sky130_fd_sc_hd__clkbuf_1_32/X
+ sky130_fd_sc_hd__clkinv_1_784/A sky130_fd_sc_hd__dfxtp_1_381/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_598 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_416/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_448/Q sky130_fd_sc_hd__nor2_4_19/B
+ sky130_fd_sc_hd__clkinv_1_795/A sky130_fd_sc_hd__dfxtp_1_384/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nor2b_1_110 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_110/Y
+ sky130_fd_sc_hd__nor2b_1_110/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__decap_12_16 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_121 sky130_fd_sc_hd__nor3_1_2/Y sky130_fd_sc_hd__nor2b_1_121/Y
+ sky130_fd_sc_hd__ha_2_45/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__decap_12_27 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_132 sky130_fd_sc_hd__clkinv_4_51/Y sky130_fd_sc_hd__nor2b_1_132/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__decap_12_38 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_143 sky130_fd_sc_hd__clkinv_4_62/Y sky130_fd_sc_hd__nor2b_1_143/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__decap_12_49 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_154 sky130_fd_sc_hd__clkinv_4_73/Y sky130_fd_sc_hd__nor2b_1_154/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__fah_1_12 sky130_fd_sc_hd__fa_2_401/B sky130_fd_sc_hd__fah_1_12/B
+ sky130_fd_sc_hd__fah_1_12/A sky130_fd_sc_hd__fa_2_402/A sky130_fd_sc_hd__fah_1_12/CI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__fah_1
Xsky130_fd_sc_hd__buf_6_0 vccd1 vssd1 sky130_fd_sc_hd__buf_6_0/X sky130_fd_sc_hd__buf_6_0/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_16 vccd1 vssd1 sky130_fd_sc_hd__buf_6_16/X sky130_fd_sc_hd__buf_6_16/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_27 vccd1 vssd1 sky130_fd_sc_hd__buf_6_27/X sky130_fd_sc_hd__buf_8_86/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_38 vccd1 vssd1 sky130_fd_sc_hd__buf_6_90/A sky130_fd_sc_hd__buf_6_38/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_49 vccd1 vssd1 sky130_fd_sc_hd__buf_6_49/X sky130_fd_sc_hd__buf_8_89/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_18 sky130_fd_sc_hd__clkinv_4_69/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_29 sky130_fd_sc_hd__clkinv_4_59/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__inv_6_0 sky130_fd_sc_hd__inv_6_0/Y sky130_fd_sc_hd__inv_6_0/A vccd1
+ vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_6
Xsky130_fd_sc_hd__nand2_1_308 sky130_fd_sc_hd__xnor2_1_60/B sky130_fd_sc_hd__nand2_1_309/Y
+ sky130_fd_sc_hd__or2_0_21/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_907 sky130_fd_sc_hd__clkinv_1_907/Y sky130_fd_sc_hd__clkinv_1_907/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_1 sky130_fd_sc_hd__nor2_4_7/Y sky130_fd_sc_hd__nor2_1_1/Y
+ sky130_fd_sc_hd__nor2_4_1/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nand2_1_319 sky130_fd_sc_hd__xnor2_1_4/B sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_918 sky130_fd_sc_hd__clkinv_1_919/A sky130_fd_sc_hd__buf_2_51/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_929 sky130_fd_sc_hd__inv_2_118/A sky130_fd_sc_hd__buf_6_17/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_104 sky130_fd_sc_hd__dfxtp_1_104/Q sky130_fd_sc_hd__dfxtp_1_105/CLK
+ sky130_fd_sc_hd__and2_0_147/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_115 sky130_fd_sc_hd__dfxtp_1_115/Q sky130_fd_sc_hd__dfxtp_1_118/CLK
+ sky130_fd_sc_hd__and2_0_203/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_126 sky130_fd_sc_hd__dfxtp_1_126/Q sky130_fd_sc_hd__dfxtp_1_126/CLK
+ sky130_fd_sc_hd__and2_0_250/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_137 sky130_fd_sc_hd__dfxtp_1_137/Q sky130_fd_sc_hd__dfxtp_1_138/CLK
+ sky130_fd_sc_hd__and2_0_156/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_148 sky130_fd_sc_hd__dfxtp_1_148/Q sky130_fd_sc_hd__dfxtp_1_152/CLK
+ sky130_fd_sc_hd__and2_0_211/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_159 sky130_fd_sc_hd__dfxtp_1_159/Q sky130_fd_sc_hd__dfxtp_1_176/CLK
+ sky130_fd_sc_hd__and2_0_102/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_460 vssd1 vccd1 sky130_fd_sc_hd__inv_2_32/Y sky130_fd_sc_hd__nand2b_1_8/Y
+ sky130_fd_sc_hd__o21ai_1_460/B1 sky130_fd_sc_hd__xor2_1_263/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_471 vssd1 vccd1 sky130_fd_sc_hd__inv_2_37/Y sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_471/B1 sky130_fd_sc_hd__xor2_1_274/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_482 vssd1 vccd1 sky130_fd_sc_hd__inv_2_33/Y sky130_fd_sc_hd__nand2b_1_9/Y
+ sky130_fd_sc_hd__o21ai_1_482/B1 sky130_fd_sc_hd__xor2_1_283/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_493 vssd1 vccd1 sky130_fd_sc_hd__buf_2_11/X sky130_fd_sc_hd__nand2b_1_14/Y
+ sky130_fd_sc_hd__o21ai_1_493/B1 sky130_fd_sc_hd__xor2_1_294/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_903 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_914 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_925 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_936 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_820 sky130_fd_sc_hd__xor2_1_683/B sky130_fd_sc_hd__nand2_1_821/Y
+ sky130_fd_sc_hd__nand2_1_820/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_947 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_831 sky130_fd_sc_hd__nand2_1_831/Y sky130_fd_sc_hd__or2_0_109/A
+ sky130_fd_sc_hd__or2_0_109/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_958 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_842 sky130_fd_sc_hd__xnor2_1_303/B sky130_fd_sc_hd__nand2_1_843/Y
+ sky130_fd_sc_hd__or2_0_112/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_969 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_853 sky130_fd_sc_hd__nand2_1_853/Y sky130_fd_sc_hd__nand2_1_855/Y
+ sky130_fd_sc_hd__nand3_1_5/C vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_864 sky130_fd_sc_hd__nor4b_2_0/B sky130_fd_sc_hd__nor4_1_4/Y
+ sky130_fd_sc_hd__nor4_1_5/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o21ai_1_20 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_13/B1 sky130_fd_sc_hd__inv_2_53/A
+ sky130_fd_sc_hd__o21ai_1_20/B1 sky130_fd_sc_hd__fa_2_118/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_31 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_0/B1 sky130_fd_sc_hd__inv_2_53/A
+ sky130_fd_sc_hd__o21ai_1_31/B1 sky130_fd_sc_hd__or2_0_24/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_42 vssd1 vccd1 sky130_fd_sc_hd__inv_2_58/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_88/Y sky130_fd_sc_hd__and2_0_6/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_53 vssd1 vccd1 sky130_fd_sc_hd__inv_2_59/Y sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__o21ai_1_53/B1 sky130_fd_sc_hd__o21ai_1_53/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_64 vssd1 vccd1 sky130_fd_sc_hd__inv_2_55/Y sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_64/B1 sky130_fd_sc_hd__o21ai_1_64/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_75 vssd1 vccd1 sky130_fd_sc_hd__inv_2_61/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__o21ai_1_75/B1 sky130_fd_sc_hd__o21ai_1_75/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_86 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_89/A2 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__o21ai_1_86/B1 sky130_fd_sc_hd__o21ai_1_86/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_97 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_99/A2 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__o21ai_1_97/B1 sky130_fd_sc_hd__o21ai_1_97/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nand2_4_2 sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__ha_2_9/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_4
Xsky130_fd_sc_hd__a222oi_1_340 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__buf_6_1/X sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__and2_0_38/A
+ sky130_fd_sc_hd__o21ai_1_565/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_280 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_280/X sky130_fd_sc_hd__clkbuf_1_280/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_351 vccd1 vssd1 sky130_fd_sc_hd__and3_4_11/X sky130_fd_sc_hd__buf_4_7/X
+ sky130_fd_sc_hd__buf_4_0/X sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__buf_2_23/X
+ sky130_fd_sc_hd__o21ai_1_580/B1 sky130_fd_sc_hd__and2b_4_8/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_291 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_292/A sky130_fd_sc_hd__buf_8_59/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_362 vccd1 vssd1 sky130_fd_sc_hd__and3_4_11/X sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__buf_8_0/X sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__o21ai_1_597/B1 sky130_fd_sc_hd__and2b_4_8/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_373 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__buf_4_7/X sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__buf_4_0/X
+ sky130_fd_sc_hd__o21ai_1_617/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_384 vccd1 vssd1 sky130_fd_sc_hd__and3_4_26/X sky130_fd_sc_hd__nor2_2_10/B
+ sky130_fd_sc_hd__buf_6_4/X sky130_fd_sc_hd__nor2_2_31/Y sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__o21ai_1_645/B1 sky130_fd_sc_hd__nor2b_1_12/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_395 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__or2_0_58/A
+ sky130_fd_sc_hd__or2_0_9/B sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__or2_0_9/A
+ sky130_fd_sc_hd__o21ai_1_658/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__buf_12_504 sky130_fd_sc_hd__buf_12_504/A sky130_fd_sc_hd__buf_12_504/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_515 sky130_fd_sc_hd__buf_12_515/A sky130_fd_sc_hd__buf_12_676/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_526 sky130_fd_sc_hd__buf_12_526/A sky130_fd_sc_hd__buf_12_526/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_537 sky130_fd_sc_hd__buf_12_537/A sky130_fd_sc_hd__buf_12_537/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_548 sky130_fd_sc_hd__buf_12_548/A sky130_fd_sc_hd__buf_12_548/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_559 sky130_fd_sc_hd__buf_12_559/A sky130_fd_sc_hd__buf_12_559/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__nand2_1_105 sky130_fd_sc_hd__o21ai_1_75/B1 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__xor2_1_313/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_704 sky130_fd_sc_hd__a221o_1_0/B2 sky130_fd_sc_hd__ha_2_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_116 sky130_fd_sc_hd__o21ai_1_96/B1 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__xor2_1_367/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_715 sky130_fd_sc_hd__nor2b_1_94/A sky130_fd_sc_hd__xor2_1_676/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_127 sky130_fd_sc_hd__nand2_1_127/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_127/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_726 sky130_fd_sc_hd__nor2b_1_105/A sky130_fd_sc_hd__xnor2_1_296/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_138 sky130_fd_sc_hd__nand2_1_138/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__xnor2_1_120/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_737 sky130_fd_sc_hd__nor2b_1_116/A sky130_fd_sc_hd__xor2_1_687/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_149 sky130_fd_sc_hd__inv_2_7/A sky130_fd_sc_hd__inv_2_54/Y
+ sky130_fd_sc_hd__nor2b_1_1/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_748 sky130_fd_sc_hd__fa_2_471/A sky130_fd_sc_hd__clkinv_1_748/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_759 sky130_fd_sc_hd__fa_2_482/A sky130_fd_sc_hd__clkinv_1_759/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__or2_0_102 sky130_fd_sc_hd__or2_0_102/A sky130_fd_sc_hd__or2_0_102/X
+ sky130_fd_sc_hd__or2_0_102/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_113 sky130_fd_sc_hd__or2_0_113/A sky130_fd_sc_hd__or2_0_113/X
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__decap_12_1209 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_9 sky130_fd_sc_hd__xor2_1_9/B sky130_fd_sc_hd__xor3_1_9/B
+ sky130_fd_sc_hd__xor2_1_9/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkinv_8_7 sky130_fd_sc_hd__clkinv_8_7/Y sky130_fd_sc_hd__clkinv_8_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__o21ai_1_290 vssd1 vccd1 sky130_fd_sc_hd__inv_2_18/Y sky130_fd_sc_hd__nand2b_1_1/Y
+ sky130_fd_sc_hd__o21ai_1_290/B1 sky130_fd_sc_hd__xor2_1_111/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_700 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_711 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_722 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_733 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_744 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_755 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_766 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_650 sky130_fd_sc_hd__xnor2_1_185/B sky130_fd_sc_hd__nand2_1_651/Y
+ sky130_fd_sc_hd__or2_0_67/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_777 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_661 sky130_fd_sc_hd__nand2_1_661/Y sky130_fd_sc_hd__or2_0_70/A
+ sky130_fd_sc_hd__or2_0_70/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_788 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_672 sky130_fd_sc_hd__xor2_1_642/B sky130_fd_sc_hd__nand2_1_673/Y
+ sky130_fd_sc_hd__nand2_1_672/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_799 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_683 sky130_fd_sc_hd__nand2_1_683/Y sky130_fd_sc_hd__or2_0_77/A
+ sky130_fd_sc_hd__or2_0_77/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_694 sky130_fd_sc_hd__xnor2_1_196/A sky130_fd_sc_hd__nand2_1_695/Y
+ sky130_fd_sc_hd__or2_0_80/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_1710 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1721 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_20 sky130_fd_sc_hd__inv_2_20/A sky130_fd_sc_hd__inv_2_20/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1732 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_31 sky130_fd_sc_hd__inv_2_31/A sky130_fd_sc_hd__inv_2_31/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1743 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_42 sky130_fd_sc_hd__inv_2_42/A sky130_fd_sc_hd__inv_2_42/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1754 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_53 sky130_fd_sc_hd__inv_2_53/A sky130_fd_sc_hd__inv_2_53/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1765 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_64 sky130_fd_sc_hd__inv_2_64/A sky130_fd_sc_hd__inv_6_0/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1776 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_75 sky130_fd_sc_hd__inv_2_77/A sky130_fd_sc_hd__inv_2_75/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1787 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_86 sky130_fd_sc_hd__inv_2_86/A sky130_fd_sc_hd__inv_2_86/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_490 la_data_out[39] sky130_fd_sc_hd__dfxtp_1_498/CLK sky130_fd_sc_hd__and2_0_364/X
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1798 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_97 sky130_fd_sc_hd__inv_4_16/Y sky130_fd_sc_hd__inv_2_97/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__ha_2_18 vssd1 vccd1 sky130_fd_sc_hd__ha_2_18/A sky130_fd_sc_hd__or2_0_111/A
+ sky130_fd_sc_hd__ha_2_18/SUM sky130_fd_sc_hd__ha_2_18/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__a222oi_1_170 vccd1 vssd1 sky130_fd_sc_hd__and3_4_8/X sky130_fd_sc_hd__buf_2_32/X
+ sky130_fd_sc_hd__buf_8_0/X sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__o21ai_1_321/B1 sky130_fd_sc_hd__nor2b_2_2/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__ha_2_29 vssd1 vccd1 la_data_out[43] sky130_fd_sc_hd__ha_2_28/B sky130_fd_sc_hd__ha_2_29/SUM
+ sky130_fd_sc_hd__ha_2_29/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__a222oi_1_181 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__nor2_1_85/B sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__nor2_2_10/B
+ sky130_fd_sc_hd__o21ai_1_165/B1 sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_192 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__buf_2_4/A
+ sky130_fd_sc_hd__buf_6_5/X sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__o21ai_1_355/B1 sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_340 sky130_fd_sc_hd__fa_2_332/A sky130_fd_sc_hd__fa_2_339/B
+ sky130_fd_sc_hd__fa_2_340/A sky130_fd_sc_hd__fa_2_340/B sky130_fd_sc_hd__fa_2_340/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_351 sky130_fd_sc_hd__fa_2_344/A sky130_fd_sc_hd__fa_2_350/B
+ sky130_fd_sc_hd__fa_2_351/A sky130_fd_sc_hd__fa_2_351/B sky130_fd_sc_hd__xor2_1_519/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_362 sky130_fd_sc_hd__or2_1_5/A sky130_fd_sc_hd__nor2_2_26/B
+ sky130_fd_sc_hd__fa_2_362/A sky130_fd_sc_hd__fa_2_362/B sky130_fd_sc_hd__fa_2_362/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_373 sky130_fd_sc_hd__fa_2_363/A sky130_fd_sc_hd__fa_2_369/B
+ sky130_fd_sc_hd__fa_2_373/A sky130_fd_sc_hd__fa_2_373/B sky130_fd_sc_hd__xor2_1_547/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_14 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_4_3/Y
+ sky130_fd_sc_hd__dfxtp_1_146/CLK sky130_fd_sc_hd__o21ai_1_1/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_384 sky130_fd_sc_hd__fa_2_381/A sky130_fd_sc_hd__fa_2_385/B
+ sky130_fd_sc_hd__fa_2_384/A sky130_fd_sc_hd__fa_2_384/B sky130_fd_sc_hd__xor2_1_566/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_25 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_2_60/A
+ sky130_fd_sc_hd__dfxtp_2_5/CLK sky130_fd_sc_hd__o21ai_2_3/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_395 sky130_fd_sc_hd__or2_1_1/A sky130_fd_sc_hd__nor2_2_29/B
+ sky130_fd_sc_hd__fa_2_395/A sky130_fd_sc_hd__fa_2_395/B sky130_fd_sc_hd__fa_2_395/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_36 sky130_fd_sc_hd__conb_1_145/LO sky130_fd_sc_hd__clkinv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_395/CLK sky130_fd_sc_hd__o21ai_1_892/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_47 sky130_fd_sc_hd__conb_1_148/LO sky130_fd_sc_hd__clkinv_2_48/Y
+ sky130_fd_sc_hd__dfxtp_1_515/CLK sky130_fd_sc_hd__nor2_1_267/B vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_105 sky130_fd_sc_hd__nor2_2_18/Y sky130_fd_sc_hd__nor2_1_105/Y
+ sky130_fd_sc_hd__nor2_1_150/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_116 sky130_fd_sc_hd__or2_0_42/B sky130_fd_sc_hd__nor2_1_116/Y
+ sky130_fd_sc_hd__or2_0_39/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_127 sky130_fd_sc_hd__and3_4_14/A sky130_fd_sc_hd__nor2_1_127/Y
+ sky130_fd_sc_hd__and3_4_14/C vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_138 sky130_fd_sc_hd__nor2_1_139/Y sky130_fd_sc_hd__nor2_1_138/Y
+ sky130_fd_sc_hd__nor2_1_142/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_14 sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__dfxtp_1_284/Q sky130_fd_sc_hd__o211ai_1_8/Y sky130_fd_sc_hd__nand2_1_13/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_149 sky130_fd_sc_hd__nor2_1_149/B sky130_fd_sc_hd__nor2_1_149/Y
+ sky130_fd_sc_hd__nor2_1_149/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_25 sky130_fd_sc_hd__nor2_4_0/Y sky130_fd_sc_hd__nor2_2_0/Y
+ sky130_fd_sc_hd__dfxtp_1_328/Q sky130_fd_sc_hd__or2_0_92/A sky130_fd_sc_hd__nand2_1_17/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_36 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__clkbuf_1_25/X
+ sky130_fd_sc_hd__nand2_1_83/B sky130_fd_sc_hd__dfxtp_1_129/Q sky130_fd_sc_hd__a22oi_1_36/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_47 sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__dfxtp_1_102/Q sky130_fd_sc_hd__dfxtp_1_70/Q sky130_fd_sc_hd__a22oi_1_47/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_58 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__clkbuf_1_25/X
+ sky130_fd_sc_hd__nand2_1_70/B sky130_fd_sc_hd__dfxtp_1_140/Q sky130_fd_sc_hd__a22oi_1_58/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_69 sky130_fd_sc_hd__clkbuf_1_24/X sky130_fd_sc_hd__clkbuf_1_23/X
+ sky130_fd_sc_hd__dfxtp_1_113/Q sky130_fd_sc_hd__dfxtp_1_81/Q sky130_fd_sc_hd__a22oi_1_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_301 sky130_fd_sc_hd__buf_12_301/A sky130_fd_sc_hd__buf_12_547/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_312 sky130_fd_sc_hd__buf_12_94/X sky130_fd_sc_hd__buf_12_479/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_323 sky130_fd_sc_hd__buf_12_39/X sky130_fd_sc_hd__buf_12_631/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_334 sky130_fd_sc_hd__buf_12_2/X sky130_fd_sc_hd__buf_12_602/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_345 sky130_fd_sc_hd__buf_12_345/A sky130_fd_sc_hd__buf_12_579/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_204 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__nor2b_1_9/Y sky130_fd_sc_hd__nor2_1_121/Y sky130_fd_sc_hd__a22oi_1_204/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_356 sky130_fd_sc_hd__buf_12_356/A sky130_fd_sc_hd__buf_12_649/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_215 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__buf_2_25/A
+ sky130_fd_sc_hd__nor2b_1_15/Y sky130_fd_sc_hd__nor2_1_178/Y sky130_fd_sc_hd__a22oi_1_215/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_367 sky130_fd_sc_hd__buf_12_51/X sky130_fd_sc_hd__buf_12_647/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_378 sky130_fd_sc_hd__buf_12_378/A sky130_fd_sc_hd__buf_12_378/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_389 sky130_fd_sc_hd__buf_12_389/A sky130_fd_sc_hd__buf_12_531/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_501 sky130_fd_sc_hd__a21oi_1_99/A2 sky130_fd_sc_hd__nand2_1_476/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_512 sky130_fd_sc_hd__nand2_1_597/A sky130_fd_sc_hd__nor2_2_29/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_523 sky130_fd_sc_hd__clkinv_1_523/Y sky130_fd_sc_hd__nor2_1_168/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_534 sky130_fd_sc_hd__o21ai_1_691/A2 sky130_fd_sc_hd__xnor2_1_139/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_545 sky130_fd_sc_hd__nand2_1_542/A sky130_fd_sc_hd__nor2_1_177/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_108 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_108/B sky130_fd_sc_hd__inv_2_32/A
+ sky130_fd_sc_hd__xnor2_1_108/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_556 sky130_fd_sc_hd__nor2_1_179/A sky130_fd_sc_hd__nand2_1_564/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_119 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_119/B sky130_fd_sc_hd__inv_2_29/A
+ sky130_fd_sc_hd__xnor2_1_119/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_567 sky130_fd_sc_hd__o21ai_1_772/B1 sky130_fd_sc_hd__nand2_1_572/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_578 sky130_fd_sc_hd__nand2_1_595/A sky130_fd_sc_hd__nor2_1_193/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_589 sky130_fd_sc_hd__o21ai_1_824/A1 sky130_fd_sc_hd__nor2_1_201/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_4_14 sky130_fd_sc_hd__clkinv_4_14/A sky130_fd_sc_hd__nand2b_1_31/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_70 sky130_fd_sc_hd__nor2_1_73/Y sky130_fd_sc_hd__nor2_1_70/Y
+ sky130_fd_sc_hd__nor2_1_71/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_25 sky130_fd_sc_hd__clkinv_4_95/Y sky130_fd_sc_hd__clkinv_4_25/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_81 sky130_fd_sc_hd__nor2_2_10/B sky130_fd_sc_hd__nor2_1_81/Y
+ sky130_fd_sc_hd__nor2_1_85/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_36 sky130_fd_sc_hd__clkinv_8_12/Y sky130_fd_sc_hd__clkinv_8_13/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_92 sky130_fd_sc_hd__buf_2_4/X sky130_fd_sc_hd__nor2_1_92/Y
+ sky130_fd_sc_hd__buf_6_5/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_47 sky130_fd_sc_hd__clkinv_4_47/A sky130_fd_sc_hd__clkinv_4_47/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_58 sky130_fd_sc_hd__clkinv_4_58/A sky130_fd_sc_hd__clkinv_4_58/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_69 sky130_fd_sc_hd__clkinv_4_69/A sky130_fd_sc_hd__clkinv_4_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_1006 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1017 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1028 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1039 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21a_1_2 sky130_fd_sc_hd__o21a_1_2/X sky130_fd_sc_hd__or2_0_32/A
+ sky130_fd_sc_hd__o21a_1_2/B1 sky130_fd_sc_hd__o21a_1_2/A2 vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__decap_12_530 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_541 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_552 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_563 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_574 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_585 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_596 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_480 sky130_fd_sc_hd__nand2_1_480/Y sky130_fd_sc_hd__or2_0_48/A
+ sky130_fd_sc_hd__or2_0_48/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_308 sky130_fd_sc_hd__fa_2_217/A sky130_fd_sc_hd__fa_2_214/B
+ sky130_fd_sc_hd__xor2_1_308/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_491 sky130_fd_sc_hd__nand2_1_491/Y sky130_fd_sc_hd__or2_0_51/A
+ sky130_fd_sc_hd__or2_0_51/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_319 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__xor2_1_319/X
+ sky130_fd_sc_hd__xor2_1_319/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nor2b_1_60 sky130_fd_sc_hd__or2_0_78/A sky130_fd_sc_hd__fa_2_481/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_71 sky130_fd_sc_hd__mux2_4_2/X sky130_fd_sc_hd__nor2b_1_71/Y
+ sky130_fd_sc_hd__mux2_4_5/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_82 sky130_fd_sc_hd__mux2_4_4/X sky130_fd_sc_hd__fa_2_492/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_93 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_93/Y
+ sky130_fd_sc_hd__nor2b_1_93/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1060 sky130_fd_sc_hd__inv_16_3/A sky130_fd_sc_hd__buf_8_73/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_1 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_1/B sky130_fd_sc_hd__buf_2_5/A
+ sky130_fd_sc_hd__xnor2_1_1/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_1071 sky130_fd_sc_hd__a221oi_1_3/B2 sky130_fd_sc_hd__a21o_2_0/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1082 sky130_fd_sc_hd__o21ai_1_918/A2 sky130_fd_sc_hd__ha_2_52/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1540 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1093 sky130_fd_sc_hd__a22o_1_78/A2 sky130_fd_sc_hd__clkinv_4_84/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1551 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1562 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1573 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1584 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1595 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_16 sky130_fd_sc_hd__buf_2_193/A sky130_fd_sc_hd__dfxtp_1_8/CLK
+ la_data_out[58] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_170 sky130_fd_sc_hd__fa_2_161/CIN sky130_fd_sc_hd__fa_2_172/A
+ sky130_fd_sc_hd__fa_2_170/A sky130_fd_sc_hd__fa_2_170/B sky130_fd_sc_hd__xor2_1_261/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_27 sky130_fd_sc_hd__ha_2_8/A sky130_fd_sc_hd__dfxtp_1_29/CLK
+ sky130_fd_sc_hd__ha_2_45/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_181 sky130_fd_sc_hd__fa_2_174/A sky130_fd_sc_hd__fa_2_182/B
+ sky130_fd_sc_hd__fa_2_181/A sky130_fd_sc_hd__fa_2_181/B sky130_fd_sc_hd__xor2_1_270/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_38 sky130_fd_sc_hd__nand2_1_76/B sky130_fd_sc_hd__dfxtp_1_45/CLK
+ sky130_fd_sc_hd__dfxtp_1_38/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_192 sky130_fd_sc_hd__fa_2_184/A sky130_fd_sc_hd__fa_2_186/A
+ sky130_fd_sc_hd__fa_2_192/A sky130_fd_sc_hd__fa_2_192/B sky130_fd_sc_hd__xor2_1_284/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_49 sky130_fd_sc_hd__nand2_1_65/B sky130_fd_sc_hd__dfxtp_1_51/CLK
+ sky130_fd_sc_hd__dfxtp_1_49/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o22ai_1_80 sky130_fd_sc_hd__xnor2_2_4/Y sky130_fd_sc_hd__xnor2_1_239/Y
+ sky130_fd_sc_hd__fa_2_441/B sky130_fd_sc_hd__xnor2_1_230/Y sky130_fd_sc_hd__o22ai_1_96/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_91 sky130_fd_sc_hd__xnor2_2_4/Y sky130_fd_sc_hd__xnor2_1_244/Y
+ sky130_fd_sc_hd__o22ai_1_91/Y sky130_fd_sc_hd__xnor2_1_239/Y sky130_fd_sc_hd__o22ai_1_96/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_sram_1kbyte_1rw1r_32x256_8_6 sky130_fd_sc_hd__buf_2_157/X sky130_fd_sc_hd__buf_2_157/X
+ sky130_fd_sc_hd__buf_12_594/X sky130_fd_sc_hd__buf_12_637/X sky130_fd_sc_hd__buf_12_625/X
+ sky130_fd_sc_hd__buf_12_600/X sky130_fd_sc_hd__buf_12_571/X sky130_fd_sc_hd__buf_12_647/X
+ sky130_fd_sc_hd__buf_12_623/X sky130_fd_sc_hd__clkinv_4_21/Y sky130_fd_sc_hd__buf_12_679/X
+ sky130_fd_sc_hd__buf_12_545/X sky130_fd_sc_hd__buf_12_565/X vccd1 sky130_fd_sc_hd__clkinv_8_18/Y
+ sky130_fd_sc_hd__clkbuf_1_229/A sky130_fd_sc_hd__clkbuf_1_147/A sky130_fd_sc_hd__clkbuf_1_233/A
+ sky130_fd_sc_hd__clkbuf_1_101/A sky130_fd_sc_hd__clkbuf_1_100/A sky130_fd_sc_hd__clkbuf_1_99/A
+ sky130_fd_sc_hd__clkbuf_1_98/A sky130_fd_sc_hd__clkbuf_1_97/A sky130_fd_sc_hd__clkbuf_1_96/A
+ sky130_fd_sc_hd__clkbuf_1_95/A sky130_fd_sc_hd__clkbuf_1_94/A sky130_fd_sc_hd__clkbuf_1_93/A
+ sky130_fd_sc_hd__clkbuf_1_92/A sky130_fd_sc_hd__clkbuf_1_91/A sky130_fd_sc_hd__clkbuf_1_90/A
+ sky130_fd_sc_hd__clkbuf_1_89/A sky130_fd_sc_hd__buf_12_570/X sky130_fd_sc_hd__clkbuf_1_108/A
+ sky130_fd_sc_hd__mux2_4_4/A1 sky130_fd_sc_hd__clkbuf_1_107/A sky130_fd_sc_hd__clkbuf_1_106/A
+ sky130_fd_sc_hd__clkbuf_1_105/A sky130_fd_sc_hd__clkbuf_1_104/A sky130_fd_sc_hd__clkbuf_1_226/A
+ sky130_fd_sc_hd__clkbuf_1_103/A sky130_fd_sc_hd__clkbuf_1_102/A sky130_fd_sc_hd__clkbuf_1_155/A
+ sky130_fd_sc_hd__clkbuf_1_154/A sky130_fd_sc_hd__clkbuf_1_152/A sky130_fd_sc_hd__clkbuf_1_151/A
+ sky130_fd_sc_hd__clkbuf_1_150/A sky130_fd_sc_hd__clkbuf_1_149/A sky130_fd_sc_hd__clkbuf_1_222/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[10] sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[11]
+ sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[12] sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[13]
+ sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[14] sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[15]
+ sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[16] sky130_fd_sc_hd__buf_12_563/X sky130_fd_sc_hd__conb_1_147/HI
+ sky130_fd_sc_hd__conb_1_147/HI sky130_fd_sc_hd__conb_1_147/HI sky130_fd_sc_hd__conb_1_147/HI
+ sky130_fd_sc_hd__clkinv_8_68/Y sky130_fd_sc_hd__clkinv_1_919/Y sky130_fd_sc_hd__clkbuf_1_320/X
+ sky130_fd_sc_hd__clkinv_1_1017/Y sky130_fd_sc_hd__clkbuf_1_313/X sky130_fd_sc_hd__clkinv_2_18/Y
+ sky130_fd_sc_hd__clkinv_1_909/Y sky130_fd_sc_hd__clkbuf_1_220/X sky130_fd_sc_hd__clkbuf_1_136/X
+ sky130_fd_sc_hd__clkbuf_1_321/X sky130_fd_sc_hd__clkinv_1_897/Y sky130_fd_sc_hd__clkinv_1_894/Y
+ sky130_fd_sc_hd__clkbuf_4_11/X sky130_fd_sc_hd__buf_2_158/X sky130_fd_sc_hd__buf_2_43/X
+ sky130_fd_sc_hd__buf_2_41/X sky130_fd_sc_hd__clkbuf_4_10/X sky130_fd_sc_hd__clkbuf_4_8/X
+ sky130_fd_sc_hd__clkbuf_4_7/X sky130_fd_sc_hd__buf_2_40/X sky130_fd_sc_hd__clkbuf_1_165/X
+ sky130_fd_sc_hd__buf_4_39/X sky130_fd_sc_hd__clkbuf_1_39/X sky130_fd_sc_hd__clkbuf_1_140/X
+ sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[0] sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[1]
+ sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[2] sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[3]
+ sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[4] sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[5]
+ sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[6] sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[7]
+ sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[8] sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[9]
+ sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[25] sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[26]
+ sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[27] sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[28]
+ sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[29] sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[30]
+ sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[31] sky130_fd_sc_hd__clkinv_1_848/Y sky130_fd_sc_hd__buf_4_38/X
+ sky130_fd_sc_hd__buf_2_183/X sky130_fd_sc_hd__buf_6_92/X sky130_fd_sc_hd__buf_2_182/X
+ sky130_fd_sc_hd__buf_2_181/X sky130_fd_sc_hd__buf_2_180/X sky130_fd_sc_hd__clkinv_1_856/Y
+ sky130_fd_sc_hd__clkbuf_1_36/X sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[17] sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[18]
+ sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[19] sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[20]
+ sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[21] sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[22]
+ sky130_fd_sc_hd__buf_12_564/X sky130_fd_sc_hd__buf_12_538/X sky130_fd_sc_hd__buf_12_651/X
+ sky130_fd_sc_hd__buf_12_558/X sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[23] sky130_sram_1kbyte_1rw1r_32x256_8_6/dout0[24]
+ vssd1 vssd1 sky130_sram_1kbyte_1rw1r_32x256_8
Xsky130_fd_sc_hd__buf_12_120 sky130_fd_sc_hd__buf_8_41/X sky130_fd_sc_hd__buf_12_433/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_131 sky130_fd_sc_hd__buf_8_37/X sky130_fd_sc_hd__buf_12_291/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_142 sky130_fd_sc_hd__buf_8_149/X sky130_fd_sc_hd__buf_12_424/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_153 sky130_fd_sc_hd__buf_12_13/X sky130_fd_sc_hd__buf_12_293/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_164 sky130_fd_sc_hd__buf_12_21/X sky130_fd_sc_hd__buf_12_164/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_4_1 sky130_fd_sc_hd__and2_0_99/B sky130_fd_sc_hd__buf_2_16/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_12_175 sky130_fd_sc_hd__buf_8_111/X sky130_fd_sc_hd__buf_12_256/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_186 sky130_fd_sc_hd__buf_2_166/X sky130_fd_sc_hd__buf_12_346/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_197 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__buf_12_197/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_320 sky130_fd_sc_hd__o21ai_1_199/A2 sky130_fd_sc_hd__xnor2_1_9/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_331 sky130_fd_sc_hd__nand2_1_188/A sky130_fd_sc_hd__nor2_1_55/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_342 sky130_fd_sc_hd__nor2_1_59/A sky130_fd_sc_hd__nand2_1_211/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_353 sky130_fd_sc_hd__o21ai_1_280/A1 sky130_fd_sc_hd__nor2_1_67/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_364 sky130_fd_sc_hd__a21oi_2_6/B1 sky130_fd_sc_hd__nand2_1_244/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_375 sky130_fd_sc_hd__nand2_1_259/A sky130_fd_sc_hd__nor2_1_83/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_386 sky130_fd_sc_hd__nand2_1_279/A sky130_fd_sc_hd__nor2_1_94/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_397 sky130_fd_sc_hd__a21oi_1_66/B1 sky130_fd_sc_hd__nand2_1_305/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_2_5 sky130_fd_sc_hd__a21oi_2_5/B1 sky130_fd_sc_hd__or2_0_8/X
+ sky130_fd_sc_hd__xnor2_1_32/B sky130_fd_sc_hd__a21oi_2_5/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_2
Xsky130_fd_sc_hd__clkinv_4_1 sky130_fd_sc_hd__clkinv_8_1/A sky130_fd_sc_hd__clkinv_4_1/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor4b_1_0 sky130_fd_sc_hd__nor4b_1_0/C sky130_fd_sc_hd__nor4b_1_0/B
+ sky130_fd_sc_hd__nor4b_1_0/A sky130_fd_sc_hd__nor4b_1_0/D_N sky130_fd_sc_hd__nor4b_1_0/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor4b_1
Xsky130_fd_sc_hd__decap_12_360 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_371 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_382 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_393 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_105 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__fa_2_76/A
+ sky130_fd_sc_hd__xor2_1_105/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_116 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__fa_2_81/B
+ sky130_fd_sc_hd__xor2_1_116/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_127 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__fa_2_95/A
+ sky130_fd_sc_hd__xor2_1_127/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_138 sky130_fd_sc_hd__fa_2_110/A sky130_fd_sc_hd__xor2_1_138/X
+ sky130_fd_sc_hd__xor2_1_138/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_149 sky130_fd_sc_hd__fa_2_110/A sky130_fd_sc_hd__nor2_2_7/B
+ sky130_fd_sc_hd__xor2_1_149/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1370 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_109 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_110/A sky130_fd_sc_hd__nand2b_2_9/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o21ai_1_801 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_861/A2 sky130_fd_sc_hd__nand2b_1_15/Y
+ sky130_fd_sc_hd__nand2_1_497/Y sky130_fd_sc_hd__xor2_1_574/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1381 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_812 vssd1 vccd1 sky130_fd_sc_hd__inv_2_52/Y sky130_fd_sc_hd__nor2_1_188/B
+ sky130_fd_sc_hd__a21oi_1_127/Y sky130_fd_sc_hd__xnor2_1_167/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1392 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_823 vssd1 vccd1 sky130_fd_sc_hd__inv_2_43/Y sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_823/B1 sky130_fd_sc_hd__xor2_1_598/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_834 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_206/Y sky130_fd_sc_hd__nand2_1_628/Y
+ sky130_fd_sc_hd__nand2_1_622/Y sky130_fd_sc_hd__o21ai_1_834/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_845 vssd1 vccd1 sky130_fd_sc_hd__inv_2_46/Y sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_845/B1 sky130_fd_sc_hd__xor2_1_618/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_856 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_2/Y sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_856/B1 sky130_fd_sc_hd__xor2_1_629/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_867 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_645/A sky130_fd_sc_hd__nor2_1_226/Y
+ sky130_fd_sc_hd__nand2_1_685/Y sky130_fd_sc_hd__xnor2_1_193/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_878 vssd1 vccd1 sky130_fd_sc_hd__nand2_1_736/Y sky130_fd_sc_hd__a21oi_1_156/Y
+ sky130_fd_sc_hd__a21oi_1_154/Y sky130_fd_sc_hd__o21ai_1_878/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_889 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_665/B sky130_fd_sc_hd__nor2_1_249/Y
+ sky130_fd_sc_hd__nand2_1_782/Y sky130_fd_sc_hd__o21ai_1_889/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nand2b_2_2 sky130_fd_sc_hd__and3_4_3/A sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__and3_4_3/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_2
Xsky130_fd_sc_hd__xor2_1_650 sky130_fd_sc_hd__xor2_1_650/B sky130_fd_sc_hd__xor2_1_650/X
+ sky130_fd_sc_hd__xor2_1_650/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_661 sky130_fd_sc_hd__xor2_1_661/B sky130_fd_sc_hd__or2_0_87/B
+ sky130_fd_sc_hd__xor2_1_661/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_672 sky130_fd_sc_hd__mux2_2_47/X sky130_fd_sc_hd__xor2_1_672/X
+ sky130_fd_sc_hd__or2_0_77/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_683 sky130_fd_sc_hd__xor2_1_683/B sky130_fd_sc_hd__xor2_1_683/X
+ sky130_fd_sc_hd__xor2_1_683/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_694 sky130_fd_sc_hd__ha_2_50/SUM sky130_fd_sc_hd__xor2_1_694/X
+ la_data_out[44] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__and2_0_107 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_96/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_107/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_15 la_data_out[112] sky130_fd_sc_hd__conb_1_127/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_118 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_98/D sky130_fd_sc_hd__o21ai_2_0/B1
+ sky130_fd_sc_hd__and2_0_118/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_26 la_data_out[101] sky130_fd_sc_hd__conb_1_116/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_129 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_68/D sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_129/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_37 la_data_out[26] sky130_fd_sc_hd__conb_1_105/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_48 la_data_out[15] sky130_fd_sc_hd__conb_1_94/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_59 la_data_out[4] sky130_fd_sc_hd__conb_1_83/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__fa_2_2 sky130_fd_sc_hd__xor3_1_2/C sky130_fd_sc_hd__fa_2_4/CIN sky130_fd_sc_hd__fa_2_2/A
+ sky130_fd_sc_hd__fa_2_2/B sky130_fd_sc_hd__fa_2_2/CIN vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a211o_1_30 vssd1 vccd1 sky130_fd_sc_hd__ha_2_1/B sky130_fd_sc_hd__dfxtp_1_93/Q
+ sky130_fd_sc_hd__nor2_1_34/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_30/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__clkinv_1_150 sky130_fd_sc_hd__nand2_2_11/A sky130_fd_sc_hd__ha_2_9/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_161 sky130_fd_sc_hd__nor2_1_34/A sky130_fd_sc_hd__dfxtp_1_157/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_172 sky130_fd_sc_hd__o22ai_1_39/B1 sky130_fd_sc_hd__dfxtp_1_190/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_4 sky130_fd_sc_hd__buf_8_4/A sky130_fd_sc_hd__buf_8_4/X vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__a22o_1_6 sky130_fd_sc_hd__inv_2_66/Y sky130_fd_sc_hd__or2_0_85/B
+ sky130_fd_sc_hd__a22o_1_6/X sky130_fd_sc_hd__a22o_1_9/B2 sky130_fd_sc_hd__a22o_1_6/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_183 sky130_fd_sc_hd__o22ai_1_21/B1 sky130_fd_sc_hd__dfxtp_1_116/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_194 sky130_fd_sc_hd__nor2_1_21/A sky130_fd_sc_hd__dfxtp_1_144/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_30 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__buf_2_105/X
+ sky130_fd_sc_hd__a22o_1_30/X sky130_fd_sc_hd__a22o_1_30/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_41 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__buf_2_116/X
+ sky130_fd_sc_hd__a22o_1_41/X sky130_fd_sc_hd__a22o_1_41/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_52 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__buf_2_126/X
+ sky130_fd_sc_hd__a22o_1_52/X sky130_fd_sc_hd__a22o_1_52/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_63 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__buf_2_184/X
+ sky130_fd_sc_hd__a22o_1_63/X sky130_fd_sc_hd__xor2_1_691/X sky130_fd_sc_hd__a22o_1_71/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_74 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__buf_2_182/X
+ sky130_fd_sc_hd__a22o_1_74/X sky130_fd_sc_hd__ha_2_20/SUM sky130_fd_sc_hd__nor2_1_269/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__nand4_1_2 sky130_fd_sc_hd__nand4_1_2/C sky130_fd_sc_hd__nand4_1_2/B
+ sky130_fd_sc_hd__nor3_1_3/C sky130_fd_sc_hd__nand4_1_2/D sky130_fd_sc_hd__nand4_1_2/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__o21ai_1_108 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_109/A2 sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__a22oi_1_164/Y sky130_fd_sc_hd__and2_0_167/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_119 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_121/A2 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_127/Y sky130_fd_sc_hd__and2_0_154/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_190 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_20 sky130_fd_sc_hd__nand2_8_1/B sky130_fd_sc_hd__nand2_1_8/B
+ sky130_fd_sc_hd__mux2_2_47/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_31 sky130_fd_sc_hd__nand2_8_4/B sky130_fd_sc_hd__nand2_1_8/B
+ sky130_fd_sc_hd__or2_0_80/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_42 sky130_fd_sc_hd__nand2_1_42/Y sky130_fd_sc_hd__nand2_1_7/B
+ sky130_fd_sc_hd__buf_4_41/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_53 sky130_fd_sc_hd__nand2_1_53/Y sky130_fd_sc_hd__nand2_1_53/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_64 sky130_fd_sc_hd__nand2_1_64/Y sky130_fd_sc_hd__nand2_1_64/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_75 sky130_fd_sc_hd__nand2_1_75/Y sky130_fd_sc_hd__nand2_1_75/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_280 vssd1 vccd1 sky130_fd_sc_hd__buf_4_41/X sky130_fd_sc_hd__xnor2_1_280/Y
+ sky130_fd_sc_hd__or2_0_79/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_86 sky130_fd_sc_hd__nand2_1_86/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__xnor2_2_1/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_291 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_291/B sky130_fd_sc_hd__xnor2_1_291/Y
+ sky130_fd_sc_hd__xnor2_1_291/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_97 sky130_fd_sc_hd__nand2_1_97/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__xor2_1_276/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_308 sky130_fd_sc_hd__or2_0_85/A sky130_fd_sc_hd__dfxtp_1_323/CLK
+ sky130_fd_sc_hd__and2_0_285/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_319 sky130_fd_sc_hd__nor2_1_237/A sky130_fd_sc_hd__dfxtp_1_319/CLK
+ sky130_fd_sc_hd__and2_0_296/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_620 vssd1 vccd1 sky130_fd_sc_hd__inv_2_29/Y sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_620/B1 sky130_fd_sc_hd__xor2_1_413/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_631 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_509/A sky130_fd_sc_hd__nor2_2_23/Y
+ sky130_fd_sc_hd__nand2_1_550/Y sky130_fd_sc_hd__xnor2_1_145/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_642 vssd1 vccd1 sky130_fd_sc_hd__nand2_2_13/Y sky130_fd_sc_hd__nand2b_1_17/Y
+ sky130_fd_sc_hd__a22oi_1_213/Y sky130_fd_sc_hd__xor3_1_25/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_653 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_9/X sky130_fd_sc_hd__nand2b_1_19/Y
+ sky130_fd_sc_hd__o21ai_1_653/B1 sky130_fd_sc_hd__xor2_1_438/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_664 vssd1 vccd1 sky130_fd_sc_hd__inv_2_45/Y sky130_fd_sc_hd__nand2b_1_21/Y
+ sky130_fd_sc_hd__o21ai_1_664/B1 sky130_fd_sc_hd__xor2_1_446/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_675 vssd1 vccd1 sky130_fd_sc_hd__inv_2_49/Y sky130_fd_sc_hd__nand2b_1_20/Y
+ sky130_fd_sc_hd__o21ai_1_675/B1 sky130_fd_sc_hd__xor2_1_456/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_686 vssd1 vccd1 sky130_fd_sc_hd__inv_2_50/Y sky130_fd_sc_hd__nand2b_1_16/Y
+ sky130_fd_sc_hd__o21ai_1_686/B1 sky130_fd_sc_hd__xor2_1_465/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_697 vssd1 vccd1 sky130_fd_sc_hd__inv_2_45/Y sky130_fd_sc_hd__nand2b_1_15/Y
+ sky130_fd_sc_hd__o21ai_1_697/B1 sky130_fd_sc_hd__xor2_1_476/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_16 sky130_fd_sc_hd__fa_2_0/A sky130_fd_sc_hd__fa_2_16/SUM sky130_fd_sc_hd__fa_2_16/A
+ sky130_fd_sc_hd__fa_2_16/B sky130_fd_sc_hd__fa_2_16/CIN vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_27 sky130_fd_sc_hd__fa_2_26/CIN sky130_fd_sc_hd__fa_2_34/B
+ sky130_fd_sc_hd__fa_2_27/A sky130_fd_sc_hd__fa_2_27/B sky130_fd_sc_hd__xor2_1_43/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_38 sky130_fd_sc_hd__fa_2_32/CIN sky130_fd_sc_hd__fa_2_40/CIN
+ sky130_fd_sc_hd__fa_2_38/A sky130_fd_sc_hd__fa_2_38/B sky130_fd_sc_hd__xor2_1_54/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_49 sky130_fd_sc_hd__fa_2_36/A sky130_fd_sc_hd__fa_2_48/B sky130_fd_sc_hd__fa_2_49/A
+ sky130_fd_sc_hd__fa_2_49/B sky130_fd_sc_hd__xor2_1_67/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_208 vccd1 vssd1 la_data_out[73] sky130_fd_sc_hd__or2_1_10/B
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__xor2_1_480 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__xor2_1_480/X
+ sky130_fd_sc_hd__xor2_1_480/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_491 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__fa_2_328/A
+ sky130_fd_sc_hd__xor2_1_491/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a222oi_1_500 vccd1 vssd1 sky130_fd_sc_hd__and3_4_18/X sky130_fd_sc_hd__or2_0_71/B
+ sky130_fd_sc_hd__buf_2_29/X sky130_fd_sc_hd__nor2_2_32/Y sky130_fd_sc_hd__buf_2_30/X
+ sky130_fd_sc_hd__o21ai_1_793/B1 sky130_fd_sc_hd__nor2b_2_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_511 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__nor2_1_85/B sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__nor2_2_10/B
+ sky130_fd_sc_hd__o21ai_1_636/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_522 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__buf_2_4/A
+ sky130_fd_sc_hd__buf_2_20/X sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__buf_2_21/X
+ sky130_fd_sc_hd__o21ai_1_823/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_533 vccd1 vssd1 sky130_fd_sc_hd__and3_4_21/X sky130_fd_sc_hd__buf_2_28/A
+ sky130_fd_sc_hd__or2_0_72/A sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__or2_0_71/B
+ sky130_fd_sc_hd__o21ai_1_842/B1 sky130_fd_sc_hd__and2b_4_12/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_544 vccd1 vssd1 sky130_fd_sc_hd__inv_2_68/Y sky130_fd_sc_hd__dfxtp_1_426/Q
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__ha_2_9/A sky130_fd_sc_hd__dfxtp_1_458/Q
+ sky130_fd_sc_hd__clkinv_1_741/A sky130_fd_sc_hd__dfxtp_1_394/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_555 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_415/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_447/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_752/A sky130_fd_sc_hd__dfxtp_1_383/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_566 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_404/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_436/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_763/A sky130_fd_sc_hd__dfxtp_1_372/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_577 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_403/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_435/Q sky130_fd_sc_hd__clkbuf_1_32/X
+ sky130_fd_sc_hd__clkinv_1_774/A sky130_fd_sc_hd__dfxtp_1_371/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_588 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_410/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_442/Q sky130_fd_sc_hd__clkbuf_1_32/X
+ sky130_fd_sc_hd__clkinv_1_785/A sky130_fd_sc_hd__dfxtp_1_378/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_599 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_417/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_449/Q sky130_fd_sc_hd__nor2_4_19/B
+ sky130_fd_sc_hd__clkinv_1_796/A sky130_fd_sc_hd__dfxtp_1_385/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nor2b_1_100 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_100/Y
+ sky130_fd_sc_hd__nor2b_1_100/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_111 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_111/Y
+ sky130_fd_sc_hd__nor2b_1_111/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__decap_12_17 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_122 sky130_fd_sc_hd__o31ai_1_0/Y sky130_fd_sc_hd__nor2b_1_122/Y
+ sky130_fd_sc_hd__and2_4_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__decap_12_28 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_133 sky130_fd_sc_hd__clkinv_4_52/Y sky130_fd_sc_hd__nor2b_1_133/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__decap_12_39 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_144 sky130_fd_sc_hd__clkinv_4_63/Y sky130_fd_sc_hd__nor2b_1_144/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_155 sky130_fd_sc_hd__clkinv_4_74/Y sky130_fd_sc_hd__nor2b_1_155/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__fah_1_13 sky130_fd_sc_hd__fa_2_393/B sky130_fd_sc_hd__fah_1_13/B
+ sky130_fd_sc_hd__fah_1_13/A sky130_fd_sc_hd__fa_2_396/A sky130_fd_sc_hd__fah_1_13/CI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__fah_1
Xsky130_fd_sc_hd__buf_6_1 vccd1 vssd1 sky130_fd_sc_hd__buf_6_1/X sky130_fd_sc_hd__buf_6_1/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_17 vccd1 vssd1 sky130_fd_sc_hd__buf_6_17/X sky130_fd_sc_hd__buf_6_17/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_28 vccd1 vssd1 sky130_fd_sc_hd__buf_6_28/X sky130_fd_sc_hd__buf_8_20/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_39 vccd1 vssd1 sky130_fd_sc_hd__buf_6_39/X sky130_fd_sc_hd__buf_8_68/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_19 sky130_fd_sc_hd__clkinv_4_65/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__inv_6_1 sky130_fd_sc_hd__inv_6_1/Y sky130_fd_sc_hd__inv_6_1/A vccd1
+ vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_6
Xsky130_fd_sc_hd__nand2_1_309 sky130_fd_sc_hd__nand2_1_309/Y sky130_fd_sc_hd__or2_0_21/A
+ sky130_fd_sc_hd__or2_0_21/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_908 sky130_fd_sc_hd__clkinv_1_909/A sky130_fd_sc_hd__buf_2_49/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_2 sky130_fd_sc_hd__nor2_1_2/B sky130_fd_sc_hd__nor2_1_2/Y
+ sky130_fd_sc_hd__nor2_1_2/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_1_919 sky130_fd_sc_hd__clkinv_1_919/Y sky130_fd_sc_hd__clkinv_1_919/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_105 sky130_fd_sc_hd__dfxtp_1_105/Q sky130_fd_sc_hd__dfxtp_1_105/CLK
+ sky130_fd_sc_hd__and2_0_153/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_116 sky130_fd_sc_hd__dfxtp_1_116/Q sky130_fd_sc_hd__dfxtp_1_118/CLK
+ sky130_fd_sc_hd__and2_0_208/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_127 sky130_fd_sc_hd__dfxtp_1_127/Q sky130_fd_sc_hd__dfxtp_1_146/CLK
+ sky130_fd_sc_hd__and2_0_106/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_138 sky130_fd_sc_hd__dfxtp_1_138/Q sky130_fd_sc_hd__dfxtp_1_138/CLK
+ sky130_fd_sc_hd__and2_0_161/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_149 sky130_fd_sc_hd__dfxtp_1_149/Q sky130_fd_sc_hd__dfxtp_1_152/CLK
+ sky130_fd_sc_hd__and2_0_216/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_450 vssd1 vccd1 sky130_fd_sc_hd__inv_2_33/Y sky130_fd_sc_hd__nand2b_1_8/Y
+ sky130_fd_sc_hd__o21ai_1_450/B1 sky130_fd_sc_hd__xor2_1_253/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_461 vssd1 vccd1 sky130_fd_sc_hd__inv_2_35/Y sky130_fd_sc_hd__nand2b_1_9/Y
+ sky130_fd_sc_hd__o21ai_1_461/B1 sky130_fd_sc_hd__xor2_1_264/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_472 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_472/A2 sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_472/B1 sky130_fd_sc_hd__xor2_1_275/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_483 vssd1 vccd1 sky130_fd_sc_hd__inv_2_31/Y sky130_fd_sc_hd__nand2b_1_8/Y
+ sky130_fd_sc_hd__o21ai_1_483/B1 sky130_fd_sc_hd__xor2_1_284/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_494 vssd1 vccd1 sky130_fd_sc_hd__buf_2_9/X sky130_fd_sc_hd__nand2b_1_8/Y
+ sky130_fd_sc_hd__o21ai_1_494/B1 sky130_fd_sc_hd__xor2_1_295/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_904 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_915 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_926 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_810 sky130_fd_sc_hd__xnor2_1_295/A sky130_fd_sc_hd__nand2_1_811/Y
+ sky130_fd_sc_hd__or2_0_104/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_937 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_821 sky130_fd_sc_hd__nand2_1_821/Y sky130_fd_sc_hd__nor2_1_261/A
+ sky130_fd_sc_hd__nor2_1_261/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_948 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_832 sky130_fd_sc_hd__xor2_1_686/B sky130_fd_sc_hd__nand2_1_833/Y
+ sky130_fd_sc_hd__nand2_1_832/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_959 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_843 sky130_fd_sc_hd__nand2_1_843/Y sky130_fd_sc_hd__or2_0_112/A
+ sky130_fd_sc_hd__or2_0_112/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_854 sky130_fd_sc_hd__nand2_1_854/Y sky130_fd_sc_hd__ha_2_46/A
+ sky130_fd_sc_hd__ha_2_46/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_865 sky130_fd_sc_hd__a21o_2_4/A2 sky130_fd_sc_hd__nand2_1_865/B
+ sky130_fd_sc_hd__a21o_2_3/B1 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o21ai_1_10 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_23/B1 sky130_fd_sc_hd__nor2_4_4/B
+ sky130_fd_sc_hd__o21ai_1_10/B1 sky130_fd_sc_hd__fa_2_64/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_21 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_12/B1 sky130_fd_sc_hd__nor2_4_4/B
+ sky130_fd_sc_hd__o21ai_1_21/B1 sky130_fd_sc_hd__fa_2_122/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_32 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_1/B1 sky130_fd_sc_hd__inv_2_53/A
+ sky130_fd_sc_hd__o21ai_1_32/B1 sky130_fd_sc_hd__o21ai_1_32/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_43 vssd1 vccd1 sky130_fd_sc_hd__inv_2_58/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_89/Y sky130_fd_sc_hd__and2_0_7/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_54 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_57/A2 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_94/Y sky130_fd_sc_hd__o21ai_1_54/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_65 vssd1 vccd1 sky130_fd_sc_hd__inv_2_55/Y sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__o21ai_1_65/B1 sky130_fd_sc_hd__o21ai_1_65/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_76 vssd1 vccd1 sky130_fd_sc_hd__inv_2_61/Y sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_76/B1 sky130_fd_sc_hd__o21ai_1_76/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_87 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_89/A2 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__o21ai_1_87/B1 sky130_fd_sc_hd__o21ai_1_87/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_98 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_98/A2 sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_98/B1 sky130_fd_sc_hd__o21ai_1_98/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nand2_4_3 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_40/A
+ sky130_fd_sc_hd__ha_2_9/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_4
Xsky130_fd_sc_hd__a222oi_1_330 vccd1 vssd1 sky130_fd_sc_hd__and3_4_11/X sky130_fd_sc_hd__buf_2_19/X
+ sky130_fd_sc_hd__buf_6_5/X sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__o21ai_1_551/B1 sky130_fd_sc_hd__and2b_4_8/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_270 vssd1 vccd1 sky130_fd_sc_hd__buf_8_113/A sky130_fd_sc_hd__inv_2_112/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_341 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__and2_0_49/A
+ sky130_fd_sc_hd__and2_0_45/A sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__and2_0_87/A
+ sky130_fd_sc_hd__o21ai_1_566/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_281 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_282/A sky130_fd_sc_hd__buf_8_57/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_352 vccd1 vssd1 sky130_fd_sc_hd__and3_4_10/X sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__buf_8_0/X sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__o21ai_1_581/B1 sky130_fd_sc_hd__and2b_4_7/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_292 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4_28/A sky130_fd_sc_hd__clkbuf_1_292/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_363 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__buf_2_31/X
+ sky130_fd_sc_hd__buf_2_19/X sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__o21ai_1_599/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_374 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__or2_0_52/B
+ sky130_fd_sc_hd__or2_0_53/A sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__o21ai_1_619/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_385 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__or2_0_61/B
+ sky130_fd_sc_hd__or2_0_58/B sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__or2_0_58/A
+ sky130_fd_sc_hd__o21ai_1_646/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_396 vccd1 vssd1 sky130_fd_sc_hd__and3_4_20/X sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__buf_4_4/X sky130_fd_sc_hd__nor2_4_16/Y sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__o21ai_1_661/B1 sky130_fd_sc_hd__and2b_4_11/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__and2_0_290 vccd1 vssd1 sky130_fd_sc_hd__and2_0_290/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_11/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_12_505 sky130_fd_sc_hd__buf_12_505/A sky130_fd_sc_hd__buf_12_611/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_516 sky130_fd_sc_hd__buf_12_516/A sky130_fd_sc_hd__buf_12_516/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_527 sky130_fd_sc_hd__buf_12_527/A sky130_fd_sc_hd__buf_12_527/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_538 sky130_fd_sc_hd__buf_12_538/A sky130_fd_sc_hd__buf_12_538/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_549 sky130_fd_sc_hd__buf_12_549/A sky130_fd_sc_hd__buf_12_549/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__nand2_1_106 sky130_fd_sc_hd__o21ai_1_78/B1 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__xnor2_1_91/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_705 sky130_fd_sc_hd__a221o_1_0/A1 sky130_fd_sc_hd__ha_2_4/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_117 sky130_fd_sc_hd__o21ai_1_97/B1 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__xor2_1_367/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_716 sky130_fd_sc_hd__nor2b_1_95/A sky130_fd_sc_hd__xnor2_1_291/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_128 sky130_fd_sc_hd__nand2_1_128/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_129/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_727 sky130_fd_sc_hd__nor2b_1_106/A sky130_fd_sc_hd__xor2_1_682/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_139 sky130_fd_sc_hd__nand2_1_139/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__xnor2_1_120/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_738 sky130_fd_sc_hd__nor2b_1_117/A sky130_fd_sc_hd__xnor2_1_302/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_749 sky130_fd_sc_hd__fa_2_472/A sky130_fd_sc_hd__clkinv_1_749/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__or2_0_103 sky130_fd_sc_hd__or2_0_103/A sky130_fd_sc_hd__or2_0_103/X
+ sky130_fd_sc_hd__or2_0_103/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__o21ai_1_280 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_2/X sky130_fd_sc_hd__o21ai_1_280/A1
+ sky130_fd_sc_hd__o21ai_1_280/B1 sky130_fd_sc_hd__xnor2_1_26/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkinv_8_8 sky130_fd_sc_hd__clkinv_8_8/Y wbs_dat_i[30] vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__o21ai_1_291 vssd1 vccd1 sky130_fd_sc_hd__inv_2_9/Y sky130_fd_sc_hd__nand2b_2_0/Y
+ sky130_fd_sc_hd__o21ai_1_291/B1 sky130_fd_sc_hd__xor2_1_112/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_701 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_712 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_723 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_734 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_745 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_756 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_640 sky130_fd_sc_hd__nand2_1_640/Y sky130_fd_sc_hd__or2_0_68/X
+ sky130_fd_sc_hd__or2_0_69/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_767 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_651 sky130_fd_sc_hd__nand2_1_651/Y sky130_fd_sc_hd__or2_0_67/A
+ sky130_fd_sc_hd__or2_0_67/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_778 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_662 sky130_fd_sc_hd__xnor2_1_188/A sky130_fd_sc_hd__nand2_1_663/Y
+ sky130_fd_sc_hd__or2_0_73/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_789 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_673 sky130_fd_sc_hd__nand2_1_673/Y sky130_fd_sc_hd__mux2_2_22/X
+ sky130_fd_sc_hd__mux2_2_42/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_684 sky130_fd_sc_hd__xor2_1_645/B sky130_fd_sc_hd__nand2_1_685/Y
+ sky130_fd_sc_hd__nand2_1_684/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_695 sky130_fd_sc_hd__nand2_1_695/Y sky130_fd_sc_hd__or2_0_80/A
+ sky130_fd_sc_hd__or2_0_80/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_1700 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1711 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_10 sky130_fd_sc_hd__inv_2_10/A sky130_fd_sc_hd__inv_2_10/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1722 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_21 sky130_fd_sc_hd__inv_2_21/A sky130_fd_sc_hd__inv_2_21/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1733 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_32 sky130_fd_sc_hd__inv_2_32/A sky130_fd_sc_hd__inv_2_32/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1744 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_43 sky130_fd_sc_hd__inv_2_43/A sky130_fd_sc_hd__inv_2_43/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1755 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_54 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__inv_2_54/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1766 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_65 sky130_fd_sc_hd__or2_0_84/B sky130_fd_sc_hd__inv_2_65/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1777 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_76 sky130_fd_sc_hd__inv_2_77/A sky130_fd_sc_hd__inv_2_76/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_480 sky130_fd_sc_hd__buf_2_175/A sky130_fd_sc_hd__dfxtp_1_480/CLK
+ sky130_fd_sc_hd__and2_0_388/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1788 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_2_0 sky130_fd_sc_hd__inv_4_8/A sky130_fd_sc_hd__nand2_2_0/A
+ sky130_fd_sc_hd__nand2_2_0/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__inv_2_87 la_data_out[41] sky130_fd_sc_hd__inv_2_89/A vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_491 sky130_fd_sc_hd__ha_2_32/A sky130_fd_sc_hd__dfxtp_1_498/CLK
+ sky130_fd_sc_hd__and2_0_369/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1799 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_98 sky130_fd_sc_hd__inv_4_17/Y sky130_fd_sc_hd__inv_2_98/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__a222oi_1_160 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__nor2_1_73/B sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__o21ai_1_308/B1 sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__ha_2_19 vssd1 vccd1 sky130_fd_sc_hd__ha_2_19/A sky130_fd_sc_hd__xor2_1_689/A
+ sky130_fd_sc_hd__ha_2_19/SUM sky130_fd_sc_hd__ha_2_19/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__a222oi_1_171 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__nor2_1_87/A sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__o21ai_1_323/B1 sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_182 vccd1 vssd1 sky130_fd_sc_hd__and3_4_8/X sky130_fd_sc_hd__or2_0_52/B
+ sky130_fd_sc_hd__or2_0_53/A sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__buf_2_32/X
+ sky130_fd_sc_hd__o21ai_1_339/B1 sky130_fd_sc_hd__nor2b_2_2/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_330 sky130_fd_sc_hd__fa_2_324/CIN sky130_fd_sc_hd__fa_2_330/SUM
+ sky130_fd_sc_hd__fa_2_330/A sky130_fd_sc_hd__fa_2_330/B sky130_fd_sc_hd__xor2_1_492/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_193 vccd1 vssd1 sky130_fd_sc_hd__and3_4_1/X sky130_fd_sc_hd__or2_0_52/B
+ sky130_fd_sc_hd__or2_0_53/A sky130_fd_sc_hd__nor2_2_9/Y sky130_fd_sc_hd__buf_2_32/X
+ sky130_fd_sc_hd__o21ai_1_357/B1 sky130_fd_sc_hd__and2b_4_3/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_341 sky130_fd_sc_hd__nor2_2_24/A sky130_fd_sc_hd__or2_1_6/B
+ sky130_fd_sc_hd__fa_2_341/A sky130_fd_sc_hd__fa_2_341/B sky130_fd_sc_hd__fa_2_341/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_352 sky130_fd_sc_hd__fa_2_348/B sky130_fd_sc_hd__fa_2_355/CIN
+ sky130_fd_sc_hd__fa_2_352/A sky130_fd_sc_hd__fa_2_352/B sky130_fd_sc_hd__fa_2_352/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_363 sky130_fd_sc_hd__fa_2_359/CIN sky130_fd_sc_hd__fa_2_368/A
+ sky130_fd_sc_hd__fa_2_363/A sky130_fd_sc_hd__fa_2_363/B sky130_fd_sc_hd__fa_2_367/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_374 sky130_fd_sc_hd__or2_1_4/A sky130_fd_sc_hd__nor2_2_25/B
+ sky130_fd_sc_hd__fa_2_374/A sky130_fd_sc_hd__fa_2_374/B sky130_fd_sc_hd__fa_2_374/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_15 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_4_0/Y
+ sky130_fd_sc_hd__dfxtp_1_190/CLK sky130_fd_sc_hd__o21ai_2_1/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_385 sky130_fd_sc_hd__fah_1_6/B sky130_fd_sc_hd__fa_2_387/CIN
+ sky130_fd_sc_hd__fa_2_385/A sky130_fd_sc_hd__fa_2_385/B sky130_fd_sc_hd__fa_2_385/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_26 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_8_4/Y
+ sky130_fd_sc_hd__dfxtp_1_275/CLK sky130_fd_sc_hd__o21ai_2_4/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_396 sky130_fd_sc_hd__fa_2_394/CIN sky130_fd_sc_hd__fah_1_9/A
+ sky130_fd_sc_hd__fa_2_396/A sky130_fd_sc_hd__fa_2_396/B sky130_fd_sc_hd__xor2_1_588/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_37 sky130_fd_sc_hd__conb_1_145/LO sky130_fd_sc_hd__clkinv_4_11/Y
+ sky130_fd_sc_hd__dfxtp_1_380/CLK sky130_fd_sc_hd__o21ai_1_892/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_48 sky130_fd_sc_hd__conb_1_148/LO sky130_fd_sc_hd__clkinv_2_48/Y
+ sky130_fd_sc_hd__dfxtp_1_520/CLK sky130_fd_sc_hd__nor2_1_267/B vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__clkinv_8_90 sky130_fd_sc_hd__clkinv_8_90/Y sky130_fd_sc_hd__clkinv_8_90/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__nor2_1_106 sky130_fd_sc_hd__nor2_1_106/B sky130_fd_sc_hd__nor2_1_106/Y
+ sky130_fd_sc_hd__nor2_1_106/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_117 sky130_fd_sc_hd__and3_1_1/B sky130_fd_sc_hd__nor2_1_117/Y
+ sky130_fd_sc_hd__and3_1_1/C vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_128 sky130_fd_sc_hd__nor2_1_131/Y sky130_fd_sc_hd__nor2_1_128/Y
+ sky130_fd_sc_hd__nor2_1_129/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_139 sky130_fd_sc_hd__nor2_1_139/B sky130_fd_sc_hd__nor2_1_139/Y
+ sky130_fd_sc_hd__nor2_1_139/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_15 sky130_fd_sc_hd__nor2_4_0/Y sky130_fd_sc_hd__nor2_2_0/Y
+ sky130_fd_sc_hd__dfxtp_1_333/Q sky130_fd_sc_hd__or2_0_89/A sky130_fd_sc_hd__nand2_1_13/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_26 sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__dfxtp_1_278/Q sky130_fd_sc_hd__o211ai_1_2/Y sky130_fd_sc_hd__nand2_2_5/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_37 sky130_fd_sc_hd__clkbuf_1_24/X sky130_fd_sc_hd__clkbuf_1_23/X
+ sky130_fd_sc_hd__dfxtp_1_97/Q sky130_fd_sc_hd__dfxtp_1_65/Q sky130_fd_sc_hd__a22oi_1_37/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_48 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__clkbuf_1_25/X
+ sky130_fd_sc_hd__nand2_1_75/B sky130_fd_sc_hd__dfxtp_1_135/Q sky130_fd_sc_hd__a22oi_1_48/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_59 sky130_fd_sc_hd__clkbuf_1_24/X sky130_fd_sc_hd__clkbuf_1_23/X
+ sky130_fd_sc_hd__dfxtp_1_108/Q sky130_fd_sc_hd__dfxtp_1_76/Q sky130_fd_sc_hd__a22oi_1_59/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_302 sky130_fd_sc_hd__buf_12_302/A sky130_fd_sc_hd__buf_12_569/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_313 sky130_fd_sc_hd__buf_12_313/A sky130_fd_sc_hd__buf_12_523/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_324 sky130_fd_sc_hd__buf_12_324/A sky130_fd_sc_hd__buf_12_609/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_335 sky130_fd_sc_hd__buf_12_335/A sky130_fd_sc_hd__buf_12_592/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_346 sky130_fd_sc_hd__buf_12_346/A sky130_fd_sc_hd__buf_12_586/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_205 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__nor2b_1_10/Y sky130_fd_sc_hd__nor2_1_127/Y sky130_fd_sc_hd__a22oi_1_205/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_357 sky130_fd_sc_hd__buf_12_357/A sky130_fd_sc_hd__buf_12_652/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_216 sky130_fd_sc_hd__or2_0_72/B sky130_fd_sc_hd__or2_0_72/A
+ sky130_fd_sc_hd__nor2b_1_16/Y sky130_fd_sc_hd__nor2_1_183/Y sky130_fd_sc_hd__a22oi_1_216/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_368 sky130_fd_sc_hd__buf_12_368/A sky130_fd_sc_hd__buf_12_482/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_379 sky130_fd_sc_hd__buf_12_35/X sky130_fd_sc_hd__buf_12_637/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_502 sky130_fd_sc_hd__xnor2_1_120/B sky130_fd_sc_hd__a21oi_1_102/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_513 sky130_fd_sc_hd__clkinv_1_513/Y sky130_fd_sc_hd__nand2_1_602/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_524 sky130_fd_sc_hd__nand2_1_514/A sky130_fd_sc_hd__nor2_1_169/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_535 sky130_fd_sc_hd__nor2_1_171/B sky130_fd_sc_hd__nand2_1_537/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_546 sky130_fd_sc_hd__a21oi_2_16/B1 sky130_fd_sc_hd__nand2_1_545/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_109 vssd1 vccd1 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__nor2_2_20/A
+ sky130_fd_sc_hd__xnor2_1_109/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_557 sky130_fd_sc_hd__nand2_1_560/A sky130_fd_sc_hd__nor2_2_26/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_568 sky130_fd_sc_hd__nor2_1_182/B sky130_fd_sc_hd__nor2_1_184/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_579 sky130_fd_sc_hd__clkinv_1_579/Y sky130_fd_sc_hd__nand2_1_606/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_60 sky130_fd_sc_hd__or2_0_61/A sky130_fd_sc_hd__nor2_1_60/Y
+ sky130_fd_sc_hd__or2_0_60/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_15 sky130_fd_sc_hd__clkinv_4_15/A sky130_fd_sc_hd__nand2_1_845/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_71 sky130_fd_sc_hd__nor2_1_73/B sky130_fd_sc_hd__nor2_1_71/Y
+ sky130_fd_sc_hd__buf_4_3/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_26 sky130_fd_sc_hd__nand2_2_5/Y sky130_fd_sc_hd__clkinv_4_26/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_82 sky130_fd_sc_hd__nor2_1_86/Y sky130_fd_sc_hd__nor2_1_82/Y
+ sky130_fd_sc_hd__nor2_1_88/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_37 sky130_fd_sc_hd__clkinv_8_14/Y sky130_fd_sc_hd__clkinv_4_37/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_93 sky130_fd_sc_hd__nor2_1_94/Y sky130_fd_sc_hd__nor2_1_93/Y
+ sky130_fd_sc_hd__nor2_1_97/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_48 sky130_fd_sc_hd__clkinv_4_48/A sky130_fd_sc_hd__clkinv_4_48/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_59 sky130_fd_sc_hd__clkinv_4_59/A sky130_fd_sc_hd__clkinv_4_59/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_1007 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1018 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1029 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21a_1_3 sky130_fd_sc_hd__o21a_1_3/X sky130_fd_sc_hd__o21a_1_3/A1
+ sky130_fd_sc_hd__o21a_1_3/B1 sky130_fd_sc_hd__o21a_1_3/A2 vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__decap_12_520 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_531 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_542 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_553 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_564 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_575 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_586 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_470 sky130_fd_sc_hd__xor2_1_411/B sky130_fd_sc_hd__nand2_1_471/Y
+ sky130_fd_sc_hd__or2_0_49/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_597 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_481 sky130_fd_sc_hd__xnor2_1_66/B sky130_fd_sc_hd__nand2_1_482/Y
+ sky130_fd_sc_hd__nand2_1_481/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_309 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__fa_2_210/A
+ sky130_fd_sc_hd__xor2_1_309/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_492 sky130_fd_sc_hd__nand2_1_492/Y sky130_fd_sc_hd__nor2_1_167/Y
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_50 sky130_fd_sc_hd__mux2_2_39/X sky130_fd_sc_hd__fa_2_476/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_61 sky130_fd_sc_hd__or2_0_78/B sky130_fd_sc_hd__nor2b_1_61/Y
+ sky130_fd_sc_hd__mux2_4_5/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_72 sky130_fd_sc_hd__or2_1_10/A sky130_fd_sc_hd__fa_2_487/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_83 la_data_out[68] sky130_fd_sc_hd__nor2b_1_83/Y sky130_fd_sc_hd__mux2_4_5/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1050 sky130_fd_sc_hd__inv_2_183/A sky130_fd_sc_hd__buf_6_20/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_94 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_94/Y
+ sky130_fd_sc_hd__nor2b_1_94/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1061 sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__buf_8_134/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_2 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_2/B sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__xnor2_1_2/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_1072 sky130_fd_sc_hd__o21ai_2_18/A1 sky130_fd_sc_hd__a21o_2_0/B1
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1530 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1083 sky130_fd_sc_hd__o21ai_1_915/A1 la_data_out[47] vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1541 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1094 sky130_fd_sc_hd__and2_0_356/A sky130_fd_sc_hd__clkinv_4_90/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1552 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1563 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1574 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1585 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1596 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__fa_2_160 sky130_fd_sc_hd__nor2_1_110/B sky130_fd_sc_hd__or2_0_28/B
+ sky130_fd_sc_hd__fa_2_160/A sky130_fd_sc_hd__fa_2_160/B sky130_fd_sc_hd__fa_2_167/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_17 sky130_fd_sc_hd__dfxtp_1_17/Q sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__dfxtp_1_17/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_171 sky130_fd_sc_hd__fa_2_166/CIN sky130_fd_sc_hd__fa_2_176/A
+ sky130_fd_sc_hd__fa_2_171/A sky130_fd_sc_hd__fa_2_171/B sky130_fd_sc_hd__xor2_1_259/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_28 sky130_fd_sc_hd__or4_1_1/B sky130_fd_sc_hd__edfxbp_1_0/CLK
+ sky130_fd_sc_hd__ha_2_46/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_182 sky130_fd_sc_hd__fa_2_175/A sky130_fd_sc_hd__fa_2_183/B
+ sky130_fd_sc_hd__fa_2_182/A sky130_fd_sc_hd__fa_2_182/B sky130_fd_sc_hd__fa_2_182/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_39 sky130_fd_sc_hd__nand2_1_75/B sky130_fd_sc_hd__dfxtp_1_45/CLK
+ sky130_fd_sc_hd__dfxtp_1_39/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_193 sky130_fd_sc_hd__or2_0_29/A sky130_fd_sc_hd__nor2_2_13/B
+ sky130_fd_sc_hd__fa_2_193/A sky130_fd_sc_hd__fa_2_193/B sky130_fd_sc_hd__fa_2_193/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o22ai_1_70 sky130_fd_sc_hd__xnor2_2_5/Y sky130_fd_sc_hd__xnor2_1_229/Y
+ sky130_fd_sc_hd__fa_2_431/B sky130_fd_sc_hd__xnor2_1_221/Y sky130_fd_sc_hd__o22ai_1_95/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_81 sky130_fd_sc_hd__xnor2_2_6/Y sky130_fd_sc_hd__xnor2_1_240/Y
+ sky130_fd_sc_hd__fa_2_441/A sky130_fd_sc_hd__xnor2_1_231/Y sky130_fd_sc_hd__o22ai_1_98/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_92 sky130_fd_sc_hd__xnor2_2_5/Y sky130_fd_sc_hd__o22ai_1_92/B1
+ sky130_fd_sc_hd__fa_2_442/B sky130_fd_sc_hd__o22ai_1_92/A1 sky130_fd_sc_hd__o22ai_1_95/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_12_110 sky130_fd_sc_hd__buf_8_140/X sky130_fd_sc_hd__buf_12_363/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_sram_1kbyte_1rw1r_32x256_8_7 sky130_fd_sc_hd__clkbuf_1_215/X sky130_fd_sc_hd__clkbuf_1_215/X
+ sky130_fd_sc_hd__buf_12_649/X sky130_fd_sc_hd__buf_12_531/X sky130_fd_sc_hd__buf_12_509/X
+ sky130_fd_sc_hd__buf_12_441/X sky130_fd_sc_hd__buf_12_653/X sky130_fd_sc_hd__buf_12_656/X
+ sky130_fd_sc_hd__buf_12_644/X sky130_fd_sc_hd__clkbuf_1_110/X sky130_fd_sc_hd__buf_12_610/X
+ sky130_fd_sc_hd__buf_12_207/X sky130_fd_sc_hd__buf_12_601/X vccd1 sky130_fd_sc_hd__clkinv_8_27/Y
+ sky130_fd_sc_hd__buf_2_96/A sky130_fd_sc_hd__buf_2_153/A sky130_fd_sc_hd__buf_2_95/A
+ sky130_fd_sc_hd__buf_2_94/A sky130_fd_sc_hd__buf_2_93/A sky130_fd_sc_hd__buf_2_92/A
+ sky130_fd_sc_hd__buf_2_91/A sky130_fd_sc_hd__buf_2_90/A sky130_fd_sc_hd__buf_2_89/A
+ sky130_fd_sc_hd__buf_2_88/A sky130_fd_sc_hd__buf_2_87/A sky130_fd_sc_hd__buf_2_86/A
+ sky130_fd_sc_hd__buf_2_85/A sky130_fd_sc_hd__buf_2_84/A sky130_fd_sc_hd__buf_2_83/A
+ sky130_fd_sc_hd__buf_6_22/A sky130_fd_sc_hd__buf_12_566/X sky130_fd_sc_hd__buf_4_24/A
+ sky130_fd_sc_hd__buf_4_25/A sky130_fd_sc_hd__buf_4_17/A sky130_fd_sc_hd__buf_4_13/A
+ sky130_fd_sc_hd__buf_2_147/A sky130_fd_sc_hd__buf_4_16/A sky130_fd_sc_hd__buf_4_18/A
+ sky130_fd_sc_hd__buf_4_15/A sky130_fd_sc_hd__buf_4_19/A sky130_fd_sc_hd__buf_2_150/A
+ sky130_fd_sc_hd__buf_4_21/A sky130_fd_sc_hd__buf_2_151/A sky130_fd_sc_hd__buf_2_148/A
+ sky130_fd_sc_hd__buf_2_149/A sky130_fd_sc_hd__buf_2_152/A sky130_fd_sc_hd__buf_4_11/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[10] sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[11]
+ sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[12] sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[13]
+ sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[14] sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[15]
+ sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[16] sky130_fd_sc_hd__buf_12_661/X sky130_fd_sc_hd__buf_12_300/X
+ sky130_fd_sc_hd__buf_12_112/X sky130_fd_sc_hd__buf_12_61/X sky130_fd_sc_hd__buf_12_200/X
+ sky130_fd_sc_hd__clkinv_8_24/Y sky130_fd_sc_hd__clkinv_1_1019/Y sky130_fd_sc_hd__clkinv_1_916/Y
+ sky130_fd_sc_hd__clkinv_2_19/Y sky130_fd_sc_hd__clkbuf_1_44/X sky130_fd_sc_hd__clkinv_1_911/Y
+ sky130_fd_sc_hd__buf_2_142/X sky130_fd_sc_hd__inv_2_104/Y sky130_fd_sc_hd__clkbuf_1_43/X
+ sky130_fd_sc_hd__clkbuf_1_316/X sky130_fd_sc_hd__inv_2_103/Y sky130_fd_sc_hd__clkinv_1_893/Y
+ sky130_fd_sc_hd__clkbuf_1_137/X sky130_fd_sc_hd__inv_2_101/Y sky130_fd_sc_hd__inv_2_100/Y
+ sky130_fd_sc_hd__inv_2_99/Y sky130_fd_sc_hd__inv_2_98/Y sky130_fd_sc_hd__clkbuf_1_218/X
+ sky130_fd_sc_hd__clkbuf_1_318/X sky130_fd_sc_hd__inv_2_97/Y sky130_fd_sc_hd__inv_2_96/Y
+ sky130_fd_sc_hd__clkbuf_1_317/X sky130_fd_sc_hd__clkbuf_1_38/X sky130_fd_sc_hd__clkbuf_1_37/X
+ sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[0] sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[1]
+ sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[2] sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[3]
+ sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[4] sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[5]
+ sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[6] sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[7]
+ sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[8] sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[9]
+ sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[25] sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[26]
+ sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[27] sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[28]
+ sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[29] sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[30]
+ sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[31] sky130_fd_sc_hd__buf_2_36/X sky130_fd_sc_hd__clkbuf_1_311/X
+ sky130_fd_sc_hd__clkbuf_1_141/X sky130_fd_sc_hd__clkinv_2_16/Y sky130_fd_sc_hd__clkbuf_1_219/X
+ sky130_fd_sc_hd__clkbuf_1_142/X sky130_fd_sc_hd__clkbuf_1_308/X sky130_fd_sc_hd__clkinv_1_854/Y
+ sky130_fd_sc_hd__clkinv_1_850/Y sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[17] sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[18]
+ sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[19] sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[20]
+ sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[21] sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[22]
+ sky130_fd_sc_hd__buf_12_523/X sky130_fd_sc_hd__buf_12_677/X sky130_fd_sc_hd__buf_12_533/X
+ sky130_fd_sc_hd__buf_12_628/X sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[23] sky130_sram_1kbyte_1rw1r_32x256_8_7/dout0[24]
+ vssd1 vssd1 sky130_sram_1kbyte_1rw1r_32x256_8
Xsky130_fd_sc_hd__buf_12_121 sky130_fd_sc_hd__buf_8_24/X sky130_fd_sc_hd__buf_12_121/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_132 sky130_fd_sc_hd__buf_8_35/X sky130_fd_sc_hd__buf_12_395/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_143 sky130_fd_sc_hd__buf_12_28/X sky130_fd_sc_hd__buf_12_378/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_154 sky130_fd_sc_hd__buf_12_23/X sky130_fd_sc_hd__buf_12_287/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_165 sky130_fd_sc_hd__buf_12_44/X sky130_fd_sc_hd__buf_12_284/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_4_2 sky130_fd_sc_hd__nor2_1_2/B sky130_fd_sc_hd__nor2_1_37/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_12_176 sky130_fd_sc_hd__buf_8_156/X sky130_fd_sc_hd__buf_12_264/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_187 sky130_fd_sc_hd__buf_2_159/X sky130_fd_sc_hd__buf_12_401/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_198 sky130_fd_sc_hd__buf_6_37/X sky130_fd_sc_hd__buf_12_446/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_310 sky130_fd_sc_hd__nand2_1_248/A sky130_fd_sc_hd__nor2_1_43/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_321 sky130_fd_sc_hd__nor2_1_49/B sky130_fd_sc_hd__nand2_1_183/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_332 sky130_fd_sc_hd__a21oi_2_1/B1 sky130_fd_sc_hd__nand2_1_191/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_343 sky130_fd_sc_hd__a21oi_1_45/A1 sky130_fd_sc_hd__o21a_1_0/A2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_354 sky130_fd_sc_hd__a21oi_2_4/B1 sky130_fd_sc_hd__nand2_1_223/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_365 sky130_fd_sc_hd__o21ai_1_327/A2 sky130_fd_sc_hd__nand2_1_250/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_376 sky130_fd_sc_hd__nand2_1_263/A sky130_fd_sc_hd__nor2_1_85/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_387 sky130_fd_sc_hd__nand2_1_281/A sky130_fd_sc_hd__nor2_1_95/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_398 sky130_fd_sc_hd__xnor2_1_57/B sky130_fd_sc_hd__a21oi_1_67/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_2_6 sky130_fd_sc_hd__a21oi_2_6/B1 sky130_fd_sc_hd__or2_0_11/X
+ sky130_fd_sc_hd__o21ai_2_7/Y sky130_fd_sc_hd__a21oi_2_6/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_2
Xsky130_fd_sc_hd__clkinv_4_2 sky130_fd_sc_hd__clkinv_4_2/A sky130_fd_sc_hd__clkinv_4_2/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__or2_0_90 sky130_fd_sc_hd__or2_0_90/A sky130_fd_sc_hd__or2_0_90/X
+ sky130_fd_sc_hd__or2_0_90/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__decap_12_350 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_361 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_372 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_383 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_394 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_106 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__fa_2_79/CIN
+ sky130_fd_sc_hd__xor2_1_106/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_117 sky130_fd_sc_hd__xor2_1_117/B sky130_fd_sc_hd__xor2_1_117/X
+ sky130_fd_sc_hd__a21oi_2_5/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_128 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__fa_2_93/CIN
+ sky130_fd_sc_hd__xor2_1_128/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_139 sky130_fd_sc_hd__fa_2_122/A sky130_fd_sc_hd__fa_2_100/A
+ sky130_fd_sc_hd__xor2_1_139/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1360 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1371 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_802 vssd1 vccd1 sky130_fd_sc_hd__inv_2_45/Y sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_802/B1 sky130_fd_sc_hd__xor2_1_576/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1382 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_813 vssd1 vccd1 sky130_fd_sc_hd__buf_2_12/X sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__o21ai_1_813/B1 sky130_fd_sc_hd__xor2_1_588/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1393 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_824 vssd1 vccd1 sky130_fd_sc_hd__inv_2_52/Y sky130_fd_sc_hd__o21ai_1_824/A1
+ sky130_fd_sc_hd__o21ai_1_824/B1 sky130_fd_sc_hd__xnor2_1_172/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_835 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_612/B sky130_fd_sc_hd__nor2_1_209/Y
+ sky130_fd_sc_hd__nand2_1_628/Y sky130_fd_sc_hd__xnor2_1_175/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_846 vssd1 vccd1 sky130_fd_sc_hd__nand2_2_13/Y sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__a22oi_1_221/Y sky130_fd_sc_hd__xor2_1_619/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_857 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_861/A2 sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__nand2_1_502/Y sky130_fd_sc_hd__xor2_1_630/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_868 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_646/A sky130_fd_sc_hd__nor2_1_227/Y
+ sky130_fd_sc_hd__nand2_1_689/Y sky130_fd_sc_hd__xnor2_1_194/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_879 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_656/A sky130_fd_sc_hd__nor2_1_239/Y
+ sky130_fd_sc_hd__nand2_1_744/Y sky130_fd_sc_hd__xnor2_1_209/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nand2b_2_3 sky130_fd_sc_hd__nor2_4_12/B sky130_fd_sc_hd__nand2b_2_3/Y
+ sky130_fd_sc_hd__nor2_4_12/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_2
Xsky130_fd_sc_hd__xor2_1_640 sky130_fd_sc_hd__xor2_1_640/B sky130_fd_sc_hd__xor2_1_640/X
+ sky130_fd_sc_hd__xor2_1_640/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_651 sky130_fd_sc_hd__xor2_1_651/B sky130_fd_sc_hd__xor2_1_651/X
+ sky130_fd_sc_hd__xor2_1_651/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_662 sky130_fd_sc_hd__xor2_1_662/B sky130_fd_sc_hd__xor2_1_662/X
+ sky130_fd_sc_hd__xor2_1_662/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_673 sky130_fd_sc_hd__mux2_2_38/X sky130_fd_sc_hd__xor2_1_673/X
+ sky130_fd_sc_hd__or2_0_78/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_684 sky130_fd_sc_hd__xor2_1_684/B sky130_fd_sc_hd__xor2_1_684/X
+ sky130_fd_sc_hd__xor2_1_684/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_695 la_data_out[49] sky130_fd_sc_hd__nand4_1_3/A sky130_fd_sc_hd__ha_2_56/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__and2_0_108 vccd1 vssd1 sky130_fd_sc_hd__and2_0_108/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_108/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_16 la_data_out[111] sky130_fd_sc_hd__conb_1_126/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_119 vccd1 vssd1 sky130_fd_sc_hd__and2_0_119/X sky130_fd_sc_hd__o21ai_2_0/B1
+ sky130_fd_sc_hd__and2_0_119/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_27 la_data_out[100] sky130_fd_sc_hd__conb_1_115/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_38 la_data_out[25] sky130_fd_sc_hd__conb_1_104/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_49 la_data_out[14] sky130_fd_sc_hd__conb_1_93/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__fa_2_3 sky130_fd_sc_hd__xor3_1_2/A sky130_fd_sc_hd__fa_2_4/B sky130_fd_sc_hd__fa_2_3/A
+ sky130_fd_sc_hd__fa_2_3/B sky130_fd_sc_hd__fa_2_3/CIN vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a211o_1_20 vssd1 vccd1 sky130_fd_sc_hd__fa_2_224/A sky130_fd_sc_hd__dfxtp_1_83/Q
+ sky130_fd_sc_hd__nor2_1_24/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_20/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__a211o_1_31 vssd1 vccd1 sky130_fd_sc_hd__xor3_1_15/A sky130_fd_sc_hd__dfxtp_1_94/Q
+ sky130_fd_sc_hd__nor2_1_35/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_31/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__clkinv_1_140 user_irq[2] sky130_fd_sc_hd__conb_1_2/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_151 sky130_fd_sc_hd__o22ai_1_32/B1 sky130_fd_sc_hd__dfxtp_1_188/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_162 sky130_fd_sc_hd__o21ai_1_5/A2 sky130_fd_sc_hd__dfxtp_1_125/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_173 sky130_fd_sc_hd__nor2_1_35/A sky130_fd_sc_hd__dfxtp_1_158/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_5 sky130_fd_sc_hd__buf_8_5/A sky130_fd_sc_hd__buf_8_5/X vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__a22o_1_7 sky130_fd_sc_hd__inv_2_66/Y sky130_fd_sc_hd__or2_0_95/B
+ sky130_fd_sc_hd__a22o_1_7/X sky130_fd_sc_hd__a22o_1_9/B2 sky130_fd_sc_hd__a22o_1_7/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_184 sky130_fd_sc_hd__o22ai_1_43/B1 sky130_fd_sc_hd__dfxtp_1_179/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_195 sky130_fd_sc_hd__o22ai_1_17/B1 sky130_fd_sc_hd__dfxtp_1_112/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_20 sky130_fd_sc_hd__inv_2_66/Y sky130_fd_sc_hd__xor2_1_660/X
+ sky130_fd_sc_hd__a22o_1_20/X sky130_fd_sc_hd__nor2_1_233/Y sky130_fd_sc_hd__xor2_1_652/X
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_31 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__buf_2_106/X
+ sky130_fd_sc_hd__a22o_1_31/X sky130_fd_sc_hd__a22o_1_31/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_42 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__buf_2_117/X
+ sky130_fd_sc_hd__a22o_1_42/X sky130_fd_sc_hd__a22o_1_42/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_53 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__buf_2_127/X
+ sky130_fd_sc_hd__a22o_1_53/X sky130_fd_sc_hd__a22o_1_53/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_64 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__buf_2_40/A
+ sky130_fd_sc_hd__a22o_1_64/X sky130_fd_sc_hd__ha_2_33/SUM sky130_fd_sc_hd__a22o_1_71/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_75 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__buf_6_92/X
+ sky130_fd_sc_hd__a22o_1_75/X sky130_fd_sc_hd__ha_2_21/SUM sky130_fd_sc_hd__nor2_1_269/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__nand4_1_3 sky130_fd_sc_hd__nand4_1_3/C sky130_fd_sc_hd__nand4_1_3/B
+ sky130_fd_sc_hd__nor4b_1_0/C sky130_fd_sc_hd__nand4_1_3/D sky130_fd_sc_hd__nand4_1_3/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__o21ai_1_109 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_109/A2 sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__a22oi_1_165/Y sky130_fd_sc_hd__and2_0_166/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_180 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_10 sky130_fd_sc_hd__nand2_1_10/Y sky130_fd_sc_hd__a22oi_1_2/Y
+ sky130_fd_sc_hd__a22oi_1_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_191 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_21 sky130_fd_sc_hd__nand2_8_1/A sky130_fd_sc_hd__nand2_1_7/B
+ sky130_fd_sc_hd__mux2_2_27/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_32 sky130_fd_sc_hd__buf_2_31/A sky130_fd_sc_hd__nand2_1_33/Y
+ sky130_fd_sc_hd__nand2_1_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_43 sky130_fd_sc_hd__nand2_1_1/B sky130_fd_sc_hd__nand2_1_8/B
+ sky130_fd_sc_hd__or2_0_82/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_54 sky130_fd_sc_hd__nand2_1_54/Y sky130_fd_sc_hd__nand2_1_54/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_65 sky130_fd_sc_hd__nand2_1_65/Y sky130_fd_sc_hd__nand2_1_65/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_270 vssd1 vccd1 la_data_out[85] sky130_fd_sc_hd__xnor2_1_270/Y
+ la_data_out[71] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_76 sky130_fd_sc_hd__nand2_1_76/Y sky130_fd_sc_hd__nand2_1_76/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_281 vssd1 vccd1 sky130_fd_sc_hd__buf_2_207/X sky130_fd_sc_hd__xnor2_1_281/Y
+ sky130_fd_sc_hd__or2_0_80/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_87 sky130_fd_sc_hd__nand2_1_87/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__xnor2_2_1/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_292 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_292/B sky130_fd_sc_hd__xnor2_1_292/Y
+ sky130_fd_sc_hd__xnor2_1_292/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_98 sky130_fd_sc_hd__nand2_1_98/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__xnor2_1_82/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_309 sky130_fd_sc_hd__or2_0_95/A sky130_fd_sc_hd__dfxtp_1_323/CLK
+ sky130_fd_sc_hd__and2_0_286/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_610 vssd1 vccd1 sky130_fd_sc_hd__buf_2_7/X sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_610/B1 sky130_fd_sc_hd__xor2_1_401/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1190 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_621 vssd1 vccd1 sky130_fd_sc_hd__inv_2_28/Y sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_621/B1 sky130_fd_sc_hd__xor2_1_414/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_632 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_526/A sky130_fd_sc_hd__nor2_2_26/Y
+ sky130_fd_sc_hd__nand2_1_561/Y sky130_fd_sc_hd__xnor2_1_149/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_643 vssd1 vccd1 sky130_fd_sc_hd__inv_2_47/Y sky130_fd_sc_hd__nand2b_1_21/Y
+ sky130_fd_sc_hd__o21ai_1_643/B1 sky130_fd_sc_hd__xor2_1_430/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_654 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_3/Y sky130_fd_sc_hd__nand2b_1_20/Y
+ sky130_fd_sc_hd__o21ai_1_654/B1 sky130_fd_sc_hd__xor2_1_439/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_665 vssd1 vccd1 sky130_fd_sc_hd__inv_2_43/Y sky130_fd_sc_hd__nand2b_1_21/Y
+ sky130_fd_sc_hd__o21ai_1_665/B1 sky130_fd_sc_hd__xor2_1_448/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_676 vssd1 vccd1 sky130_fd_sc_hd__xor2_2_2/X sky130_fd_sc_hd__nand2b_1_15/Y
+ sky130_fd_sc_hd__o21ai_1_676/B1 sky130_fd_sc_hd__xor2_1_457/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_687 vssd1 vccd1 sky130_fd_sc_hd__inv_2_47/Y sky130_fd_sc_hd__nand2b_1_15/Y
+ sky130_fd_sc_hd__o21ai_1_687/B1 sky130_fd_sc_hd__xor2_1_466/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_698 vssd1 vccd1 sky130_fd_sc_hd__inv_2_51/Y sky130_fd_sc_hd__nand2b_1_16/Y
+ sky130_fd_sc_hd__o21ai_1_698/B1 sky130_fd_sc_hd__xor2_1_477/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_17 sky130_fd_sc_hd__or2_0_0/A sky130_fd_sc_hd__nor2_2_2/A sky130_fd_sc_hd__fa_2_17/A
+ sky130_fd_sc_hd__fa_2_17/B sky130_fd_sc_hd__fa_2_17/CIN vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_28 sky130_fd_sc_hd__fa_2_19/CIN sky130_fd_sc_hd__fa_2_30/A
+ sky130_fd_sc_hd__fa_2_28/A sky130_fd_sc_hd__fa_2_28/B sky130_fd_sc_hd__xor2_1_48/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_39 sky130_fd_sc_hd__fa_2_32/A sky130_fd_sc_hd__fa_2_40/B sky130_fd_sc_hd__fa_2_39/A
+ sky130_fd_sc_hd__fa_2_39/B sky130_fd_sc_hd__xor2_1_57/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_209 vccd1 vssd1 la_data_out[78] sky130_fd_sc_hd__mux2_4_4/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__xor2_1_470 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__fa_2_309/B
+ sky130_fd_sc_hd__xor2_1_470/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_481 sky130_fd_sc_hd__fa_2_379/A sky130_fd_sc_hd__fa_2_320/B
+ sky130_fd_sc_hd__xor2_1_481/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_492 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__xor2_1_492/X
+ sky130_fd_sc_hd__xor2_1_492/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a222oi_1_501 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__buf_2_21/X
+ sky130_fd_sc_hd__nor2_1_87/A sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__o21ai_1_795/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_512 vccd1 vssd1 sky130_fd_sc_hd__and3_4_18/X sky130_fd_sc_hd__or2_0_72/B
+ sky130_fd_sc_hd__or2_0_72/A sky130_fd_sc_hd__nor2_2_32/Y sky130_fd_sc_hd__or2_0_71/B
+ sky130_fd_sc_hd__o21ai_1_809/B1 sky130_fd_sc_hd__nor2b_2_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_523 vccd1 vssd1 sky130_fd_sc_hd__and3_4_20/X sky130_fd_sc_hd__or2_0_72/B
+ sky130_fd_sc_hd__or2_0_72/A sky130_fd_sc_hd__nor2_4_16/Y sky130_fd_sc_hd__or2_0_71/B
+ sky130_fd_sc_hd__o21ai_1_825/B1 sky130_fd_sc_hd__and2b_4_11/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_534 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__buf_8_0/A
+ sky130_fd_sc_hd__buf_4_6/X sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__buf_4_1/X
+ sky130_fd_sc_hd__o21ai_1_843/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_545 vccd1 vssd1 sky130_fd_sc_hd__inv_2_68/Y sky130_fd_sc_hd__dfxtp_1_425/Q
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__ha_2_9/A sky130_fd_sc_hd__dfxtp_1_457/Q
+ sky130_fd_sc_hd__clkinv_1_742/A sky130_fd_sc_hd__dfxtp_1_393/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_556 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_414/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_446/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_753/A sky130_fd_sc_hd__dfxtp_1_382/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_567 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_403/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_435/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_764/A sky130_fd_sc_hd__dfxtp_1_371/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_578 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_409/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_441/Q sky130_fd_sc_hd__clkbuf_1_32/X
+ sky130_fd_sc_hd__clkinv_1_775/A sky130_fd_sc_hd__dfxtp_1_377/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_589 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_398/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_430/Q sky130_fd_sc_hd__clkbuf_1_32/X
+ sky130_fd_sc_hd__clkinv_1_786/A sky130_fd_sc_hd__dfxtp_1_366/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nor2b_1_101 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_101/Y
+ sky130_fd_sc_hd__nor2b_1_101/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_112 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_112/Y
+ sky130_fd_sc_hd__nor2b_1_112/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__decap_12_18 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_123 la_data_out[45] sky130_fd_sc_hd__maj3_1_0/B sky130_fd_sc_hd__ha_2_52/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__decap_12_29 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_134 sky130_fd_sc_hd__clkinv_4_53/Y sky130_fd_sc_hd__nor2b_1_134/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_145 sky130_fd_sc_hd__clkinv_4_64/Y sky130_fd_sc_hd__nor2b_1_145/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_156 sky130_fd_sc_hd__clkinv_4_75/Y sky130_fd_sc_hd__nor2b_1_156/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__fah_1_14 sky130_fd_sc_hd__fah_1_13/CI sky130_fd_sc_hd__fah_1_14/B
+ sky130_fd_sc_hd__fah_1_14/A sky130_fd_sc_hd__fa_2_398/A sky130_fd_sc_hd__fah_1_14/CI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__fah_1
Xsky130_fd_sc_hd__buf_6_2 vccd1 vssd1 sky130_fd_sc_hd__buf_6_2/X sky130_fd_sc_hd__buf_6_2/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_18 vccd1 vssd1 sky130_fd_sc_hd__buf_8_55/A sky130_fd_sc_hd__buf_6_18/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_29 vccd1 vssd1 sky130_fd_sc_hd__buf_6_29/X sky130_fd_sc_hd__buf_8_47/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__sdlclkp_4_0 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_8_1/Y
+ sky130_fd_sc_hd__dfxtp_1_46/CLK sky130_fd_sc_hd__o21ai_1_0/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__clkinv_1_909 sky130_fd_sc_hd__clkinv_1_909/Y sky130_fd_sc_hd__clkinv_1_909/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_3 sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__nor2_1_3/Y
+ sky130_fd_sc_hd__nor2_4_1/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__dfxtp_1_106 sky130_fd_sc_hd__dfxtp_1_106/Q sky130_fd_sc_hd__dfxtp_1_99/CLK
+ sky130_fd_sc_hd__and2_0_158/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_117 sky130_fd_sc_hd__dfxtp_1_117/Q sky130_fd_sc_hd__dfxtp_1_118/CLK
+ sky130_fd_sc_hd__and2_0_212/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_128 sky130_fd_sc_hd__dfxtp_1_128/Q sky130_fd_sc_hd__dfxtp_1_146/CLK
+ sky130_fd_sc_hd__and2_0_115/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_139 sky130_fd_sc_hd__dfxtp_1_139/Q sky130_fd_sc_hd__dfxtp_1_141/CLK
+ sky130_fd_sc_hd__and2_0_168/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_440 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_476/A2 sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_440/B1 sky130_fd_sc_hd__xor2_1_245/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_451 vssd1 vccd1 sky130_fd_sc_hd__inv_2_31/Y sky130_fd_sc_hd__nand2b_1_14/Y
+ sky130_fd_sc_hd__o21ai_1_451/B1 sky130_fd_sc_hd__xor2_1_254/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_462 vssd1 vccd1 sky130_fd_sc_hd__buf_2_11/X sky130_fd_sc_hd__nand2b_1_13/Y
+ sky130_fd_sc_hd__o21ai_1_462/B1 sky130_fd_sc_hd__xor2_1_265/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_473 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_7/X sky130_fd_sc_hd__nand2_1_363/Y
+ sky130_fd_sc_hd__a21oi_1_78/Y sky130_fd_sc_hd__xnor2_1_79/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_3_0 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__o21ai_1_484 vssd1 vccd1 sky130_fd_sc_hd__inv_2_36/Y sky130_fd_sc_hd__nand2b_2_3/Y
+ sky130_fd_sc_hd__o21ai_1_484/B1 sky130_fd_sc_hd__xor2_1_285/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_495 vssd1 vccd1 sky130_fd_sc_hd__inv_2_37/Y sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_495/B1 sky130_fd_sc_hd__xor2_1_297/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_905 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_916 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_800 sky130_fd_sc_hd__xor2_1_678/B sky130_fd_sc_hd__nand2_1_801/Y
+ sky130_fd_sc_hd__nand2_1_800/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_927 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_811 sky130_fd_sc_hd__nand2_1_811/Y sky130_fd_sc_hd__or2_0_104/A
+ sky130_fd_sc_hd__or2_0_104/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_938 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_822 sky130_fd_sc_hd__xnor2_1_298/A sky130_fd_sc_hd__nand2_1_823/Y
+ sky130_fd_sc_hd__or2_0_107/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_949 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_833 sky130_fd_sc_hd__nand2_1_833/Y sky130_fd_sc_hd__nor2_1_264/A
+ sky130_fd_sc_hd__nor2_1_264/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_844 sky130_fd_sc_hd__buf_2_128/A sky130_fd_sc_hd__dfxtp_1_20/Q
+ sky130_fd_sc_hd__dfxtp_1_1/Q vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_855 sky130_fd_sc_hd__nand2_1_855/Y sky130_fd_sc_hd__nand2_1_856/Y
+ sky130_fd_sc_hd__nand3_1_5/C vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_866 sky130_fd_sc_hd__a21o_2_3/A2 sky130_fd_sc_hd__nand2_1_866/B
+ sky130_fd_sc_hd__a21o_2_2/B1 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o21ai_1_11 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_22/B1 sky130_fd_sc_hd__nor2_4_4/B
+ sky130_fd_sc_hd__o21ai_1_11/B1 sky130_fd_sc_hd__fa_2_72/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_22 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_11/B1 sky130_fd_sc_hd__nor2_4_4/B
+ sky130_fd_sc_hd__o21ai_1_22/B1 sky130_fd_sc_hd__fa_2_125/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_33 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_2/B1 sky130_fd_sc_hd__inv_2_53/A
+ sky130_fd_sc_hd__o21ai_1_33/B1 sky130_fd_sc_hd__o21ai_1_33/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_44 vssd1 vccd1 sky130_fd_sc_hd__inv_2_58/Y sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_44/B1 sky130_fd_sc_hd__o21ai_1_44/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_55 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_57/A2 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_95/Y sky130_fd_sc_hd__o21ai_1_55/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_66 vssd1 vccd1 sky130_fd_sc_hd__inv_2_56/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__o21ai_1_66/B1 sky130_fd_sc_hd__o21ai_1_66/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_77 vssd1 vccd1 sky130_fd_sc_hd__inv_2_61/Y sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__o21ai_1_77/B1 sky130_fd_sc_hd__o21ai_1_77/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_88 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_89/A2 sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__o21ai_1_88/B1 sky130_fd_sc_hd__o21ai_1_88/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_99 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_99/A2 sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__o21ai_1_99/B1 sky130_fd_sc_hd__o21ai_1_99/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nand2_4_4 sky130_fd_sc_hd__nand2_4_4/Y sky130_fd_sc_hd__or2_0_25/X
+ sky130_fd_sc_hd__xnor2_1_4/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_4
Xsky130_fd_sc_hd__a222oi_1_320 vccd1 vssd1 sky130_fd_sc_hd__and3_4_16/X sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__buf_8_0/X sky130_fd_sc_hd__nor2_2_19/Y sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__o21ai_1_537/B1 sky130_fd_sc_hd__nor2b_2_3/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_260 vssd1 vccd1 sky130_fd_sc_hd__buf_12_39/A sky130_fd_sc_hd__clkbuf_1_260/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_331 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__and2_0_38/A
+ sky130_fd_sc_hd__and2_0_49/A sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__and2_0_45/A
+ sky130_fd_sc_hd__o21ai_1_552/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_271 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_271/X sky130_fd_sc_hd__inv_2_179/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_342 vccd1 vssd1 sky130_fd_sc_hd__and3_4_10/X sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__buf_4_7/X sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__buf_4_0/X
+ sky130_fd_sc_hd__o21ai_1_568/B1 sky130_fd_sc_hd__and2b_4_7/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_282 vssd1 vccd1 sky130_fd_sc_hd__buf_8_111/A sky130_fd_sc_hd__clkbuf_1_282/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_353 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__buf_6_1/X sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__and2_0_38/A
+ sky130_fd_sc_hd__o21ai_1_584/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_293 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_294/A sky130_fd_sc_hd__buf_8_154/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_364 vccd1 vssd1 sky130_fd_sc_hd__and3_4_11/X sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__inv_6_0/Y sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__o21ai_1_603/B1 sky130_fd_sc_hd__and2b_4_8/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_375 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__buf_6_2/X sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__buf_4_7/X
+ sky130_fd_sc_hd__o21ai_1_620/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_386 vccd1 vssd1 sky130_fd_sc_hd__and3_4_21/X sky130_fd_sc_hd__or2_0_60/B
+ sky130_fd_sc_hd__or2_0_60/A sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__or2_0_61/A
+ sky130_fd_sc_hd__o21ai_1_647/B1 sky130_fd_sc_hd__and2b_4_12/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_397 vccd1 vssd1 sky130_fd_sc_hd__and3_1_2/X sky130_fd_sc_hd__buf_2_25/A
+ sky130_fd_sc_hd__inv_6_0/Y sky130_fd_sc_hd__nor2_1_174/Y sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__o21ai_1_662/B1 sky130_fd_sc_hd__nor2b_1_14/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a21oi_2_10 sky130_fd_sc_hd__a21oi_2_10/B1 sky130_fd_sc_hd__or2_0_33/X
+ sky130_fd_sc_hd__xnor2_1_86/B sky130_fd_sc_hd__xor2_1_296/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_2
Xsky130_fd_sc_hd__and2_0_280 vccd1 vssd1 sky130_fd_sc_hd__and2_0_280/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__fa_2_417/SUM vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_291 vccd1 vssd1 sky130_fd_sc_hd__and2_0_291/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_12/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_12_506 sky130_fd_sc_hd__buf_12_506/A sky130_fd_sc_hd__buf_12_530/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_517 sky130_fd_sc_hd__buf_12_517/A sky130_fd_sc_hd__buf_12_517/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_528 sky130_fd_sc_hd__buf_12_528/A sky130_fd_sc_hd__buf_12_528/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_539 sky130_fd_sc_hd__buf_12_539/A sky130_fd_sc_hd__buf_12_539/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__nand2_1_107 sky130_fd_sc_hd__o21ai_1_79/B1 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__xnor2_1_91/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_706 sky130_fd_sc_hd__nand4_1_0/D sky130_fd_sc_hd__ha_2_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_118 sky130_fd_sc_hd__nand2_1_118/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__xnor2_1_98/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_717 sky130_fd_sc_hd__nor2b_1_96/A sky130_fd_sc_hd__xor2_1_677/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_129 sky130_fd_sc_hd__nand2_1_129/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_129/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_728 sky130_fd_sc_hd__nor2b_1_107/A sky130_fd_sc_hd__xnor2_1_297/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_739 sky130_fd_sc_hd__nor2b_1_118/A sky130_fd_sc_hd__xor2_1_688/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__or2_0_104 sky130_fd_sc_hd__or2_0_104/A sky130_fd_sc_hd__or2_0_104/X
+ sky130_fd_sc_hd__or2_0_104/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__o21ai_1_270 vssd1 vccd1 sky130_fd_sc_hd__inv_2_14/Y sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__o21ai_1_270/B1 sky130_fd_sc_hd__xor2_1_92/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_281 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_300/B1 sky130_fd_sc_hd__nor2_1_67/A
+ sky130_fd_sc_hd__nor2_1_66/Y sky130_fd_sc_hd__o21ai_1_281/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkinv_8_9 sky130_fd_sc_hd__clkinv_8_9/Y wbs_dat_i[29] vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__o21ai_1_292 vssd1 vccd1 sky130_fd_sc_hd__inv_2_13/Y sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__o21ai_1_292/B1 sky130_fd_sc_hd__xor2_1_113/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_702 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_713 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_724 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_735 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_746 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_630 sky130_fd_sc_hd__nand2_1_630/Y sky130_fd_sc_hd__buf_2_27/X
+ sky130_fd_sc_hd__buf_2_15/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_757 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_641 sky130_fd_sc_hd__xor2_1_624/B sky130_fd_sc_hd__nand2_1_642/Y
+ sky130_fd_sc_hd__or2_0_69/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_768 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_652 sky130_fd_sc_hd__xnor2_2_2/B sky130_fd_sc_hd__nand2_1_653/Y
+ sky130_fd_sc_hd__nand2_1_652/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_779 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_663 sky130_fd_sc_hd__nand2_1_663/Y sky130_fd_sc_hd__or2_0_73/A
+ sky130_fd_sc_hd__or2_0_73/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_674 sky130_fd_sc_hd__xnor2_1_191/A sky130_fd_sc_hd__nand2_1_675/Y
+ sky130_fd_sc_hd__or2_0_76/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_685 sky130_fd_sc_hd__nand2_1_685/Y sky130_fd_sc_hd__mux2_2_27/X
+ sky130_fd_sc_hd__mux2_2_47/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_696 sky130_fd_sc_hd__xor2_1_648/B sky130_fd_sc_hd__nand2_1_697/Y
+ sky130_fd_sc_hd__nand2_1_696/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_1701 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1712 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_11 sky130_fd_sc_hd__inv_2_11/A sky130_fd_sc_hd__inv_2_11/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1723 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_22 sky130_fd_sc_hd__inv_2_22/A sky130_fd_sc_hd__inv_2_22/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1734 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_33 sky130_fd_sc_hd__inv_2_33/A sky130_fd_sc_hd__inv_2_33/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1745 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_44 sky130_fd_sc_hd__inv_2_44/A sky130_fd_sc_hd__inv_2_44/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1756 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_55 sky130_fd_sc_hd__inv_2_55/A sky130_fd_sc_hd__inv_2_55/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1767 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_66 sky130_fd_sc_hd__inv_2_66/A sky130_fd_sc_hd__inv_2_66/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_470 sky130_fd_sc_hd__ha_2_53/A sky130_fd_sc_hd__dfxtp_1_515/CLK
+ sky130_fd_sc_hd__and2_0_359/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1778 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_77 sky130_fd_sc_hd__inv_2_77/A sky130_fd_sc_hd__inv_2_77/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_481 la_data_out[48] sky130_fd_sc_hd__dfxtp_1_489/CLK sky130_fd_sc_hd__and2_0_366/X
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1789 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_2_1 sky130_fd_sc_hd__nand2_2_1/Y sky130_fd_sc_hd__nand2_2_1/A
+ sky130_fd_sc_hd__nand2_2_1/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__inv_2_88 la_data_out[41] sky130_fd_sc_hd__inv_2_90/A vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_492 la_data_out[41] sky130_fd_sc_hd__dfxtp_1_498/CLK sky130_fd_sc_hd__and2_0_368/X
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_99 sky130_fd_sc_hd__inv_4_18/Y sky130_fd_sc_hd__inv_2_99/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__a222oi_1_150 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__buf_4_2/X sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__o21ai_1_295/B1 sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_161 vccd1 vssd1 sky130_fd_sc_hd__and3_4_7/X sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__inv_6_0/Y sky130_fd_sc_hd__nor2_2_7/Y sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__o21ai_1_310/B1 sky130_fd_sc_hd__nor2b_2_1/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_172 vccd1 vssd1 sky130_fd_sc_hd__and3_4_2/X sky130_fd_sc_hd__nor2_2_4/B
+ sky130_fd_sc_hd__buf_2_4/A sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__o21ai_1_324/B1 sky130_fd_sc_hd__and2b_4_4/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_320 sky130_fd_sc_hd__fa_2_314/CIN sky130_fd_sc_hd__fa_2_322/CIN
+ sky130_fd_sc_hd__fa_2_320/A sky130_fd_sc_hd__fa_2_320/B sky130_fd_sc_hd__xor2_1_480/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_183 vccd1 vssd1 sky130_fd_sc_hd__and3_4_1/X sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__buf_4_6/X sky130_fd_sc_hd__nor2_2_9/Y sky130_fd_sc_hd__and2_0_25/A
+ sky130_fd_sc_hd__o21ai_1_340/B1 sky130_fd_sc_hd__and2b_4_3/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_331 sky130_fd_sc_hd__fa_2_318/A sky130_fd_sc_hd__fa_2_330/B
+ sky130_fd_sc_hd__fa_2_331/A sky130_fd_sc_hd__fa_2_331/B sky130_fd_sc_hd__xor2_1_493/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_194 vccd1 vssd1 sky130_fd_sc_hd__and3_4_2/X sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__buf_4_6/X sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__and2_0_25/A
+ sky130_fd_sc_hd__o21ai_1_358/B1 sky130_fd_sc_hd__and2b_4_4/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_342 sky130_fd_sc_hd__fa_2_337/CIN sky130_fd_sc_hd__fa_2_348/A
+ sky130_fd_sc_hd__fa_2_342/A sky130_fd_sc_hd__fa_2_342/B sky130_fd_sc_hd__fa_2_342/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_353 sky130_fd_sc_hd__fa_2_342/CIN sky130_fd_sc_hd__fa_2_353/SUM
+ sky130_fd_sc_hd__fa_2_353/A sky130_fd_sc_hd__fa_2_353/B sky130_fd_sc_hd__xor2_1_523/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_364 sky130_fd_sc_hd__fa_2_360/CIN sky130_fd_sc_hd__fa_2_367/B
+ sky130_fd_sc_hd__fa_2_364/A sky130_fd_sc_hd__fa_2_364/B sky130_fd_sc_hd__xor2_1_540/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_375 sky130_fd_sc_hd__fa_2_371/CIN sky130_fd_sc_hd__fah_1_7/A
+ sky130_fd_sc_hd__fa_2_375/A sky130_fd_sc_hd__fa_2_375/B sky130_fd_sc_hd__xor2_1_554/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_16 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_8_3/Y
+ sky130_fd_sc_hd__clkinv_2_8/A sky130_fd_sc_hd__o21ai_2_1/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_386 sky130_fd_sc_hd__fah_1_6/A sky130_fd_sc_hd__fa_2_387/A
+ sky130_fd_sc_hd__fa_2_386/A sky130_fd_sc_hd__fa_2_386/B sky130_fd_sc_hd__xor2_1_570/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_27 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_8_5/Y
+ sky130_fd_sc_hd__dfxtp_1_264/CLK sky130_fd_sc_hd__o21ai_2_4/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_397 sky130_fd_sc_hd__fa_2_395/B sky130_fd_sc_hd__fah_1_9/CI
+ sky130_fd_sc_hd__fa_2_397/A sky130_fd_sc_hd__fa_2_397/B sky130_fd_sc_hd__xor2_1_586/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_38 sky130_fd_sc_hd__conb_1_145/LO sky130_fd_sc_hd__clkinv_4_11/Y
+ sky130_fd_sc_hd__dfxtp_1_375/CLK sky130_fd_sc_hd__o21ai_1_892/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_49 sky130_fd_sc_hd__conb_1_148/LO sky130_fd_sc_hd__clkinv_8_67/A
+ sky130_fd_sc_hd__dfxtp_1_509/CLK sky130_fd_sc_hd__o21ai_1_913/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__clkinv_8_80 sky130_fd_sc_hd__clkinv_8_81/A sky130_fd_sc_hd__clkinv_8_80/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__nor2_1_107 sky130_fd_sc_hd__nor2_1_112/A sky130_fd_sc_hd__nor2_1_107/Y
+ sky130_fd_sc_hd__nor2_1_107/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_118 sky130_fd_sc_hd__nor2_1_118/B sky130_fd_sc_hd__nor2_1_118/Y
+ sky130_fd_sc_hd__nor2_1_120/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_129 sky130_fd_sc_hd__nor2_1_73/B sky130_fd_sc_hd__nor2_1_129/Y
+ sky130_fd_sc_hd__buf_4_3/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_16 sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__dfxtp_1_283/Q sky130_fd_sc_hd__o211ai_1_7/Y sky130_fd_sc_hd__nand2_1_14/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_27 sky130_fd_sc_hd__nor2_4_0/Y sky130_fd_sc_hd__nor2_2_0/Y
+ sky130_fd_sc_hd__dfxtp_1_327/Q sky130_fd_sc_hd__nor2_1_241/A sky130_fd_sc_hd__nand2_2_5/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_38 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__clkbuf_1_25/X
+ sky130_fd_sc_hd__nand2_1_80/B sky130_fd_sc_hd__dfxtp_1_130/Q sky130_fd_sc_hd__a22oi_1_38/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_49 sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__dfxtp_1_103/Q sky130_fd_sc_hd__dfxtp_1_71/Q sky130_fd_sc_hd__a22oi_1_49/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_303 sky130_fd_sc_hd__buf_12_303/A sky130_fd_sc_hd__buf_12_303/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_314 sky130_fd_sc_hd__bufinv_8_0/Y sky130_fd_sc_hd__buf_12_490/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_325 sky130_fd_sc_hd__buf_12_325/A sky130_fd_sc_hd__buf_12_325/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_336 sky130_fd_sc_hd__buf_12_41/X sky130_fd_sc_hd__buf_12_587/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_347 sky130_fd_sc_hd__buf_12_347/A sky130_fd_sc_hd__buf_12_585/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_206 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__nor2b_1_11/Y sky130_fd_sc_hd__nor2_1_130/Y sky130_fd_sc_hd__a22oi_1_206/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_358 sky130_fd_sc_hd__buf_12_358/A sky130_fd_sc_hd__buf_12_644/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_217 sky130_fd_sc_hd__or2_0_72/B sky130_fd_sc_hd__or2_0_72/A
+ sky130_fd_sc_hd__nor2b_1_17/Y sky130_fd_sc_hd__nor2_1_186/Y sky130_fd_sc_hd__a22oi_1_217/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_369 sky130_fd_sc_hd__buf_12_369/A sky130_fd_sc_hd__buf_12_505/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_503 sky130_fd_sc_hd__clkinv_1_503/Y sky130_fd_sc_hd__nand2_1_480/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_514 sky130_fd_sc_hd__nand2_1_602/A sky130_fd_sc_hd__nor2_2_28/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_525 sky130_fd_sc_hd__nand2_1_517/A sky130_fd_sc_hd__nor2_2_22/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_536 sky130_fd_sc_hd__nor2_1_171/A sky130_fd_sc_hd__nand2_1_543/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_547 sky130_fd_sc_hd__o21ai_1_723/A2 sky130_fd_sc_hd__xnor2_1_146/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_558 sky130_fd_sc_hd__o21ai_1_751/A2 sky130_fd_sc_hd__xnor2_1_152/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_569 sky130_fd_sc_hd__a21oi_2_18/B1 sky130_fd_sc_hd__nand2_1_576/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_50 sky130_fd_sc_hd__nor2_1_51/B sky130_fd_sc_hd__nor2_1_50/Y
+ sky130_fd_sc_hd__nor2_1_50/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_61 sky130_fd_sc_hd__and3_4_4/A sky130_fd_sc_hd__nor2_1_61/Y
+ sky130_fd_sc_hd__and3_4_4/C vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_16 sky130_fd_sc_hd__inv_2_114/Y sky130_fd_sc_hd__buf_8_99/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_72 sky130_fd_sc_hd__and3_4_6/A sky130_fd_sc_hd__nor2_1_72/Y
+ sky130_fd_sc_hd__and3_4_6/C vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_27 sky130_fd_sc_hd__clkinv_4_27/A sky130_fd_sc_hd__clkinv_4_27/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_83 sky130_fd_sc_hd__nor2_1_83/B sky130_fd_sc_hd__nor2_1_83/Y
+ sky130_fd_sc_hd__nor2_1_83/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_38 sky130_fd_sc_hd__clkinv_8_17/A sky130_fd_sc_hd__clkinv_4_38/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_94 sky130_fd_sc_hd__nor2_1_94/B sky130_fd_sc_hd__nor2_1_94/Y
+ sky130_fd_sc_hd__nor2_1_94/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_49 sky130_fd_sc_hd__clkinv_4_49/A sky130_fd_sc_hd__clkinv_4_49/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_1008 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1019 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21a_1_4 sky130_fd_sc_hd__o21a_1_4/X sky130_fd_sc_hd__or2_0_55/A
+ sky130_fd_sc_hd__o21a_1_4/B1 sky130_fd_sc_hd__o21a_1_4/A2 vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__decap_12_510 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_521 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_532 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_543 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_554 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_565 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_576 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_460 sky130_fd_sc_hd__xor2_1_403/A sky130_fd_sc_hd__nand2_1_461/Y
+ sky130_fd_sc_hd__nand2_1_460/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_587 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_471 sky130_fd_sc_hd__nand2_1_471/Y sky130_fd_sc_hd__or2_0_49/A
+ sky130_fd_sc_hd__or2_0_49/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_598 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_482 sky130_fd_sc_hd__nand2_1_482/Y sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__inv_6_0/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_493 sky130_fd_sc_hd__nand2_1_493/Y sky130_fd_sc_hd__nor2_1_174/Y
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_40 sky130_fd_sc_hd__or2_0_74/A sky130_fd_sc_hd__fa_2_471/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_51 sky130_fd_sc_hd__mux2_2_8/X sky130_fd_sc_hd__nor2b_1_51/Y
+ sky130_fd_sc_hd__buf_2_214/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_62 sky130_fd_sc_hd__mux2_2_38/X sky130_fd_sc_hd__fa_2_482/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_73 sky130_fd_sc_hd__or2_1_10/B sky130_fd_sc_hd__nor2b_1_73/Y
+ sky130_fd_sc_hd__mux2_4_5/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1040 sky130_fd_sc_hd__clkinv_4_34/A sky130_fd_sc_hd__inv_2_113/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_84 sky130_fd_sc_hd__or2_0_84/B sky130_fd_sc_hd__or2_0_112/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1051 sky130_fd_sc_hd__inv_2_184/A sky130_fd_sc_hd__clkbuf_1_269/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_95 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_95/Y
+ sky130_fd_sc_hd__nor2b_1_95/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1062 sky130_fd_sc_hd__inv_16_5/A sky130_fd_sc_hd__buf_8_151/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_3 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_3/B sky130_fd_sc_hd__buf_2_3/A
+ sky130_fd_sc_hd__xnor2_1_3/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_1520 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1073 sky130_fd_sc_hd__o21ai_1_914/A2 sky130_fd_sc_hd__ha_2_45/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1531 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1084 sky130_fd_sc_hd__maj3_1_3/B la_data_out[50] vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1542 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1095 sky130_fd_sc_hd__and2_0_354/A sky130_fd_sc_hd__inv_2_105/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1553 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1564 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1575 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1586 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1597 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__fa_2_150 sky130_fd_sc_hd__xor3_1_16/B sky130_fd_sc_hd__fa_2_150/SUM
+ sky130_fd_sc_hd__fa_2_150/A sky130_fd_sc_hd__fa_2_150/B sky130_fd_sc_hd__fa_2_150/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_161 sky130_fd_sc_hd__fa_2_154/B sky130_fd_sc_hd__fa_2_164/A
+ sky130_fd_sc_hd__fa_2_161/A sky130_fd_sc_hd__fa_2_161/B sky130_fd_sc_hd__fa_2_161/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and3_4_0 sky130_fd_sc_hd__and3_4_0/A sky130_fd_sc_hd__nor2_4_8/B
+ sky130_fd_sc_hd__or2b_2_0/A sky130_fd_sc_hd__and3_4_0/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__dfxtp_1_18 sky130_fd_sc_hd__dfxtp_1_18/Q sky130_fd_sc_hd__dfxtp_1_8/CLK
+ la_data_out[57] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_172 sky130_fd_sc_hd__fa_2_165/A sky130_fd_sc_hd__fa_2_171/B
+ sky130_fd_sc_hd__fa_2_172/A sky130_fd_sc_hd__fa_2_172/B sky130_fd_sc_hd__fa_2_172/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_29 sky130_fd_sc_hd__ha_2_9/B sky130_fd_sc_hd__dfxtp_1_29/CLK
+ sky130_fd_sc_hd__ha_2_46/B vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_183 sky130_fd_sc_hd__fa_2_177/B sky130_fd_sc_hd__fa_2_185/CIN
+ sky130_fd_sc_hd__fa_2_183/A sky130_fd_sc_hd__fa_2_183/B sky130_fd_sc_hd__fa_2_183/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_194 sky130_fd_sc_hd__fa_2_189/CIN sky130_fd_sc_hd__fa_2_201/A
+ sky130_fd_sc_hd__fa_2_194/A sky130_fd_sc_hd__fa_2_194/B sky130_fd_sc_hd__fa_2_199/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o22ai_1_60 sky130_fd_sc_hd__nor2_1_7/A sky130_fd_sc_hd__o22ai_1_3/A2
+ sky130_fd_sc_hd__o22ai_1_60/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_71 sky130_fd_sc_hd__nor2b_1_20/A sky130_fd_sc_hd__xnor2_1_226/Y
+ sky130_fd_sc_hd__fa_2_431/A sky130_fd_sc_hd__xnor2_1_222/Y sky130_fd_sc_hd__o22ai_1_78/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_82 sky130_fd_sc_hd__xnor2_2_5/Y sky130_fd_sc_hd__xnor2_1_243/Y
+ sky130_fd_sc_hd__o22ai_1_82/Y sky130_fd_sc_hd__xnor2_1_232/Y sky130_fd_sc_hd__o22ai_1_95/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_93 sky130_fd_sc_hd__xnor2_2_6/Y sky130_fd_sc_hd__xnor2_1_246/Y
+ sky130_fd_sc_hd__fa_2_442/A sky130_fd_sc_hd__xnor2_1_240/Y sky130_fd_sc_hd__o22ai_1_98/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_4_40 vccd1 vssd1 sky130_fd_sc_hd__buf_4_40/X wbs_dat_i[0] vssd1
+ vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_12_100 sky130_fd_sc_hd__buf_8_34/X sky130_fd_sc_hd__buf_12_100/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_111 sky130_fd_sc_hd__buf_8_102/X sky130_fd_sc_hd__buf_12_388/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_sram_1kbyte_1rw1r_32x256_8_8 sky130_fd_sc_hd__inv_8_1/Y sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__buf_12_630/X sky130_fd_sc_hd__buf_12_572/X sky130_fd_sc_hd__buf_12_667/X
+ sky130_fd_sc_hd__buf_12_636/X sky130_fd_sc_hd__buf_12_401/X sky130_fd_sc_hd__buf_12_673/X
+ sky130_fd_sc_hd__buf_12_648/X sky130_fd_sc_hd__clkinv_1_956/Y sky130_fd_sc_hd__buf_12_657/X
+ sky130_fd_sc_hd__buf_12_589/X sky130_fd_sc_hd__buf_12_591/X vccd1 sky130_fd_sc_hd__clkinv_8_16/Y
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[16] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[17]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[18] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[19]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[20] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[21]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[22] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[23]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[24] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[25]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[26] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[27]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[28] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[29]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[30] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[31]
+ sky130_fd_sc_hd__buf_12_557/X sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[1] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[2]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[3] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[4]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[5] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[6]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[7] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[8]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[9] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[10]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[11] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[12]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[13] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[14]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[15] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout1[0]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[10] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[11]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[12] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[13]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[14] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[15]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[16] sky130_fd_sc_hd__buf_12_530/X sky130_fd_sc_hd__buf_12_115/X
+ sky130_fd_sc_hd__buf_12_92/X sky130_fd_sc_hd__buf_12_14/X sky130_fd_sc_hd__buf_12_158/X
+ sky130_fd_sc_hd__clkinv_8_21/Y sky130_fd_sc_hd__clkbuf_4_19/X sky130_fd_sc_hd__clkbuf_4_19/X
+ sky130_fd_sc_hd__clkbuf_4_19/X sky130_fd_sc_hd__clkbuf_4_19/X sky130_fd_sc_hd__clkbuf_4_19/X
+ sky130_fd_sc_hd__clkbuf_4_19/X sky130_fd_sc_hd__clkbuf_4_19/X sky130_fd_sc_hd__clkbuf_4_19/X
+ sky130_fd_sc_hd__clkbuf_4_19/X sky130_fd_sc_hd__clkbuf_4_19/X sky130_fd_sc_hd__clkbuf_1_67/A
+ sky130_fd_sc_hd__clkbuf_1_67/A sky130_fd_sc_hd__clkbuf_4_16/A sky130_fd_sc_hd__buf_6_11/A
+ sky130_fd_sc_hd__buf_6_11/A sky130_fd_sc_hd__buf_6_11/A sky130_fd_sc_hd__buf_6_11/A
+ sky130_fd_sc_hd__buf_6_11/A sky130_fd_sc_hd__buf_6_11/A sky130_fd_sc_hd__buf_6_11/X
+ sky130_fd_sc_hd__buf_6_11/X sky130_fd_sc_hd__buf_6_11/X sky130_fd_sc_hd__buf_6_11/X
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[0] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[1]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[2] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[3]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[4] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[5]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[6] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[7]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[8] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[9]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[25] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[26]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[27] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[28]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[29] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[30]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[31] sky130_fd_sc_hd__buf_6_11/X sky130_fd_sc_hd__buf_6_11/X
+ sky130_fd_sc_hd__buf_6_11/X sky130_fd_sc_hd__buf_6_11/X sky130_fd_sc_hd__buf_6_11/X
+ sky130_fd_sc_hd__buf_6_11/X sky130_fd_sc_hd__buf_6_11/X sky130_fd_sc_hd__buf_6_11/X
+ sky130_fd_sc_hd__buf_6_11/X sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[17] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[18]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[19] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[20]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[21] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[22]
+ sky130_fd_sc_hd__buf_12_521/X sky130_fd_sc_hd__buf_12_582/X sky130_fd_sc_hd__buf_12_590/X
+ sky130_fd_sc_hd__buf_12_477/X sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[23] sky130_sram_1kbyte_1rw1r_32x256_8_8/dout0[24]
+ sky130_sram_1kbyte_1rw1r_32x256_8_8/sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/gnd_uq26
+ vssd1 sky130_sram_1kbyte_1rw1r_32x256_8
Xsky130_fd_sc_hd__buf_12_122 sky130_fd_sc_hd__buf_12_32/X sky130_fd_sc_hd__buf_12_448/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_133 sky130_fd_sc_hd__buf_12_46/X sky130_fd_sc_hd__buf_12_355/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_144 sky130_fd_sc_hd__buf_12_22/X sky130_fd_sc_hd__buf_12_390/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_155 sky130_fd_sc_hd__buf_8_48/X sky130_fd_sc_hd__buf_12_155/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_166 sky130_fd_sc_hd__buf_12_25/X sky130_fd_sc_hd__buf_12_276/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_4_3 sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__nor2_1_36/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_12_177 sky130_fd_sc_hd__buf_8_127/X sky130_fd_sc_hd__buf_12_421/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_188 sky130_fd_sc_hd__buf_6_26/X sky130_fd_sc_hd__buf_12_353/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_199 sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__buf_12_382/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_300 sky130_fd_sc_hd__and2_0_221/A sky130_fd_sc_hd__a222oi_1_44/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_311 sky130_fd_sc_hd__a21oi_1_50/B1 sky130_fd_sc_hd__nand2_1_249/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_322 sky130_fd_sc_hd__nor2_1_49/A sky130_fd_sc_hd__nand2_1_189/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_333 sky130_fd_sc_hd__o21ai_1_237/A2 sky130_fd_sc_hd__xnor2_1_16/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_344 sky130_fd_sc_hd__nand2_1_203/A sky130_fd_sc_hd__or2_0_5/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_355 sky130_fd_sc_hd__o21ai_1_295/A2 sky130_fd_sc_hd__xnor2_1_29/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_366 sky130_fd_sc_hd__nor2_1_76/B sky130_fd_sc_hd__nor2_1_78/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_377 sky130_fd_sc_hd__nand2_1_265/A sky130_fd_sc_hd__nor2_1_86/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_388 sky130_fd_sc_hd__xor2_1_187/B sky130_fd_sc_hd__o21ai_1_372/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_399 sky130_fd_sc_hd__a21oi_1_67/B1 sky130_fd_sc_hd__nand2_1_309/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_2_7 sky130_fd_sc_hd__a21oi_2_7/B1 sky130_fd_sc_hd__or2_0_28/X
+ sky130_fd_sc_hd__xnor2_1_73/B sky130_fd_sc_hd__a21oi_2_7/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_2
Xsky130_fd_sc_hd__clkinv_4_3 sky130_fd_sc_hd__clkinv_8_3/A sky130_fd_sc_hd__clkinv_4_3/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__or2_0_80 sky130_fd_sc_hd__or2_0_80/A sky130_fd_sc_hd__or2_0_80/X
+ sky130_fd_sc_hd__or2_0_80/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_91 sky130_fd_sc_hd__or2_0_91/A sky130_fd_sc_hd__or2_0_91/X
+ sky130_fd_sc_hd__or2_0_91/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__decap_12_340 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_351 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_362 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_373 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_384 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_395 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_107 sky130_fd_sc_hd__xor2_1_6/B sky130_fd_sc_hd__fa_2_79/B
+ sky130_fd_sc_hd__xor2_1_107/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_290 sky130_fd_sc_hd__nand2_1_290/Y sky130_fd_sc_hd__nor2_1_98/A
+ sky130_fd_sc_hd__nor2_1_98/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_118 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__fa_2_88/CIN
+ sky130_fd_sc_hd__xor2_1_118/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_129 sky130_fd_sc_hd__fa_2_110/A sky130_fd_sc_hd__fa_2_94/B
+ sky130_fd_sc_hd__xor2_1_129/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1350 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1361 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1372 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_803 vssd1 vccd1 sky130_fd_sc_hd__inv_2_51/Y sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_803/B1 sky130_fd_sc_hd__xor2_1_577/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1383 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_814 vssd1 vccd1 sky130_fd_sc_hd__inv_2_46/Y sky130_fd_sc_hd__nand2b_2_6/Y
+ sky130_fd_sc_hd__o21ai_1_814/B1 sky130_fd_sc_hd__xor2_1_589/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1394 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_825 vssd1 vccd1 sky130_fd_sc_hd__buf_2_13/X sky130_fd_sc_hd__nand2b_2_6/Y
+ sky130_fd_sc_hd__o21ai_1_825/B1 sky130_fd_sc_hd__xor2_1_599/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_836 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_2/Y sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__o21ai_1_836/B1 sky130_fd_sc_hd__xor2_1_607/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_847 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_2/Y sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_847/B1 sky130_fd_sc_hd__xor2_1_620/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_858 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_219/Y sky130_fd_sc_hd__o21a_1_5/X
+ sky130_fd_sc_hd__nand2_1_655/Y sky130_fd_sc_hd__xnor2_1_185/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_869 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_647/A sky130_fd_sc_hd__nor2_1_228/Y
+ sky130_fd_sc_hd__nand2_1_693/Y sky130_fd_sc_hd__xnor2_1_195/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nand2b_2_4 sky130_fd_sc_hd__nor2_4_13/B sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__nor2_4_13/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_2
Xsky130_fd_sc_hd__xor2_1_630 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__xor2_1_630/X
+ sky130_fd_sc_hd__xor2_1_630/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_641 sky130_fd_sc_hd__xor2_1_641/B sky130_fd_sc_hd__xor2_1_641/X
+ sky130_fd_sc_hd__xor2_1_641/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_652 sky130_fd_sc_hd__xor2_1_652/B sky130_fd_sc_hd__xor2_1_652/X
+ sky130_fd_sc_hd__xor2_1_652/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_663 sky130_fd_sc_hd__xor2_1_663/B sky130_fd_sc_hd__or2_0_90/B
+ sky130_fd_sc_hd__xor2_1_663/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_674 sky130_fd_sc_hd__xor2_1_674/B sky130_fd_sc_hd__xor2_1_674/X
+ sky130_fd_sc_hd__xor2_1_675/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_685 sky130_fd_sc_hd__xor2_1_685/B sky130_fd_sc_hd__xor2_1_685/X
+ sky130_fd_sc_hd__xor2_1_685/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_696 sky130_fd_sc_hd__ha_2_57/SUM sky130_fd_sc_hd__xor2_1_696/X
+ la_data_out[53] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__and2_0_109 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_64/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_109/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_17 la_data_out[110] sky130_fd_sc_hd__conb_1_125/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_28 la_data_out[99] sky130_fd_sc_hd__conb_1_114/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_39 la_data_out[24] sky130_fd_sc_hd__conb_1_103/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__fa_2_4 sky130_fd_sc_hd__xor3_1_1/A sky130_fd_sc_hd__fa_2_5/B sky130_fd_sc_hd__fa_2_4/A
+ sky130_fd_sc_hd__fa_2_4/B sky130_fd_sc_hd__fa_2_4/CIN vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a211o_1_10 vssd1 vccd1 sky130_fd_sc_hd__fa_2_267/A sky130_fd_sc_hd__dfxtp_1_73/Q
+ sky130_fd_sc_hd__nor2_1_14/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_10/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__a211o_1_21 vssd1 vccd1 sky130_fd_sc_hd__fa_2_217/B sky130_fd_sc_hd__dfxtp_1_84/Q
+ sky130_fd_sc_hd__nor2_1_25/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_21/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__clkinv_1_130 io_oeb[9] sky130_fd_sc_hd__conb_1_12/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_141 user_irq[1] sky130_fd_sc_hd__conb_1_1/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_152 sky130_fd_sc_hd__nor2_1_33/A sky130_fd_sc_hd__dfxtp_1_156/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_163 sky130_fd_sc_hd__o22ai_1_36/B1 sky130_fd_sc_hd__dfxtp_1_185/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_174 sky130_fd_sc_hd__o21ai_1_9/A2 sky130_fd_sc_hd__dfxtp_1_126/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_6 sky130_fd_sc_hd__buf_8_6/A sky130_fd_sc_hd__buf_8_6/X vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__a22o_1_8 sky130_fd_sc_hd__inv_2_66/Y sky130_fd_sc_hd__a22o_1_8/A2
+ sky130_fd_sc_hd__a22o_1_8/X sky130_fd_sc_hd__a22o_1_9/B2 sky130_fd_sc_hd__a22o_1_8/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_185 sky130_fd_sc_hd__nor2_1_24/A sky130_fd_sc_hd__dfxtp_1_147/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_10 sky130_fd_sc_hd__inv_2_66/Y sky130_fd_sc_hd__nor2_1_240/B
+ sky130_fd_sc_hd__a22o_1_10/X sky130_fd_sc_hd__a22o_1_9/B2 sky130_fd_sc_hd__xor2_1_657/X
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_21 sky130_fd_sc_hd__inv_2_66/Y sky130_fd_sc_hd__xor2_1_659/X
+ sky130_fd_sc_hd__a22o_1_21/X sky130_fd_sc_hd__nor2_1_233/Y sky130_fd_sc_hd__a22o_1_21/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_196 sky130_fd_sc_hd__o22ai_1_47/B1 sky130_fd_sc_hd__dfxtp_1_175/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_32 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__buf_2_107/X
+ sky130_fd_sc_hd__a22o_1_32/X sky130_fd_sc_hd__a22o_1_32/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_43 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__buf_2_118/X
+ sky130_fd_sc_hd__a22o_1_43/X sky130_fd_sc_hd__a22o_1_43/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_54 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__buf_2_45/A
+ sky130_fd_sc_hd__a22o_1_54/X sky130_fd_sc_hd__xor2_1_690/X sky130_fd_sc_hd__a22o_1_71/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_65 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__clkbuf_4_7/A
+ sky130_fd_sc_hd__a22o_1_65/X sky130_fd_sc_hd__ha_2_34/SUM sky130_fd_sc_hd__a22o_1_71/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_76 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__buf_2_183/X
+ sky130_fd_sc_hd__a22o_1_76/X sky130_fd_sc_hd__ha_2_22/SUM sky130_fd_sc_hd__nor2_1_269/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__nand4_1_4 sky130_fd_sc_hd__nor3_1_5/Y sky130_fd_sc_hd__nor4_1_2/Y
+ sky130_fd_sc_hd__nor4b_2_0/C sky130_fd_sc_hd__nor4_1_1/Y sky130_fd_sc_hd__nor4_1_3/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__clkinv_2_0 sky130_fd_sc_hd__clkinv_2_0/Y sky130_fd_sc_hd__clkinv_2_0/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__decap_12_170 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_181 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_11 sky130_fd_sc_hd__nand2_1_11/Y sky130_fd_sc_hd__a22oi_1_8/Y
+ sky130_fd_sc_hd__a22oi_1_9/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_192 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_22 sky130_fd_sc_hd__nand2_8_2/B sky130_fd_sc_hd__nand2_1_8/B
+ sky130_fd_sc_hd__or2_0_78/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_33 sky130_fd_sc_hd__nand2_1_33/Y sky130_fd_sc_hd__nand2_1_8/B
+ sky130_fd_sc_hd__mux2_2_48/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_44 sky130_fd_sc_hd__inv_2_64/A sky130_fd_sc_hd__nand2_1_45/Y
+ sky130_fd_sc_hd__nand2_1_46/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_55 sky130_fd_sc_hd__nand2_1_55/Y sky130_fd_sc_hd__nand2_1_55/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_260 vssd1 vccd1 la_data_out[77] sky130_fd_sc_hd__xnor2_1_260/Y
+ sky130_fd_sc_hd__mux2_2_24/X vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_66 sky130_fd_sc_hd__nand2_1_66/Y sky130_fd_sc_hd__nand2_1_66/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_271 vssd1 vccd1 la_data_out[67] sky130_fd_sc_hd__xnor2_1_271/Y
+ sky130_fd_sc_hd__or2_0_78/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_77 sky130_fd_sc_hd__nand2_1_77/Y sky130_fd_sc_hd__nand2_1_77/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_282 vssd1 vccd1 la_data_out[79] sky130_fd_sc_hd__xnor2_1_282/Y
+ sky130_fd_sc_hd__or2_0_78/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_88 sky130_fd_sc_hd__nand2_1_88/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__xor2_1_234/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_293 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_293/B sky130_fd_sc_hd__xnor2_1_293/Y
+ sky130_fd_sc_hd__xnor2_1_293/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_99 sky130_fd_sc_hd__nand2_1_99/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__xnor2_1_82/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o21ai_1_600 vssd1 vccd1 sky130_fd_sc_hd__inv_2_42/Y sky130_fd_sc_hd__nor2_2_18/Y
+ sky130_fd_sc_hd__nand2_1_453/Y sky130_fd_sc_hd__xnor2_1_112/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1180 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_611 vssd1 vccd1 sky130_fd_sc_hd__inv_2_29/Y sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_611/B1 sky130_fd_sc_hd__xor2_1_402/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1191 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_622 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_66/A sky130_fd_sc_hd__nor2_1_161/Y
+ sky130_fd_sc_hd__nand2_1_482/Y sky130_fd_sc_hd__xnor2_1_121/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_633 vssd1 vccd1 sky130_fd_sc_hd__nor2_2_29/Y sky130_fd_sc_hd__nand2_1_602/B
+ sky130_fd_sc_hd__nand2_1_598/Y sky130_fd_sc_hd__o21ai_1_633/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_644 vssd1 vccd1 sky130_fd_sc_hd__inv_2_44/Y sky130_fd_sc_hd__nand2b_1_20/Y
+ sky130_fd_sc_hd__o21ai_1_644/B1 sky130_fd_sc_hd__xor2_1_431/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_655 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_691/A2 sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_655/B1 sky130_fd_sc_hd__xor2_1_440/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_666 vssd1 vccd1 sky130_fd_sc_hd__buf_2_13/X sky130_fd_sc_hd__nand2b_1_18/Y
+ sky130_fd_sc_hd__o21ai_1_666/B1 sky130_fd_sc_hd__xor2_1_449/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_677 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_713/A2 sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_677/B1 sky130_fd_sc_hd__xor2_1_458/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_688 vssd1 vccd1 sky130_fd_sc_hd__inv_2_44/Y sky130_fd_sc_hd__nand2b_1_21/Y
+ sky130_fd_sc_hd__o21ai_1_688/B1 sky130_fd_sc_hd__xor2_1_467/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_699 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_9/X sky130_fd_sc_hd__nand2b_1_20/Y
+ sky130_fd_sc_hd__o21ai_1_699/B1 sky130_fd_sc_hd__xor2_1_478/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_18 sky130_fd_sc_hd__nor2_2_2/B sky130_fd_sc_hd__or2_0_1/B sky130_fd_sc_hd__fa_2_18/A
+ sky130_fd_sc_hd__fa_2_18/B sky130_fd_sc_hd__fa_2_25/SUM vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_29 sky130_fd_sc_hd__fa_2_24/CIN sky130_fd_sc_hd__fa_2_34/A
+ sky130_fd_sc_hd__fa_2_29/A sky130_fd_sc_hd__fa_2_29/B sky130_fd_sc_hd__xor2_1_46/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__xor2_1_460 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__fa_2_302/A
+ sky130_fd_sc_hd__xor2_1_460/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_471 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__fa_2_309/A
+ sky130_fd_sc_hd__xor2_1_471/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_482 sky130_fd_sc_hd__fah_1_14/A sky130_fd_sc_hd__fa_2_320/A
+ sky130_fd_sc_hd__xor2_1_482/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_493 sky130_fd_sc_hd__fa_2_379/A sky130_fd_sc_hd__xor2_1_493/X
+ sky130_fd_sc_hd__xor2_1_493/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a222oi_1_502 vccd1 vssd1 sky130_fd_sc_hd__and3_4_21/X sky130_fd_sc_hd__buf_2_15/X
+ sky130_fd_sc_hd__buf_2_4/A sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__buf_2_20/X
+ sky130_fd_sc_hd__o21ai_1_796/B1 sky130_fd_sc_hd__and2b_4_12/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_513 vccd1 vssd1 sky130_fd_sc_hd__and3_4_20/X sky130_fd_sc_hd__buf_2_29/X
+ sky130_fd_sc_hd__buf_2_30/X sky130_fd_sc_hd__nor2_4_16/Y sky130_fd_sc_hd__buf_2_26/X
+ sky130_fd_sc_hd__o21ai_1_810/B1 sky130_fd_sc_hd__and2b_4_11/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__dfxtp_4_0 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_4_0/D sky130_fd_sc_hd__dfxtp_4_3/CLK
+ sky130_fd_sc_hd__fa_2_414/A vssd1 vccd1 sky130_fd_sc_hd__dfxtp_4
Xsky130_fd_sc_hd__a222oi_1_524 vccd1 vssd1 sky130_fd_sc_hd__and3_4_21/X sky130_fd_sc_hd__buf_2_29/X
+ sky130_fd_sc_hd__buf_2_30/X sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__buf_4_7/X
+ sky130_fd_sc_hd__o21ai_1_826/B1 sky130_fd_sc_hd__and2b_4_12/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_535 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__buf_4_1/X
+ sky130_fd_sc_hd__buf_4_0/A sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__buf_2_27/A
+ sky130_fd_sc_hd__o21ai_1_844/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_546 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_424/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_456/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_743/A sky130_fd_sc_hd__dfxtp_1_392/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_557 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_413/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_445/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_754/A sky130_fd_sc_hd__dfxtp_1_381/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_568 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_402/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_434/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_765/A sky130_fd_sc_hd__dfxtp_1_370/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_579 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_411/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_443/Q sky130_fd_sc_hd__clkbuf_1_32/X
+ sky130_fd_sc_hd__clkinv_1_776/A sky130_fd_sc_hd__dfxtp_1_379/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nor2b_1_102 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_102/Y
+ sky130_fd_sc_hd__nor2b_1_102/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_113 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_113/Y
+ sky130_fd_sc_hd__nor2b_1_113/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__decap_12_19 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_124 la_data_out[54] sky130_fd_sc_hd__maj3_1_2/B sky130_fd_sc_hd__ha_2_60/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_135 sky130_fd_sc_hd__clkinv_4_54/Y sky130_fd_sc_hd__nor2b_1_135/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_146 sky130_fd_sc_hd__clkinv_4_65/Y sky130_fd_sc_hd__nor2b_1_146/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_157 sky130_fd_sc_hd__clkinv_4_76/Y sky130_fd_sc_hd__nor2b_1_157/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__fah_1_15 sky130_fd_sc_hd__fah_1_12/CI sky130_fd_sc_hd__fah_1_15/B
+ sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__fa_2_404/A sky130_fd_sc_hd__fah_1_15/CI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__fah_1
Xsky130_fd_sc_hd__buf_6_3 vccd1 vssd1 sky130_fd_sc_hd__buf_6_3/X sky130_fd_sc_hd__buf_6_3/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_19 vccd1 vssd1 sky130_fd_sc_hd__buf_6_19/X sky130_fd_sc_hd__buf_6_19/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__clkinv_2_60 sky130_fd_sc_hd__clkinv_2_60/Y sky130_fd_sc_hd__clkinv_2_60/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__sdlclkp_4_1 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_8_3/Y
+ sky130_fd_sc_hd__dfxtp_1_57/CLK sky130_fd_sc_hd__o21ai_1_0/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_4 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_4/Y
+ sky130_fd_sc_hd__nor2_1_4/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__dfxtp_1_107 sky130_fd_sc_hd__dfxtp_1_107/Q sky130_fd_sc_hd__dfxtp_1_99/CLK
+ sky130_fd_sc_hd__and2_0_163/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_118 sky130_fd_sc_hd__dfxtp_1_118/Q sky130_fd_sc_hd__dfxtp_1_118/CLK
+ sky130_fd_sc_hd__and2_0_218/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_129 sky130_fd_sc_hd__dfxtp_1_129/Q sky130_fd_sc_hd__dfxtp_1_146/CLK
+ sky130_fd_sc_hd__and2_0_120/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_430 vssd1 vccd1 sky130_fd_sc_hd__inv_2_29/Y sky130_fd_sc_hd__nand2b_1_12/Y
+ sky130_fd_sc_hd__o21ai_1_430/B1 sky130_fd_sc_hd__xor2_1_237/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_441 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_505/A2 sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_441/B1 sky130_fd_sc_hd__xor2_1_246/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_452 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_486/A2 sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_452/B1 sky130_fd_sc_hd__xor2_1_256/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_463 vssd1 vccd1 sky130_fd_sc_hd__buf_2_9/X sky130_fd_sc_hd__nand2b_1_14/Y
+ sky130_fd_sc_hd__o21ai_1_463/B1 sky130_fd_sc_hd__xor2_1_266/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_474 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_119/Y sky130_fd_sc_hd__nor2_1_120/Y
+ sky130_fd_sc_hd__nand2_1_371/Y sky130_fd_sc_hd__o21ai_1_474/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_3_1 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__o21ai_1_485 vssd1 vccd1 sky130_fd_sc_hd__inv_2_41/Y sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_485/B1 sky130_fd_sc_hd__xor2_1_286/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_496 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_496/A2 sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_496/B1 sky130_fd_sc_hd__xor2_1_298/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_906 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_917 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_801 sky130_fd_sc_hd__nand2_1_801/Y sky130_fd_sc_hd__nor2_1_256/A
+ sky130_fd_sc_hd__nor2_1_256/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_928 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_812 sky130_fd_sc_hd__xor2_1_681/B sky130_fd_sc_hd__nand2_1_813/Y
+ sky130_fd_sc_hd__nand2_1_812/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_939 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_823 sky130_fd_sc_hd__nand2_1_823/Y sky130_fd_sc_hd__or2_0_107/A
+ sky130_fd_sc_hd__or2_0_107/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_834 sky130_fd_sc_hd__xnor2_1_301/A sky130_fd_sc_hd__nand2_1_835/Y
+ sky130_fd_sc_hd__or2_0_110/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_845 sky130_fd_sc_hd__nand2_1_845/Y sky130_fd_sc_hd__nand2b_1_31/B
+ sky130_fd_sc_hd__nand2_1_845/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_856 sky130_fd_sc_hd__nand2_1_856/Y sky130_fd_sc_hd__nor2_1_268/B
+ sky130_fd_sc_hd__nor2_1_275/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o21ai_1_12 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_21/B1 sky130_fd_sc_hd__nor2_4_4/B
+ sky130_fd_sc_hd__o21ai_1_12/B1 sky130_fd_sc_hd__fa_2_75/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_23 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_10/B1 sky130_fd_sc_hd__nor2_4_4/B
+ sky130_fd_sc_hd__o21ai_1_23/B1 sky130_fd_sc_hd__fa_2_127/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_34 vssd1 vccd1 sky130_fd_sc_hd__inv_2_62/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_84/Y sky130_fd_sc_hd__and2_0_2/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_45 vssd1 vccd1 sky130_fd_sc_hd__inv_2_58/Y sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__o21ai_1_45/B1 sky130_fd_sc_hd__and2_0_8/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_56 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_57/A2 sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_56/B1 sky130_fd_sc_hd__o21ai_1_56/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_67 vssd1 vccd1 sky130_fd_sc_hd__inv_2_56/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__o21ai_1_67/B1 sky130_fd_sc_hd__o21ai_1_67/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_290 sky130_fd_sc_hd__fa_2_198/A sky130_fd_sc_hd__xor2_1_290/X
+ sky130_fd_sc_hd__xor2_1_290/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__o21ai_1_78 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_81/A2 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__o21ai_1_78/B1 sky130_fd_sc_hd__o21ai_1_78/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_89 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_89/A2 sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_89/B1 sky130_fd_sc_hd__o21ai_1_89/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_310 vccd1 vssd1 sky130_fd_sc_hd__and3_4_17/X sky130_fd_sc_hd__buf_4_0/X
+ sky130_fd_sc_hd__buf_2_23/X sky130_fd_sc_hd__nor2_2_20/Y sky130_fd_sc_hd__buf_2_31/X
+ sky130_fd_sc_hd__o21ai_1_525/B1 sky130_fd_sc_hd__nor2b_2_4/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_250 vssd1 vccd1 sky130_fd_sc_hd__buf_12_43/A sky130_fd_sc_hd__buf_2_156/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_321 vccd1 vssd1 sky130_fd_sc_hd__and3_4_10/X sky130_fd_sc_hd__buf_2_31/X
+ sky130_fd_sc_hd__buf_2_19/X sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__o21ai_1_539/B1 sky130_fd_sc_hd__and2b_4_7/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_261 vssd1 vccd1 sky130_fd_sc_hd__buf_12_45/A sky130_fd_sc_hd__buf_6_17/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_332 vccd1 vssd1 sky130_fd_sc_hd__and3_4_16/X sky130_fd_sc_hd__or2_0_52/B
+ sky130_fd_sc_hd__or2_0_53/A sky130_fd_sc_hd__nor2_2_19/Y sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__o21ai_1_553/B1 sky130_fd_sc_hd__nor2b_2_3/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_272 vssd1 vccd1 sky130_fd_sc_hd__buf_8_150/A sky130_fd_sc_hd__clkbuf_1_50/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_343 vccd1 vssd1 sky130_fd_sc_hd__and3_4_11/X sky130_fd_sc_hd__buf_2_23/X
+ sky130_fd_sc_hd__buf_2_31/X sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__buf_2_19/X
+ sky130_fd_sc_hd__o21ai_1_569/B1 sky130_fd_sc_hd__and2b_4_8/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_283 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_284/A sky130_fd_sc_hd__buf_12_64/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_354 vccd1 vssd1 sky130_fd_sc_hd__and3_4_11/X sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__buf_4_7/X sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__buf_4_0/X
+ sky130_fd_sc_hd__o21ai_1_586/B1 sky130_fd_sc_hd__and2b_4_8/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_294 vssd1 vccd1 sky130_fd_sc_hd__buf_8_155/A sky130_fd_sc_hd__clkbuf_1_294/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_365 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__buf_4_7/X sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__buf_4_0/X
+ sky130_fd_sc_hd__o21ai_1_605/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_376 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__buf_8_0/X sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__o21ai_1_621/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_387 vccd1 vssd1 sky130_fd_sc_hd__and3_4_18/X sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__buf_4_3/X sky130_fd_sc_hd__nor2_2_32/Y sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__o21ai_1_648/B1 sky130_fd_sc_hd__nor2b_2_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_398 vccd1 vssd1 sky130_fd_sc_hd__and3_4_25/X sky130_fd_sc_hd__buf_2_20/X
+ sky130_fd_sc_hd__buf_2_21/X sky130_fd_sc_hd__nor2_1_186/Y sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__o21ai_1_664/B1 sky130_fd_sc_hd__nor2b_1_17/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__buf_4_0 vccd1 vssd1 sky130_fd_sc_hd__buf_4_0/X sky130_fd_sc_hd__buf_4_0/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__and2_0_270 vccd1 vssd1 sky130_fd_sc_hd__and2_0_270/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__xor2_1_643/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__a21oi_2_11 sky130_fd_sc_hd__a21oi_2_11/B1 sky130_fd_sc_hd__or2_0_35/X
+ sky130_fd_sc_hd__o21ai_2_9/Y sky130_fd_sc_hd__xor2_1_330/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_2
Xsky130_fd_sc_hd__and2_0_281 vccd1 vssd1 sky130_fd_sc_hd__and2_0_281/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__fa_2_416/SUM vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_292 vccd1 vssd1 sky130_fd_sc_hd__and2_0_292/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_13/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_12_507 sky130_fd_sc_hd__buf_12_507/A sky130_fd_sc_hd__buf_12_564/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_518 sky130_fd_sc_hd__buf_12_518/A sky130_fd_sc_hd__buf_12_518/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_529 sky130_fd_sc_hd__buf_12_529/A sky130_fd_sc_hd__buf_12_529/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__inv_4_0 sky130_fd_sc_hd__inv_4_0/Y sky130_fd_sc_hd__inv_4_0/A vccd1
+ vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__nand2_1_108 sky130_fd_sc_hd__o21ai_1_82/B1 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__xor2_1_330/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_707 sky130_fd_sc_hd__a221oi_1_0/A1 sky130_fd_sc_hd__ha_2_6/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_119 sky130_fd_sc_hd__nand2_1_119/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__xnor2_1_98/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_718 sky130_fd_sc_hd__nor2b_1_97/A sky130_fd_sc_hd__xnor2_1_292/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_729 sky130_fd_sc_hd__nor2b_1_108/A sky130_fd_sc_hd__xor2_1_683/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__or2_0_105 sky130_fd_sc_hd__or2_0_105/A sky130_fd_sc_hd__or2_0_105/X
+ sky130_fd_sc_hd__or2_0_105/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__o21ai_1_260 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_295/A2 sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__o21ai_1_260/B1 sky130_fd_sc_hd__xor2_1_84/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_271 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_2/X sky130_fd_sc_hd__nand2_1_214/Y
+ sky130_fd_sc_hd__a21oi_1_47/Y sky130_fd_sc_hd__xnor2_1_24/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_282 vssd1 vccd1 sky130_fd_sc_hd__buf_2_3/X sky130_fd_sc_hd__nand2b_1_6/Y
+ sky130_fd_sc_hd__o21ai_1_282/B1 sky130_fd_sc_hd__xor2_1_102/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_293 vssd1 vccd1 sky130_fd_sc_hd__buf_2_2/X sky130_fd_sc_hd__nand2b_1_6/Y
+ sky130_fd_sc_hd__o21ai_1_293/B1 sky130_fd_sc_hd__xor2_1_114/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_703 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_714 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_725 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_736 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_620 sky130_fd_sc_hd__nand2_1_620/Y sky130_fd_sc_hd__buf_2_20/X
+ sky130_fd_sc_hd__buf_2_4/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_747 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_631 sky130_fd_sc_hd__xor2_1_616/A sky130_fd_sc_hd__nand2_1_632/Y
+ sky130_fd_sc_hd__nand2_1_631/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_758 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_642 sky130_fd_sc_hd__nand2_1_642/Y sky130_fd_sc_hd__or2_0_69/A
+ sky130_fd_sc_hd__or2_0_69/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_769 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_653 sky130_fd_sc_hd__nand2_1_653/Y sky130_fd_sc_hd__buf_2_29/X
+ sky130_fd_sc_hd__or2_0_71/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_664 sky130_fd_sc_hd__xor2_1_640/B sky130_fd_sc_hd__nand2_1_665/Y
+ sky130_fd_sc_hd__nand2_1_664/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_2_0 la_data_in[1] la_oenb[1] sky130_fd_sc_hd__nor2b_2_0/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_2
Xsky130_fd_sc_hd__nand2_1_675 sky130_fd_sc_hd__nand2_1_675/Y sky130_fd_sc_hd__or2_0_76/A
+ sky130_fd_sc_hd__or2_0_76/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_686 sky130_fd_sc_hd__xnor2_1_194/A sky130_fd_sc_hd__nand2_1_687/Y
+ sky130_fd_sc_hd__or2_0_78/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_697 sky130_fd_sc_hd__nand2_1_697/Y sky130_fd_sc_hd__mux2_4_2/X
+ sky130_fd_sc_hd__mux2_2_48/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_1702 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1713 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_12 sky130_fd_sc_hd__inv_2_12/A sky130_fd_sc_hd__inv_2_12/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1724 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_23 sky130_fd_sc_hd__inv_2_23/A sky130_fd_sc_hd__inv_2_23/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1735 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_34 sky130_fd_sc_hd__inv_2_34/A sky130_fd_sc_hd__inv_2_34/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1746 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_45 sky130_fd_sc_hd__inv_2_45/A sky130_fd_sc_hd__inv_2_45/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1757 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_56 sky130_fd_sc_hd__inv_2_56/A sky130_fd_sc_hd__inv_2_56/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_460 sky130_fd_sc_hd__buf_2_63/A sky130_fd_sc_hd__clkinv_2_46/Y
+ sky130_fd_sc_hd__nand2_1_845/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1768 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_67 sky130_fd_sc_hd__inv_2_67/A sky130_fd_sc_hd__inv_2_67/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_471 sky130_fd_sc_hd__nor2_1_277/B sky130_fd_sc_hd__edfxbp_1_0/CLK
+ sky130_fd_sc_hd__nor2b_1_122/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1779 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_78 sky130_fd_sc_hd__inv_2_79/A sky130_fd_sc_hd__inv_2_78/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_482 sky130_fd_sc_hd__ha_2_39/A sky130_fd_sc_hd__dfxtp_1_489/CLK
+ sky130_fd_sc_hd__and2_0_367/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_2_2 sky130_fd_sc_hd__nand2_2_2/Y sky130_fd_sc_hd__nand2_2_2/A
+ sky130_fd_sc_hd__nand2_2_2/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__inv_2_89 sky130_fd_sc_hd__inv_2_89/A sky130_fd_sc_hd__inv_2_89/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_493 la_data_out[42] sky130_fd_sc_hd__dfxtp_1_498/CLK sky130_fd_sc_hd__and2_0_378/X
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2b_1_30 sky130_fd_sc_hd__inv_2_152/A sky130_fd_sc_hd__dfxtp_1_1/Q
+ sky130_fd_sc_hd__dfxtp_1_20/Q vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a222oi_1_140 vccd1 vssd1 sky130_fd_sc_hd__and3_4_2/X sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__nor2_2_10/B sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__buf_6_4/X
+ sky130_fd_sc_hd__o21ai_1_285/B1 sky130_fd_sc_hd__and2b_4_4/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_151 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__nor2_2_10/B
+ sky130_fd_sc_hd__buf_6_4/X sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__o21ai_1_297/B1 sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_162 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__nor2_2_10/B sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__buf_6_4/X
+ sky130_fd_sc_hd__o21ai_1_312/B1 sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_310 sky130_fd_sc_hd__fa_2_301/CIN sky130_fd_sc_hd__fa_2_312/A
+ sky130_fd_sc_hd__fa_2_310/A sky130_fd_sc_hd__fa_2_310/B sky130_fd_sc_hd__xor2_1_474/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_173 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__nor2_2_10/B
+ sky130_fd_sc_hd__buf_6_4/X sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__o21ai_1_325/B1 sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_321 sky130_fd_sc_hd__fa_2_314/A sky130_fd_sc_hd__fa_2_322/B
+ sky130_fd_sc_hd__fa_2_321/A sky130_fd_sc_hd__fa_2_321/B sky130_fd_sc_hd__xor2_1_483/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_184 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__nor2_2_4/B
+ sky130_fd_sc_hd__buf_2_4/A sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__o21ai_1_342/B1 sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_332 sky130_fd_sc_hd__fa_2_324/A sky130_fd_sc_hd__fa_2_326/A
+ sky130_fd_sc_hd__fa_2_332/A sky130_fd_sc_hd__fa_2_332/B sky130_fd_sc_hd__xor2_1_497/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_195 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__nor2_2_5/A
+ sky130_fd_sc_hd__nor2_2_5/B sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__nor2_2_4/B
+ sky130_fd_sc_hd__o21ai_1_359/B1 sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_343 sky130_fd_sc_hd__fa_2_336/CIN sky130_fd_sc_hd__fa_2_342/A
+ sky130_fd_sc_hd__fa_2_343/A sky130_fd_sc_hd__fa_2_343/B sky130_fd_sc_hd__xor2_1_515/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_354 sky130_fd_sc_hd__fa_2_346/B sky130_fd_sc_hd__fa_2_351/A
+ sky130_fd_sc_hd__fa_2_354/A sky130_fd_sc_hd__fa_2_354/B sky130_fd_sc_hd__fa_2_354/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_365 sky130_fd_sc_hd__fa_2_359/A sky130_fd_sc_hd__fa_2_366/A
+ sky130_fd_sc_hd__fa_2_365/A sky130_fd_sc_hd__fa_2_365/B sky130_fd_sc_hd__xor2_1_536/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_376 sky130_fd_sc_hd__fa_2_370/A sky130_fd_sc_hd__fa_2_375/B
+ sky130_fd_sc_hd__fa_2_376/A sky130_fd_sc_hd__fa_2_376/B sky130_fd_sc_hd__fa_2_376/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_17 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_4_1/Y
+ sky130_fd_sc_hd__dfxtp_1_170/CLK sky130_fd_sc_hd__o21ai_2_1/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_387 sky130_fd_sc_hd__nor2_2_27/A sky130_fd_sc_hd__or2_1_3/B
+ sky130_fd_sc_hd__fa_2_387/A sky130_fd_sc_hd__fa_2_387/B sky130_fd_sc_hd__fa_2_387/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_28 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_8_5/Y
+ sky130_fd_sc_hd__dfxtp_1_269/CLK sky130_fd_sc_hd__o21ai_2_4/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_398 sky130_fd_sc_hd__fa_2_397/A sky130_fd_sc_hd__fah_1_8/A
+ sky130_fd_sc_hd__fa_2_398/A sky130_fd_sc_hd__fa_2_398/B sky130_fd_sc_hd__fa_2_398/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_39 sky130_fd_sc_hd__conb_1_145/LO sky130_fd_sc_hd__clkinv_4_11/Y
+ sky130_fd_sc_hd__dfxtp_1_371/CLK sky130_fd_sc_hd__o21ai_1_892/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__clkinv_8_70 sky130_fd_sc_hd__clkinv_8_71/A sky130_fd_sc_hd__clkinv_8_70/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_81 sky130_fd_sc_hd__clkinv_8_82/A sky130_fd_sc_hd__clkinv_8_81/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_90 sky130_fd_sc_hd__buf_8_95/X sky130_fd_sc_hd__buf_12_90/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__nor2_1_108 sky130_fd_sc_hd__nor2_1_113/B sky130_fd_sc_hd__nor2_1_108/Y
+ sky130_fd_sc_hd__nor2_1_108/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_119 sky130_fd_sc_hd__nor2_1_119/B sky130_fd_sc_hd__nor2_1_119/Y
+ sky130_fd_sc_hd__nor2_1_119/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_17 sky130_fd_sc_hd__nor2_4_0/Y sky130_fd_sc_hd__nor2_2_0/Y
+ sky130_fd_sc_hd__dfxtp_1_332/Q sky130_fd_sc_hd__or2_0_88/A sky130_fd_sc_hd__nand2_1_14/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_28 sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__dfxtp_1_277/Q sky130_fd_sc_hd__o211ai_1_1/Y sky130_fd_sc_hd__nand2_2_6/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_39 sky130_fd_sc_hd__clkbuf_1_24/X sky130_fd_sc_hd__clkbuf_1_23/X
+ sky130_fd_sc_hd__dfxtp_1_98/Q sky130_fd_sc_hd__dfxtp_1_66/Q sky130_fd_sc_hd__a22oi_1_39/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_304 sky130_fd_sc_hd__buf_12_85/X sky130_fd_sc_hd__buf_12_475/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_315 sky130_fd_sc_hd__buf_12_315/A sky130_fd_sc_hd__buf_12_544/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_326 sky130_fd_sc_hd__buf_12_326/A sky130_fd_sc_hd__buf_12_478/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_337 sky130_fd_sc_hd__buf_12_337/A sky130_fd_sc_hd__buf_12_601/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_348 sky130_fd_sc_hd__buf_12_348/A sky130_fd_sc_hd__buf_12_492/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_207 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__nor2b_2_3/Y sky130_fd_sc_hd__nor2_2_19/Y sky130_fd_sc_hd__a22oi_1_207/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_359 sky130_fd_sc_hd__buf_12_359/A sky130_fd_sc_hd__buf_12_669/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_218 sky130_fd_sc_hd__or2_0_72/B sky130_fd_sc_hd__or2_0_72/A
+ sky130_fd_sc_hd__nor2b_1_12/Y sky130_fd_sc_hd__nor2_2_31/Y sky130_fd_sc_hd__a22oi_1_218/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_504 sky130_fd_sc_hd__nand2_1_477/A sky130_fd_sc_hd__nor2_1_160/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_515 sky130_fd_sc_hd__xnor2_2_2/A sky130_fd_sc_hd__nand2_1_503/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_526 sky130_fd_sc_hd__o21ai_1_671/A2 sky130_fd_sc_hd__xnor2_1_135/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_537 sky130_fd_sc_hd__nand2_1_531/A sky130_fd_sc_hd__nor2_1_173/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_548 sky130_fd_sc_hd__nor2_1_176/A sky130_fd_sc_hd__nand2_1_554/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_559 sky130_fd_sc_hd__o21ai_1_752/B1 sky130_fd_sc_hd__o21ai_1_753/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_40 sky130_fd_sc_hd__ha_2_9/SUM sky130_fd_sc_hd__nor2_1_40/Y
+ sky130_fd_sc_hd__nor2_1_40/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_51 sky130_fd_sc_hd__nor2_1_51/B sky130_fd_sc_hd__nor2_1_51/Y
+ sky130_fd_sc_hd__nor2_1_55/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_62 sky130_fd_sc_hd__nor2_1_62/B sky130_fd_sc_hd__nor2_1_62/Y
+ sky130_fd_sc_hd__nor2_1_62/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_17 sky130_fd_sc_hd__a21o_2_1/X sky130_fd_sc_hd__inv_2_126/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_73 sky130_fd_sc_hd__nor2_1_73/B sky130_fd_sc_hd__nor2_1_73/Y
+ sky130_fd_sc_hd__buf_6_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_28 sky130_fd_sc_hd__nand2_1_9/Y sky130_fd_sc_hd__clkinv_4_28/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_84 sky130_fd_sc_hd__nor2_1_90/Y sky130_fd_sc_hd__nor2_1_84/Y
+ sky130_fd_sc_hd__nor2_1_87/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_39 sky130_fd_sc_hd__clkinv_8_72/A sky130_fd_sc_hd__clkinv_4_40/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_95 sky130_fd_sc_hd__nor2_2_4/B sky130_fd_sc_hd__nor2_1_95/Y
+ sky130_fd_sc_hd__buf_2_4/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_12_1009 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21a_1_5 sky130_fd_sc_hd__o21a_1_5/X sky130_fd_sc_hd__o21a_1_5/A1
+ sky130_fd_sc_hd__o21a_1_5/B1 sky130_fd_sc_hd__o21a_1_5/A2 vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__decap_12_500 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_511 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_522 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_533 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_544 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_555 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_566 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_450 sky130_fd_sc_hd__xnor2_1_113/A sky130_fd_sc_hd__nand2_1_451/Y
+ sky130_fd_sc_hd__nand2_1_450/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_577 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_461 sky130_fd_sc_hd__nand2_1_461/Y sky130_fd_sc_hd__nor2_1_155/A
+ sky130_fd_sc_hd__nor2_1_155/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_588 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_472 sky130_fd_sc_hd__nand2_1_472/Y sky130_fd_sc_hd__nand2_1_482/Y
+ sky130_fd_sc_hd__nand2_1_478/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_599 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_483 sky130_fd_sc_hd__nand2_1_483/Y sky130_fd_sc_hd__xnor2_1_67/B
+ sky130_fd_sc_hd__nand2_1_487/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_494 sky130_fd_sc_hd__nand2_1_494/Y sky130_fd_sc_hd__nor2_1_178/Y
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_30 sky130_fd_sc_hd__fa_2_417/B sky130_fd_sc_hd__fa_2_465/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_41 sky130_fd_sc_hd__or2_0_74/B sky130_fd_sc_hd__nor2b_1_41/Y
+ sky130_fd_sc_hd__buf_2_214/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_52 sky130_fd_sc_hd__or2_1_11/A sky130_fd_sc_hd__fa_2_477/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_63 sky130_fd_sc_hd__mux2_2_24/X sky130_fd_sc_hd__nor2b_1_63/Y
+ sky130_fd_sc_hd__mux2_4_5/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1030 sky130_fd_sc_hd__clkinv_1_1031/A sky130_fd_sc_hd__inv_2_86/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_74 sky130_fd_sc_hd__xnor2_2_5/A sky130_fd_sc_hd__fa_2_488/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1041 sky130_fd_sc_hd__buf_8_112/A sky130_fd_sc_hd__inv_2_168/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_85 sky130_fd_sc_hd__or2_0_84/A sky130_fd_sc_hd__nor2b_1_85/Y
+ sky130_fd_sc_hd__mux2_4_5/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1052 sky130_fd_sc_hd__inv_2_185/A sky130_fd_sc_hd__ha_2_34/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1510 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_96 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_96/Y
+ sky130_fd_sc_hd__nor2b_1_96/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1063 sky130_fd_sc_hd__bufinv_8_1/A sky130_fd_sc_hd__buf_8_129/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_4 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_4/B sky130_fd_sc_hd__buf_2_2/A
+ sky130_fd_sc_hd__xnor2_1_4/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_1521 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1074 sky130_fd_sc_hd__nor2_1_278/B sky130_fd_sc_hd__nor2_4_0/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1532 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1085 sky130_fd_sc_hd__maj3_1_2/C sky130_fd_sc_hd__ha_2_59/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1543 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1096 sky130_fd_sc_hd__and2_0_361/A sky130_fd_sc_hd__inv_2_107/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1554 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1565 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1576 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1587 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_290 sky130_fd_sc_hd__a22oi_1_2/B2 sky130_fd_sc_hd__dfxtp_1_2/CLK
+ sky130_fd_sc_hd__and2_0_266/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1598 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__mux2_4_0 sky130_fd_sc_hd__or2_0_82/B sky130_fd_sc_hd__mux2_8_1/S
+ sky130_fd_sc_hd__buf_6_12/X sky130_fd_sc_hd__mux2_4_0/A1 vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__mux2_4
Xsky130_fd_sc_hd__fa_2_140 sky130_fd_sc_hd__fa_2_139/B sky130_fd_sc_hd__or2_0_22/A
+ sky130_fd_sc_hd__fa_2_140/A sky130_fd_sc_hd__fa_2_140/B sky130_fd_sc_hd__fa_2_140/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_151 sky130_fd_sc_hd__fa_2_150/B sky130_fd_sc_hd__fa_2_152/CIN
+ sky130_fd_sc_hd__fa_2_151/A sky130_fd_sc_hd__fa_2_151/B sky130_fd_sc_hd__xor2_1_235/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_162 sky130_fd_sc_hd__fa_2_158/B sky130_fd_sc_hd__fa_2_168/B
+ sky130_fd_sc_hd__fa_2_162/A sky130_fd_sc_hd__fa_2_162/B sky130_fd_sc_hd__xor2_1_245/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and3_4_1 sky130_fd_sc_hd__nor2_2_9/B sky130_fd_sc_hd__nor2_2_9/A
+ sky130_fd_sc_hd__and3_4_1/C sky130_fd_sc_hd__and3_4_1/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__dfxtp_1_19 sky130_fd_sc_hd__buf_2_189/A sky130_fd_sc_hd__edfxbp_1_0/CLK
+ la_data_out[35] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_173 sky130_fd_sc_hd__fa_2_166/A sky130_fd_sc_hd__fa_2_174/B
+ sky130_fd_sc_hd__fa_2_173/A sky130_fd_sc_hd__fa_2_173/B sky130_fd_sc_hd__xor2_1_264/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_184 sky130_fd_sc_hd__fa_2_177/A sky130_fd_sc_hd__fa_2_185/A
+ sky130_fd_sc_hd__fa_2_184/A sky130_fd_sc_hd__fa_2_184/B sky130_fd_sc_hd__fa_2_184/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_195 sky130_fd_sc_hd__fa_2_188/CIN sky130_fd_sc_hd__fa_2_194/A
+ sky130_fd_sc_hd__fa_2_195/A sky130_fd_sc_hd__fa_2_195/B sky130_fd_sc_hd__xor2_1_293/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o22ai_1_50 sky130_fd_sc_hd__nor2_1_17/A sky130_fd_sc_hd__o22ai_1_50/B1
+ sky130_fd_sc_hd__o22ai_1_50/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_61 sky130_fd_sc_hd__nor2_1_4/A sky130_fd_sc_hd__o22ai_1_0/A2
+ sky130_fd_sc_hd__o22ai_1_61/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_72 sky130_fd_sc_hd__xnor2_2_6/Y sky130_fd_sc_hd__xnor2_1_227/Y
+ sky130_fd_sc_hd__o22ai_1_72/Y sky130_fd_sc_hd__xnor2_1_223/Y sky130_fd_sc_hd__o22ai_1_98/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_190 vccd1 vssd1 sky130_fd_sc_hd__ha_2_9/A sky130_fd_sc_hd__or4_1_1/B
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_83 sky130_fd_sc_hd__xnor2_1_233/Y sky130_fd_sc_hd__xnor2_1_241/Y
+ sky130_fd_sc_hd__fa_2_440/B sky130_fd_sc_hd__inv_2_65/Y sky130_fd_sc_hd__o22ai_1_99/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_94 sky130_fd_sc_hd__xnor2_1_241/Y sky130_fd_sc_hd__xnor2_1_245/Y
+ sky130_fd_sc_hd__ha_2_13/B sky130_fd_sc_hd__inv_2_65/Y sky130_fd_sc_hd__o22ai_1_99/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_4_30 vccd1 vssd1 sky130_fd_sc_hd__buf_4_30/X sky130_fd_sc_hd__buf_4_30/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_41 vccd1 vssd1 sky130_fd_sc_hd__buf_4_41/X sky130_fd_sc_hd__buf_4_41/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_12_101 sky130_fd_sc_hd__buf_8_150/X sky130_fd_sc_hd__buf_12_101/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_112 sky130_fd_sc_hd__buf_8_4/X sky130_fd_sc_hd__buf_12_112/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_sram_1kbyte_1rw1r_32x256_8_9 sky130_fd_sc_hd__buf_2_143/X sky130_fd_sc_hd__buf_2_143/X
+ sky130_fd_sc_hd__buf_12_676/X sky130_fd_sc_hd__buf_12_634/X sky130_fd_sc_hd__buf_12_443/X
+ sky130_fd_sc_hd__buf_12_675/X sky130_fd_sc_hd__buf_12_669/X sky130_fd_sc_hd__buf_12_642/X
+ sky130_fd_sc_hd__buf_12_616/X sky130_fd_sc_hd__nand2b_2_10/Y sky130_fd_sc_hd__buf_12_638/X
+ sky130_fd_sc_hd__buf_12_593/X sky130_fd_sc_hd__buf_12_633/X vccd1 sky130_fd_sc_hd__clkinv_2_45/Y
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[16] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[17]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[18] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[19]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[20] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[21]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[22] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[23]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[24] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[25]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[26] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[27]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[28] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[29]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[30] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[31]
+ sky130_fd_sc_hd__buf_12_527/X sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[1] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[2]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[3] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[4]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[5] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[6]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[7] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[8]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[9] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[10]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[11] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[12]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[13] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[14]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[15] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout1[0]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[10] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[11]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[12] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[13]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[14] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[15]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[16] sky130_fd_sc_hd__buf_12_553/X sky130_fd_sc_hd__buf_12_100/X
+ sky130_fd_sc_hd__buf_12_95/X sky130_fd_sc_hd__buf_12_162/X sky130_fd_sc_hd__buf_12_161/X
+ sky130_fd_sc_hd__dfxtp_1_0/CLK sky130_fd_sc_hd__buf_2_140/X sky130_fd_sc_hd__buf_2_140/X
+ sky130_fd_sc_hd__buf_2_140/X sky130_fd_sc_hd__buf_2_140/A sky130_fd_sc_hd__buf_2_140/A
+ sky130_fd_sc_hd__buf_2_140/A sky130_fd_sc_hd__buf_2_140/A sky130_fd_sc_hd__buf_2_140/A
+ sky130_fd_sc_hd__buf_2_140/A sky130_fd_sc_hd__buf_2_140/A sky130_fd_sc_hd__buf_2_140/A
+ sky130_fd_sc_hd__buf_2_140/A sky130_fd_sc_hd__buf_2_140/A sky130_fd_sc_hd__buf_2_140/A
+ sky130_fd_sc_hd__buf_2_140/A sky130_fd_sc_hd__buf_2_140/A sky130_fd_sc_hd__buf_2_140/A
+ sky130_fd_sc_hd__buf_2_140/A sky130_fd_sc_hd__buf_2_140/A sky130_fd_sc_hd__buf_2_140/A
+ sky130_fd_sc_hd__buf_6_7/A sky130_fd_sc_hd__buf_6_7/A sky130_fd_sc_hd__buf_6_7/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[0] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[1]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[2] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[3]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[4] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[5]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[6] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[7]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[8] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[9]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[25] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[26]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[27] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[28]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[29] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[30]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[31] sky130_fd_sc_hd__buf_6_7/A sky130_fd_sc_hd__buf_6_7/A
+ sky130_fd_sc_hd__buf_6_7/A sky130_fd_sc_hd__buf_6_7/A sky130_fd_sc_hd__buf_6_7/A
+ sky130_fd_sc_hd__buf_6_7/A sky130_fd_sc_hd__buf_6_7/A sky130_fd_sc_hd__buf_6_7/A
+ sky130_fd_sc_hd__buf_6_7/A sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[17] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[18]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[19] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[20]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[21] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[22]
+ sky130_fd_sc_hd__buf_8_165/X sky130_fd_sc_hd__buf_12_619/X sky130_fd_sc_hd__buf_12_607/X
+ sky130_fd_sc_hd__buf_12_519/X sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[23] sky130_sram_1kbyte_1rw1r_32x256_8_9/dout0[24]
+ sky130_sram_1kbyte_1rw1r_32x256_8_9/sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/gnd_uq26
+ vssd1 sky130_sram_1kbyte_1rw1r_32x256_8
Xsky130_fd_sc_hd__buf_12_123 sky130_fd_sc_hd__buf_8_40/X sky130_fd_sc_hd__buf_12_123/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_134 sky130_fd_sc_hd__buf_8_45/X sky130_fd_sc_hd__buf_12_402/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_145 sky130_fd_sc_hd__buf_12_30/X sky130_fd_sc_hd__buf_12_439/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_156 sky130_fd_sc_hd__buf_12_56/X sky130_fd_sc_hd__buf_12_310/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_167 sky130_fd_sc_hd__buf_12_16/X sky130_fd_sc_hd__buf_12_167/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_90 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_44/A1 sky130_fd_sc_hd__clkbuf_1_90/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_4_4 sky130_fd_sc_hd__nor2_2_5/A sky130_fd_sc_hd__buf_4_0/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_12_178 sky130_fd_sc_hd__buf_8_105/X sky130_fd_sc_hd__buf_12_278/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_189 sky130_fd_sc_hd__buf_4_31/X sky130_fd_sc_hd__buf_12_443/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_301 sky130_fd_sc_hd__and2_0_248/A sky130_fd_sc_hd__a222oi_1_45/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_312 sky130_fd_sc_hd__a21oi_1_35/B1 sky130_fd_sc_hd__nand2_1_168/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_323 sky130_fd_sc_hd__a21oi_2_0/B1 sky130_fd_sc_hd__nand2_1_180/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_334 sky130_fd_sc_hd__nand2_1_195/A sky130_fd_sc_hd__nor2_1_58/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_345 sky130_fd_sc_hd__nand2_1_206/A sky130_fd_sc_hd__nor2_1_62/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_356 sky130_fd_sc_hd__nor2_1_66/A sky130_fd_sc_hd__nand2_1_231/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_367 sky130_fd_sc_hd__nand2_1_246/A sky130_fd_sc_hd__nor2_1_77/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_378 sky130_fd_sc_hd__a21oi_1_58/B1 sky130_fd_sc_hd__nand2_1_274/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_389 sky130_fd_sc_hd__nand2_1_285/A sky130_fd_sc_hd__nor2_1_97/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_2_8 sky130_fd_sc_hd__a21oi_2_8/B1 sky130_fd_sc_hd__or2_0_29/X
+ sky130_fd_sc_hd__xnor2_1_78/B sky130_fd_sc_hd__a21oi_2_8/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_2
Xsky130_fd_sc_hd__or2_0_70 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__or2_0_70/X
+ sky130_fd_sc_hd__or2_0_70/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__clkinv_4_4 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkinv_4_4/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__or2_0_81 sky130_fd_sc_hd__or2_0_81/A sky130_fd_sc_hd__or2_0_81/X
+ la_data_out[71] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_92 sky130_fd_sc_hd__or2_0_92/A sky130_fd_sc_hd__or2_0_92/X
+ sky130_fd_sc_hd__or2_0_92/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__decap_12_330 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_341 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_352 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_363 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_374 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_385 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_396 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_280 sky130_fd_sc_hd__nand2_1_280/Y sky130_fd_sc_hd__nor2_1_94/A
+ sky130_fd_sc_hd__nor2_1_94/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_108 sky130_fd_sc_hd__xor2_1_9/B sky130_fd_sc_hd__fa_2_79/A
+ sky130_fd_sc_hd__xor2_1_108/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_291 sky130_fd_sc_hd__xnor2_1_1/B sky130_fd_sc_hd__nand2_1_292/Y
+ sky130_fd_sc_hd__nand2_1_291/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_890 sky130_fd_sc_hd__clkinv_1_890/Y sky130_fd_sc_hd__clkinv_4_88/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xor2_1_119 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__fa_2_88/B
+ sky130_fd_sc_hd__xor2_1_119/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1340 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1351 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_90 sky130_fd_sc_hd__conb_1_90/LO sky130_fd_sc_hd__conb_1_90/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1362 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1373 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_804 vssd1 vccd1 sky130_fd_sc_hd__inv_2_52/Y sky130_fd_sc_hd__nand2_1_594/Y
+ sky130_fd_sc_hd__a21oi_1_122/Y sky130_fd_sc_hd__xnor2_1_165/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1384 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_815 vssd1 vccd1 sky130_fd_sc_hd__nand2_2_13/Y sky130_fd_sc_hd__nand2b_1_16/Y
+ sky130_fd_sc_hd__a22oi_1_220/Y sky130_fd_sc_hd__xor2_1_590/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1395 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_826 vssd1 vccd1 sky130_fd_sc_hd__inv_2_48/Y sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__o21ai_1_826/B1 sky130_fd_sc_hd__xor2_1_600/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_837 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_9/X sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_837/B1 sky130_fd_sc_hd__xor2_1_610/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_848 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_861/A2 sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__nand2_1_500/Y sky130_fd_sc_hd__xor2_1_621/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_859 vssd1 vccd1 sky130_fd_sc_hd__buf_2_13/X sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_859/B1 sky130_fd_sc_hd__xor2_1_633/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nand2b_2_5 sky130_fd_sc_hd__nor2_4_14/B sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__nor2_4_14/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_2
Xsky130_fd_sc_hd__xor2_1_620 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__fa_2_411/B
+ sky130_fd_sc_hd__xor2_1_620/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_631 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__nor2_4_18/B
+ sky130_fd_sc_hd__xor2_1_631/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_642 sky130_fd_sc_hd__xor2_1_642/B sky130_fd_sc_hd__xor2_1_642/X
+ sky130_fd_sc_hd__xor2_1_642/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_653 sky130_fd_sc_hd__xor2_1_653/B sky130_fd_sc_hd__xor2_1_653/X
+ sky130_fd_sc_hd__xor2_1_653/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_664 sky130_fd_sc_hd__xor2_1_664/B sky130_fd_sc_hd__xor2_1_664/X
+ sky130_fd_sc_hd__xor2_1_664/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_675 sky130_fd_sc_hd__xor2_1_675/B sky130_fd_sc_hd__xor2_1_675/X
+ sky130_fd_sc_hd__xor2_1_675/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_686 sky130_fd_sc_hd__xor2_1_686/B sky130_fd_sc_hd__xor2_1_686/X
+ sky130_fd_sc_hd__xor2_1_686/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_697 sky130_fd_sc_hd__a21o_2_4/B1 sky130_fd_sc_hd__xor2_1_697/X
+ wbs_adr_i[10] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkinv_1_18 la_data_out[109] sky130_fd_sc_hd__conb_1_124/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_29 la_data_out[98] sky130_fd_sc_hd__conb_1_113/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__fa_2_5 sky130_fd_sc_hd__xor3_1_0/B sky130_fd_sc_hd__fa_2_5/SUM sky130_fd_sc_hd__fa_2_5/A
+ sky130_fd_sc_hd__fa_2_5/B sky130_fd_sc_hd__fa_2_5/CIN vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a211o_1_11 vssd1 vccd1 sky130_fd_sc_hd__fa_2_265/A sky130_fd_sc_hd__dfxtp_1_74/Q
+ sky130_fd_sc_hd__nor2_1_15/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_11/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__a211o_1_22 vssd1 vccd1 sky130_fd_sc_hd__fa_2_214/A sky130_fd_sc_hd__dfxtp_1_85/Q
+ sky130_fd_sc_hd__nor2_1_26/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_22/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__clkinv_1_120 io_oeb[19] sky130_fd_sc_hd__conb_1_22/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_131 io_oeb[8] sky130_fd_sc_hd__conb_1_11/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_142 user_irq[0] sky130_fd_sc_hd__conb_1_0/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_153 sky130_fd_sc_hd__o21ai_1_2/A2 sky130_fd_sc_hd__dfxtp_1_124/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_164 sky130_fd_sc_hd__nor2_1_30/A sky130_fd_sc_hd__dfxtp_1_153/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_175 sky130_fd_sc_hd__o22ai_1_40/B1 sky130_fd_sc_hd__dfxtp_1_182/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_7 sky130_fd_sc_hd__buf_8_7/A sky130_fd_sc_hd__buf_8_7/X vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__a22o_1_9 sky130_fd_sc_hd__inv_2_66/Y sky130_fd_sc_hd__or2_0_92/B
+ sky130_fd_sc_hd__a22o_1_9/X sky130_fd_sc_hd__a22o_1_9/B2 sky130_fd_sc_hd__a22o_1_9/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_186 sky130_fd_sc_hd__o22ai_1_20/B1 sky130_fd_sc_hd__dfxtp_1_115/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_11 sky130_fd_sc_hd__inv_2_66/Y sky130_fd_sc_hd__or2_0_91/B
+ sky130_fd_sc_hd__a22o_1_11/X sky130_fd_sc_hd__a22o_1_9/B2 sky130_fd_sc_hd__a22o_1_11/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_22 sky130_fd_sc_hd__buf_2_63/A sky130_fd_sc_hd__buf_2_97/X
+ sky130_fd_sc_hd__a22o_1_22/X sky130_fd_sc_hd__a22o_1_22/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_197 sky130_fd_sc_hd__nor2_1_20/A sky130_fd_sc_hd__dfxtp_1_143/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_33 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__buf_2_108/X
+ sky130_fd_sc_hd__a22o_1_33/X sky130_fd_sc_hd__a22o_1_33/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_44 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__buf_2_119/X
+ sky130_fd_sc_hd__a22o_1_44/X sky130_fd_sc_hd__a22o_1_44/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_55 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__buf_2_46/A
+ sky130_fd_sc_hd__a22o_1_55/X sky130_fd_sc_hd__ha_2_26/SUM sky130_fd_sc_hd__a22o_1_71/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_66 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__clkbuf_4_8/A
+ sky130_fd_sc_hd__a22o_1_66/X sky130_fd_sc_hd__ha_2_35/SUM sky130_fd_sc_hd__a22o_1_71/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_77 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__buf_4_38/X
+ sky130_fd_sc_hd__a22o_1_77/X sky130_fd_sc_hd__ha_2_23/SUM sky130_fd_sc_hd__nor2_1_269/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_2_1 sky130_fd_sc_hd__clkinv_2_1/Y sky130_fd_sc_hd__clkinv_2_1/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__nor2_1_280 sky130_fd_sc_hd__maj3_1_3/X sky130_fd_sc_hd__nor2_1_280/Y
+ sky130_fd_sc_hd__ha_2_55/SUM vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_12_160 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_171 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_182 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_12 sky130_fd_sc_hd__nand2_1_12/Y sky130_fd_sc_hd__nand2_1_12/B
+ sky130_fd_sc_hd__nand2_1_12/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_193 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_23 sky130_fd_sc_hd__nand2_8_2/A sky130_fd_sc_hd__nand2_1_7/B
+ sky130_fd_sc_hd__or2_0_78/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_34 sky130_fd_sc_hd__nand2_1_0/B sky130_fd_sc_hd__nand2_1_8/B
+ sky130_fd_sc_hd__or2_1_10/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_45 sky130_fd_sc_hd__nand2_1_45/Y sky130_fd_sc_hd__nand2_1_8/B
+ sky130_fd_sc_hd__mux2_4_4/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_250 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_4/B sky130_fd_sc_hd__xnor2_1_250/Y
+ sky130_fd_sc_hd__or2_0_82/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_56 sky130_fd_sc_hd__nand2_1_56/Y sky130_fd_sc_hd__nand2_1_56/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_261 vssd1 vccd1 la_data_out[81] sky130_fd_sc_hd__xnor2_1_261/Y
+ sky130_fd_sc_hd__mux2_4_2/X vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_67 sky130_fd_sc_hd__nand2_1_67/Y sky130_fd_sc_hd__nand2_1_67/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_272 vssd1 vccd1 la_data_out[68] sky130_fd_sc_hd__xnor2_1_272/Y
+ sky130_fd_sc_hd__or2_0_78/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_78 sky130_fd_sc_hd__nand2_1_78/Y sky130_fd_sc_hd__nand2_1_78/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_283 vssd1 vccd1 la_data_out[71] sky130_fd_sc_hd__xnor2_1_283/Y
+ sky130_fd_sc_hd__or2_0_79/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_89 sky130_fd_sc_hd__nand2_1_89/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__xor2_1_234/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_294 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_294/B sky130_fd_sc_hd__xnor2_1_294/Y
+ sky130_fd_sc_hd__xnor2_1_294/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_1170 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_601 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_152/Y sky130_fd_sc_hd__nand2_1_457/Y
+ sky130_fd_sc_hd__nand2_1_451/Y sky130_fd_sc_hd__o21ai_1_601/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1181 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_612 vssd1 vccd1 sky130_fd_sc_hd__buf_2_8/X sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_612/B1 sky130_fd_sc_hd__xor2_1_404/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1192 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_623 vssd1 vccd1 sky130_fd_sc_hd__nand2_2_12/Y sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__a22oi_1_212/Y sky130_fd_sc_hd__xor2_1_415/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_634 vssd1 vccd1 sky130_fd_sc_hd__inv_2_44/Y sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_634/B1 sky130_fd_sc_hd__xor2_1_586/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_645 vssd1 vccd1 sky130_fd_sc_hd__inv_2_50/Y sky130_fd_sc_hd__nand2b_1_15/Y
+ sky130_fd_sc_hd__o21ai_1_645/B1 sky130_fd_sc_hd__xor2_1_432/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_656 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_723/A2 sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__o21ai_1_656/B1 sky130_fd_sc_hd__xor2_1_441/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_667 vssd1 vccd1 sky130_fd_sc_hd__inv_2_48/Y sky130_fd_sc_hd__nand2b_1_19/Y
+ sky130_fd_sc_hd__o21ai_1_667/B1 sky130_fd_sc_hd__xor2_1_450/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_678 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_742/A2 sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__o21ai_1_678/B1 sky130_fd_sc_hd__xor2_1_459/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_689 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_723/A2 sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_689/B1 sky130_fd_sc_hd__xor2_1_469/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_19 sky130_fd_sc_hd__fa_2_12/B sky130_fd_sc_hd__fa_2_22/A sky130_fd_sc_hd__fa_2_19/A
+ sky130_fd_sc_hd__fa_2_19/B sky130_fd_sc_hd__fa_2_19/CIN vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__xor2_1_450 sky130_fd_sc_hd__fa_2_338/A sky130_fd_sc_hd__fa_2_291/A
+ sky130_fd_sc_hd__xor2_1_450/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_461 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__xor2_1_461/X
+ sky130_fd_sc_hd__xor2_1_461/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_472 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__xor2_1_472/X
+ sky130_fd_sc_hd__xor2_1_472/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_483 sky130_fd_sc_hd__xor2_1_548/B sky130_fd_sc_hd__xor2_1_483/X
+ sky130_fd_sc_hd__xor2_1_483/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_494 sky130_fd_sc_hd__fa_2_357/A sky130_fd_sc_hd__fa_2_331/B
+ sky130_fd_sc_hd__xor2_1_494/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a222oi_1_503 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__nor2_2_10/B
+ sky130_fd_sc_hd__buf_6_4/X sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__o21ai_1_797/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_514 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__buf_2_15/X
+ sky130_fd_sc_hd__buf_2_4/A sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__buf_2_20/X
+ sky130_fd_sc_hd__o21ai_1_634/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__dfxtp_4_1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_4_1/D sky130_fd_sc_hd__clkinv_4_6/Y
+ sky130_fd_sc_hd__or2_0_24/A vssd1 vccd1 sky130_fd_sc_hd__dfxtp_4
Xsky130_fd_sc_hd__a222oi_1_525 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__buf_4_0/A
+ sky130_fd_sc_hd__buf_2_27/X sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__buf_2_15/X
+ sky130_fd_sc_hd__o21ai_1_827/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_536 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__buf_8_0/A sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__o21ai_1_845/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_547 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_423/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_455/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_744/A sky130_fd_sc_hd__dfxtp_1_391/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_558 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_412/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_444/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_755/A sky130_fd_sc_hd__dfxtp_1_380/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_569 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_401/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_433/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_766/A sky130_fd_sc_hd__dfxtp_1_369/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nor2b_1_103 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_103/Y
+ sky130_fd_sc_hd__nor2b_1_103/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_114 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_114/Y
+ sky130_fd_sc_hd__nor2b_1_114/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_125 sky130_fd_sc_hd__nor2b_1_125/B_N sky130_fd_sc_hd__nor2b_1_125/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_136 sky130_fd_sc_hd__clkinv_4_55/Y sky130_fd_sc_hd__nor2b_1_136/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_147 sky130_fd_sc_hd__clkinv_4_66/Y sky130_fd_sc_hd__nor2b_1_147/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__fah_1_16 sky130_fd_sc_hd__or2_1_3/A sky130_fd_sc_hd__fah_1_16/B
+ sky130_fd_sc_hd__fah_1_16/A sky130_fd_sc_hd__or2_1_1/B sky130_fd_sc_hd__fah_1_16/CI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__fah_1
Xsky130_fd_sc_hd__buf_6_4 vccd1 vssd1 sky130_fd_sc_hd__buf_6_4/X sky130_fd_sc_hd__buf_6_4/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__clkinv_2_50 sky130_fd_sc_hd__buf_4_42/A wbs_dat_i[20] vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__sdlclkp_4_2 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_2_5/Y
+ sky130_fd_sc_hd__dfxtp_1_51/CLK sky130_fd_sc_hd__o21ai_1_0/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_5 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_5/Y
+ sky130_fd_sc_hd__nor2_1_5/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__dfxtp_1_108 sky130_fd_sc_hd__dfxtp_1_108/Q sky130_fd_sc_hd__dfxtp_1_99/CLK
+ sky130_fd_sc_hd__and2_0_167/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_119 sky130_fd_sc_hd__dfxtp_1_119/Q sky130_fd_sc_hd__dfxtp_1_122/CLK
+ sky130_fd_sc_hd__and2_0_223/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_420 vssd1 vccd1 sky130_fd_sc_hd__inv_2_40/Y sky130_fd_sc_hd__nand2b_1_9/Y
+ sky130_fd_sc_hd__o21ai_1_420/B1 sky130_fd_sc_hd__xor2_1_229/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_431 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_496/A2 sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_431/B1 sky130_fd_sc_hd__xor2_1_238/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_442 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_442/A2 sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_442/B1 sky130_fd_sc_hd__xor2_1_247/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_453 vssd1 vccd1 sky130_fd_sc_hd__inv_2_41/Y sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_453/B1 sky130_fd_sc_hd__xor2_1_257/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_464 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_0/Y sky130_fd_sc_hd__nand2b_2_3/Y
+ sky130_fd_sc_hd__o21ai_1_464/B1 sky130_fd_sc_hd__xor2_1_267/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_475 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_505/A2 sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_475/B1 sky130_fd_sc_hd__xor2_1_277/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_3_2 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__o21ai_1_486 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_486/A2 sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_486/B1 sky130_fd_sc_hd__xor2_1_287/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_497 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_7/X sky130_fd_sc_hd__or2_0_32/B
+ sky130_fd_sc_hd__o21a_1_2/A2 sky130_fd_sc_hd__xnor2_1_85/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_907 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_918 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_802 sky130_fd_sc_hd__xnor2_1_293/A sky130_fd_sc_hd__nand2_1_803/Y
+ sky130_fd_sc_hd__or2_0_102/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_929 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_813 sky130_fd_sc_hd__nand2_1_813/Y sky130_fd_sc_hd__nor2_1_259/A
+ sky130_fd_sc_hd__nor2_1_259/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_824 sky130_fd_sc_hd__xor2_1_684/B sky130_fd_sc_hd__nand2_1_825/Y
+ sky130_fd_sc_hd__nand2_1_824/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_835 sky130_fd_sc_hd__nand2_1_835/Y sky130_fd_sc_hd__or2_0_110/A
+ sky130_fd_sc_hd__or2_0_110/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_846 sky130_fd_sc_hd__nand2_1_846/Y la_data_out[36] la_data_out[56]
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_857 sky130_fd_sc_hd__nor2_1_267/B sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_71/B1 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o21ai_1_13 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_20/B1 sky130_fd_sc_hd__inv_2_53/A
+ sky130_fd_sc_hd__o21ai_1_13/B1 sky130_fd_sc_hd__fa_2_82/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_24 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_9/B1 sky130_fd_sc_hd__nor2_4_4/B
+ sky130_fd_sc_hd__o21ai_1_24/B1 sky130_fd_sc_hd__fa_2_130/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_35 vssd1 vccd1 sky130_fd_sc_hd__inv_2_62/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_85/Y sky130_fd_sc_hd__and2_0_3/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_46 vssd1 vccd1 sky130_fd_sc_hd__inv_2_63/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_90/Y sky130_fd_sc_hd__o21ai_1_46/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_57 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_57/A2 sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__o21ai_1_57/B1 sky130_fd_sc_hd__o21ai_1_57/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_280 sky130_fd_sc_hd__fa_2_239/A sky130_fd_sc_hd__xor2_1_280/X
+ sky130_fd_sc_hd__xor2_1_280/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__o21ai_1_68 vssd1 vccd1 sky130_fd_sc_hd__inv_2_56/Y sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_68/B1 sky130_fd_sc_hd__o21ai_1_68/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_291 sky130_fd_sc_hd__fa_2_198/A sky130_fd_sc_hd__and3_4_13/A
+ sky130_fd_sc_hd__xor2_1_291/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__o21ai_1_79 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_81/A2 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__o21ai_1_79/B1 sky130_fd_sc_hd__o21ai_1_79/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_300 vccd1 vssd1 sky130_fd_sc_hd__and3_4_11/X sky130_fd_sc_hd__and2_0_45/A
+ sky130_fd_sc_hd__and2_0_87/A sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__o21ai_1_512/B1 sky130_fd_sc_hd__and2b_4_8/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_240 vssd1 vccd1 sky130_fd_sc_hd__inv_2_176/A sky130_fd_sc_hd__buf_8_70/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_311 vccd1 vssd1 sky130_fd_sc_hd__and3_4_10/X sky130_fd_sc_hd__buf_2_19/X
+ sky130_fd_sc_hd__buf_6_5/X sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__o21ai_1_526/B1 sky130_fd_sc_hd__and2b_4_7/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_251 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1_962/A sky130_fd_sc_hd__buf_4_8/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_322 vccd1 vssd1 sky130_fd_sc_hd__and3_4_11/X sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__buf_6_1/X sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__and2_0_38/A
+ sky130_fd_sc_hd__o21ai_1_540/B1 sky130_fd_sc_hd__and2b_4_8/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_262 vssd1 vccd1 sky130_fd_sc_hd__buf_12_41/A sky130_fd_sc_hd__buf_8_108/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_333 vccd1 vssd1 sky130_fd_sc_hd__and3_4_17/X sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__buf_6_2/X sky130_fd_sc_hd__nor2_2_20/Y sky130_fd_sc_hd__buf_4_7/X
+ sky130_fd_sc_hd__o21ai_1_554/B1 sky130_fd_sc_hd__nor2b_2_4/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_273 vssd1 vccd1 sky130_fd_sc_hd__buf_8_148/A sky130_fd_sc_hd__clkbuf_1_273/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_344 vccd1 vssd1 sky130_fd_sc_hd__and3_4_11/X sky130_fd_sc_hd__buf_4_0/X
+ sky130_fd_sc_hd__buf_2_23/X sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__buf_2_31/X
+ sky130_fd_sc_hd__o21ai_1_571/B1 sky130_fd_sc_hd__and2b_4_8/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_284 vssd1 vccd1 sky130_fd_sc_hd__buf_6_26/A sky130_fd_sc_hd__clkbuf_1_284/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_355 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__buf_2_23/X
+ sky130_fd_sc_hd__buf_2_31/X sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__buf_2_19/X
+ sky130_fd_sc_hd__o21ai_1_587/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_295 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_296/A sky130_fd_sc_hd__buf_4_30/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_366 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__buf_2_23/X
+ sky130_fd_sc_hd__buf_2_31/X sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__buf_2_19/X
+ sky130_fd_sc_hd__o21ai_1_606/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_377 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__inv_6_0/Y sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__o21ai_1_624/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_388 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__or2_0_9/B
+ sky130_fd_sc_hd__or2_0_9/A sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__or2_0_4/B
+ sky130_fd_sc_hd__o21ai_1_649/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_399 vccd1 vssd1 sky130_fd_sc_hd__and3_4_25/X sky130_fd_sc_hd__buf_2_4/A
+ sky130_fd_sc_hd__buf_2_20/X sky130_fd_sc_hd__nor2_1_186/Y sky130_fd_sc_hd__buf_2_21/X
+ sky130_fd_sc_hd__o21ai_1_665/B1 sky130_fd_sc_hd__nor2b_1_17/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__buf_4_1 vccd1 vssd1 sky130_fd_sc_hd__buf_4_1/X sky130_fd_sc_hd__buf_4_7/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__and2_0_260 vccd1 vssd1 sky130_fd_sc_hd__and2_0_260/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__xor2_1_648/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_271 vccd1 vssd1 sky130_fd_sc_hd__and2_0_271/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__and2_0_271/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__a21oi_2_12 sky130_fd_sc_hd__a21oi_2_12/B1 sky130_fd_sc_hd__or2_0_37/X
+ sky130_fd_sc_hd__xnor2_1_98/B sky130_fd_sc_hd__xor2_1_346/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_2
Xsky130_fd_sc_hd__and2_0_282 vccd1 vssd1 sky130_fd_sc_hd__and2_0_282/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__fa_2_415/SUM vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_293 vccd1 vssd1 sky130_fd_sc_hd__and2_0_293/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_14/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_12_508 sky130_fd_sc_hd__buf_12_508/A sky130_fd_sc_hd__buf_12_619/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_519 sky130_fd_sc_hd__buf_12_519/A sky130_fd_sc_hd__buf_12_519/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__inv_4_1 sky130_fd_sc_hd__inv_4_1/Y sky130_fd_sc_hd__inv_4_1/A vccd1
+ vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__nand2_1_109 sky130_fd_sc_hd__o21ai_1_83/B1 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__xor2_1_330/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_708 sky130_fd_sc_hd__nand4_1_0/C sky130_fd_sc_hd__or4_1_1/C
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_719 sky130_fd_sc_hd__nor2b_1_98/A sky130_fd_sc_hd__xor2_1_678/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__or2_0_106 sky130_fd_sc_hd__or2_0_106/A sky130_fd_sc_hd__or2_0_106/X
+ sky130_fd_sc_hd__or2_0_106/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__o21ai_1_250 vssd1 vccd1 sky130_fd_sc_hd__inv_2_10/Y sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__o21ai_1_250/B1 sky130_fd_sc_hd__xor2_1_73/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_261 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_261/A2 sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__o21ai_1_261/B1 sky130_fd_sc_hd__xor2_1_85/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_272 vssd1 vccd1 sky130_fd_sc_hd__buf_2_5/X sky130_fd_sc_hd__nand2b_1_7/Y
+ sky130_fd_sc_hd__o21ai_1_272/B1 sky130_fd_sc_hd__xor2_1_93/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_283 vssd1 vccd1 sky130_fd_sc_hd__inv_2_26/Y sky130_fd_sc_hd__nand2b_1_5/Y
+ sky130_fd_sc_hd__nand2_1_155/Y sky130_fd_sc_hd__xor2_1_103/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_294 vssd1 vccd1 sky130_fd_sc_hd__inv_2_16/Y sky130_fd_sc_hd__nand2b_1_7/Y
+ sky130_fd_sc_hd__o21ai_1_294/B1 sky130_fd_sc_hd__xor2_1_115/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_704 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_715 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_726 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_610 sky130_fd_sc_hd__xnor2_1_170/A sky130_fd_sc_hd__nand2_1_611/Y
+ sky130_fd_sc_hd__nand2_1_610/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_737 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_621 sky130_fd_sc_hd__xnor2_1_175/A sky130_fd_sc_hd__nand2_1_622/Y
+ sky130_fd_sc_hd__nand2_1_621/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_748 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_632 sky130_fd_sc_hd__nand2_1_632/Y sky130_fd_sc_hd__nor2_1_211/A
+ sky130_fd_sc_hd__nor2_1_211/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_759 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_643 sky130_fd_sc_hd__nand2_1_643/Y sky130_fd_sc_hd__nand2_1_653/Y
+ sky130_fd_sc_hd__nand2_1_649/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_654 sky130_fd_sc_hd__xor2_1_632/A sky130_fd_sc_hd__nand2_1_655/Y
+ sky130_fd_sc_hd__nand2_1_654/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_665 sky130_fd_sc_hd__nand2_1_665/Y sky130_fd_sc_hd__mux2_2_15/X
+ sky130_fd_sc_hd__mux2_2_35/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_2_1 sky130_fd_sc_hd__nor2_2_7/A sky130_fd_sc_hd__and3_4_7/B
+ sky130_fd_sc_hd__nor2b_2_1/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_2
Xsky130_fd_sc_hd__nand2_1_676 sky130_fd_sc_hd__xor2_1_643/B sky130_fd_sc_hd__nand2_1_677/Y
+ sky130_fd_sc_hd__nand2_1_676/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_687 sky130_fd_sc_hd__nand2_1_687/Y sky130_fd_sc_hd__or2_0_78/A
+ sky130_fd_sc_hd__or2_0_78/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_698 sky130_fd_sc_hd__xnor2_1_197/A sky130_fd_sc_hd__nand2_1_699/Y
+ sky130_fd_sc_hd__or2_1_10/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_1703 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1714 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_13 sky130_fd_sc_hd__inv_2_13/A sky130_fd_sc_hd__inv_2_13/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1725 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_24 sky130_fd_sc_hd__inv_2_24/A sky130_fd_sc_hd__inv_2_24/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1736 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_35 sky130_fd_sc_hd__inv_2_35/A sky130_fd_sc_hd__inv_2_35/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1747 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_46 sky130_fd_sc_hd__inv_2_46/A sky130_fd_sc_hd__inv_2_46/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_450 sky130_fd_sc_hd__dfxtp_1_450/Q sky130_fd_sc_hd__dfxtp_1_451/CLK
+ sky130_fd_sc_hd__nor2b_1_97/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1758 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_57 sky130_fd_sc_hd__inv_2_57/A sky130_fd_sc_hd__inv_2_57/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_461 sky130_fd_sc_hd__mux2_8_0/S sky130_fd_sc_hd__edfxbp_1_0/CLK
+ la_data_out[47] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1769 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_68 sky130_fd_sc_hd__inv_2_68/A sky130_fd_sc_hd__inv_2_68/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_472 sky130_fd_sc_hd__dfxtp_1_472/Q sky130_fd_sc_hd__dfxtp_1_479/CLK
+ sky130_fd_sc_hd__and2_0_383/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_79 sky130_fd_sc_hd__inv_2_79/A sky130_fd_sc_hd__inv_2_79/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_483 la_data_out[50] sky130_fd_sc_hd__dfxtp_1_489/CLK sky130_fd_sc_hd__and2_0_375/X
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_2_3 sky130_fd_sc_hd__nand2_2_3/Y sky130_fd_sc_hd__nand2_2_3/A
+ sky130_fd_sc_hd__nand2_2_3/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__dfxtp_1_494 la_data_out[43] sky130_fd_sc_hd__dfxtp_1_498/CLK sky130_fd_sc_hd__and2_0_379/X
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2b_1_20 sky130_fd_sc_hd__nand2b_1_20/Y sky130_fd_sc_hd__and3_4_24/C
+ sky130_fd_sc_hd__and3_4_24/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__nand2b_1_31 sky130_fd_sc_hd__nand2b_1_31/Y sky130_fd_sc_hd__nand2_1_845/A
+ sky130_fd_sc_hd__nand2b_1_31/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a222oi_1_130 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__buf_4_5/X sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__o21ai_1_270/B1 sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_141 vccd1 vssd1 sky130_fd_sc_hd__and3_4_7/X sky130_fd_sc_hd__buf_4_6/X
+ sky130_fd_sc_hd__buf_4_1/X sky130_fd_sc_hd__nor2_2_7/Y sky130_fd_sc_hd__nor2_2_5/A
+ sky130_fd_sc_hd__o21ai_1_286/B1 sky130_fd_sc_hd__nor2b_2_1/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_152 vccd1 vssd1 sky130_fd_sc_hd__and3_4_2/X sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__nor2_1_87/A sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__o21ai_1_298/B1 sky130_fd_sc_hd__and2b_4_4/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_300 sky130_fd_sc_hd__nor2_2_22/B sky130_fd_sc_hd__or2_1_8/B
+ sky130_fd_sc_hd__fa_2_300/A sky130_fd_sc_hd__fa_2_300/B sky130_fd_sc_hd__fa_2_307/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_163 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__buf_6_4/X
+ sky130_fd_sc_hd__buf_6_0/X sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__o21ai_1_313/B1 sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_311 sky130_fd_sc_hd__fa_2_306/CIN sky130_fd_sc_hd__fa_2_316/A
+ sky130_fd_sc_hd__fa_2_311/A sky130_fd_sc_hd__fa_2_311/B sky130_fd_sc_hd__xor2_1_472/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_174 vccd1 vssd1 sky130_fd_sc_hd__and3_4_8/X sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__buf_2_32/X sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__o21ai_1_328/B1 sky130_fd_sc_hd__nor2b_2_2/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_322 sky130_fd_sc_hd__fa_2_315/A sky130_fd_sc_hd__fa_2_323/B
+ sky130_fd_sc_hd__fa_2_322/A sky130_fd_sc_hd__fa_2_322/B sky130_fd_sc_hd__fa_2_322/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_185 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__nor2_1_87/A sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__o21ai_1_343/B1 sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_333 sky130_fd_sc_hd__or2_1_7/A sky130_fd_sc_hd__nor2_2_24/B
+ sky130_fd_sc_hd__fa_2_333/A sky130_fd_sc_hd__fa_2_333/B sky130_fd_sc_hd__fa_2_333/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_196 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__buf_4_1/X
+ sky130_fd_sc_hd__nor2_2_5/A sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__nor2_2_5/B
+ sky130_fd_sc_hd__o21ai_1_361/B1 sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_344 sky130_fd_sc_hd__fa_2_337/A sky130_fd_sc_hd__fa_2_345/A
+ sky130_fd_sc_hd__fa_2_344/A sky130_fd_sc_hd__fa_2_344/B sky130_fd_sc_hd__xor2_1_510/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_355 sky130_fd_sc_hd__nor2_2_23/A sky130_fd_sc_hd__or2_1_5/B
+ sky130_fd_sc_hd__fa_2_355/A sky130_fd_sc_hd__fa_2_355/B sky130_fd_sc_hd__fa_2_355/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_366 sky130_fd_sc_hd__fa_2_362/B sky130_fd_sc_hd__fa_2_368/CIN
+ sky130_fd_sc_hd__fa_2_366/A sky130_fd_sc_hd__fa_2_366/B sky130_fd_sc_hd__fa_2_366/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_377 sky130_fd_sc_hd__fa_2_371/A sky130_fd_sc_hd__fa_2_378/B
+ sky130_fd_sc_hd__fa_2_377/A sky130_fd_sc_hd__fa_2_377/B sky130_fd_sc_hd__xor2_1_551/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_18 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_4_3/Y
+ sky130_fd_sc_hd__dfxtp_1_176/CLK sky130_fd_sc_hd__o21ai_2_1/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_388 sky130_fd_sc_hd__fa_2_385/CIN sky130_fd_sc_hd__fah_1_16/A
+ sky130_fd_sc_hd__fa_2_388/A sky130_fd_sc_hd__fa_2_388/B sky130_fd_sc_hd__xor2_1_577/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_29 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_8_5/Y
+ sky130_fd_sc_hd__dfxtp_1_266/CLK sky130_fd_sc_hd__o21ai_2_4/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_399 sky130_fd_sc_hd__fah_1_9/B sky130_fd_sc_hd__fah_1_8/CI
+ sky130_fd_sc_hd__fa_2_399/A sky130_fd_sc_hd__fa_2_399/B sky130_fd_sc_hd__xor2_1_591/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_8_60 sky130_fd_sc_hd__clkinv_8_61/A sky130_fd_sc_hd__clkinv_8_2/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_71 sky130_fd_sc_hd__clkinv_8_72/A sky130_fd_sc_hd__clkinv_8_71/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_82 sky130_fd_sc_hd__clkinv_8_83/A sky130_fd_sc_hd__clkinv_8_82/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_80 sky130_fd_sc_hd__buf_8_153/X sky130_fd_sc_hd__buf_12_80/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_91 sky130_fd_sc_hd__buf_8_132/X sky130_fd_sc_hd__buf_12_91/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__nor2_1_109 sky130_fd_sc_hd__xnor2_1_71/Y sky130_fd_sc_hd__nor2_1_109/Y
+ sky130_fd_sc_hd__xnor2_1_68/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_18 sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__dfxtp_1_282/Q sky130_fd_sc_hd__o211ai_1_6/Y sky130_fd_sc_hd__nand2_2_4/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_29 sky130_fd_sc_hd__nor2_4_0/Y sky130_fd_sc_hd__nor2_2_0/Y
+ sky130_fd_sc_hd__dfxtp_1_326/Q sky130_fd_sc_hd__or2_0_95/A sky130_fd_sc_hd__nand2_2_6/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_305 sky130_fd_sc_hd__buf_12_305/A sky130_fd_sc_hd__buf_12_491/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_316 sky130_fd_sc_hd__buf_12_43/X sky130_fd_sc_hd__buf_12_645/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_327 sky130_fd_sc_hd__buf_12_47/X sky130_fd_sc_hd__buf_12_659/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_338 sky130_fd_sc_hd__buf_12_338/A sky130_fd_sc_hd__buf_12_536/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_349 sky130_fd_sc_hd__buf_12_90/X sky130_fd_sc_hd__buf_12_596/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_208 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__and2b_4_7/X sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__a22oi_1_208/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_219 sky130_fd_sc_hd__or2_0_72/B sky130_fd_sc_hd__or2_0_72/A
+ sky130_fd_sc_hd__and2b_4_11/X sky130_fd_sc_hd__nor2_4_16/Y sky130_fd_sc_hd__a22oi_1_219/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor3_2_0 sky130_fd_sc_hd__or4_1_0/X sky130_fd_sc_hd__nor3_2_0/Y
+ sky130_fd_sc_hd__ha_2_6/A sky130_fd_sc_hd__ha_2_3/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor3_2
Xsky130_fd_sc_hd__clkinv_1_505 sky130_fd_sc_hd__nand2_1_481/A sky130_fd_sc_hd__nor2_1_161/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_516 sky130_fd_sc_hd__a21oi_2_19/B1 sky130_fd_sc_hd__nand2_1_587/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_527 sky130_fd_sc_hd__nor2_1_168/B sky130_fd_sc_hd__nand2_1_526/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_538 sky130_fd_sc_hd__a21oi_2_15/B1 sky130_fd_sc_hd__nand2_1_534/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_549 sky130_fd_sc_hd__clkinv_1_549/Y sky130_fd_sc_hd__o21a_1_4/A2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_30 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_30/Y
+ sky130_fd_sc_hd__nor2_1_30/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_41 sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__inv_2_5/A
+ sky130_fd_sc_hd__nor2_1_2/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_52 sky130_fd_sc_hd__nor2_1_52/B sky130_fd_sc_hd__nor2_1_52/Y
+ sky130_fd_sc_hd__nor2_1_52/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_63 sky130_fd_sc_hd__nor2_1_63/B sky130_fd_sc_hd__nor2_1_63/Y
+ sky130_fd_sc_hd__nor2_1_63/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_18 sky130_fd_sc_hd__buf_8_29/A sky130_fd_sc_hd__inv_2_132/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_74 sky130_fd_sc_hd__nor2_1_74/B sky130_fd_sc_hd__nor2_1_74/Y
+ sky130_fd_sc_hd__nor2_1_74/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_29 sky130_fd_sc_hd__nand2_1_10/Y sky130_fd_sc_hd__clkinv_4_29/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_85 sky130_fd_sc_hd__nor2_1_85/B sky130_fd_sc_hd__nor2_1_85/Y
+ sky130_fd_sc_hd__nor2_1_87/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_96 sky130_fd_sc_hd__nor2_2_4/Y sky130_fd_sc_hd__nor2_1_96/Y
+ sky130_fd_sc_hd__nor2_2_5/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_12_501 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_512 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_523 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_534 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_545 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_556 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_440 sky130_fd_sc_hd__nand2_1_440/Y sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__buf_6_1/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_567 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_451 sky130_fd_sc_hd__nand2_1_451/Y sky130_fd_sc_hd__nor2_1_152/A
+ sky130_fd_sc_hd__nor2_1_152/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_578 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_462 sky130_fd_sc_hd__xnor2_1_63/B sky130_fd_sc_hd__nand2_1_463/Y
+ sky130_fd_sc_hd__nand2_1_462/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_589 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_473 sky130_fd_sc_hd__xnor2_1_119/A sky130_fd_sc_hd__nand2_1_474/Y
+ sky130_fd_sc_hd__nand2_1_473/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_484 sky130_fd_sc_hd__xor2_1_419/A sky130_fd_sc_hd__nand2_1_485/Y
+ sky130_fd_sc_hd__nand2_1_484/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_495 sky130_fd_sc_hd__nand2_1_495/Y sky130_fd_sc_hd__nor2_1_183/Y
+ sky130_fd_sc_hd__or2_0_72/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_20 sky130_fd_sc_hd__or2_0_84/A sky130_fd_sc_hd__fa_2_440/A
+ sky130_fd_sc_hd__nor2b_1_20/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_31 sky130_fd_sc_hd__fa_2_417/A sky130_fd_sc_hd__nor2b_1_31/Y
+ sky130_fd_sc_hd__buf_2_214/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_42 sky130_fd_sc_hd__mux2_2_43/X sky130_fd_sc_hd__fa_2_472/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_53 sky130_fd_sc_hd__or2_1_11/B sky130_fd_sc_hd__nor2b_1_53/Y
+ sky130_fd_sc_hd__buf_2_214/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1020 sky130_fd_sc_hd__clkinv_1_1022/A sky130_fd_sc_hd__inv_12_1/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_64 sky130_fd_sc_hd__or2_0_79/A sky130_fd_sc_hd__fa_2_483/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1031 sky130_fd_sc_hd__clkbuf_1_273/A sky130_fd_sc_hd__clkinv_1_1031/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_75 la_data_out[72] sky130_fd_sc_hd__nor2b_1_75/Y sky130_fd_sc_hd__mux2_4_5/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1042 sky130_fd_sc_hd__inv_2_175/A sky130_fd_sc_hd__inv_2_121/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1500 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_86 sky130_fd_sc_hd__or2_0_83/A sky130_fd_sc_hd__nor2b_1_86/Y
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1053 sky130_fd_sc_hd__inv_2_186/A sky130_fd_sc_hd__clkbuf_1_275/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1511 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_97 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_97/Y
+ sky130_fd_sc_hd__nor2b_1_97/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1064 sky130_fd_sc_hd__clkinv_4_44/A sky130_fd_sc_hd__buf_8_121/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_5 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_8/A sky130_fd_sc_hd__xnor2_1_5/Y
+ sky130_fd_sc_hd__xnor2_1_5/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_1522 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1075 sky130_fd_sc_hd__a22o_1_80/B2 la_data_out[57] vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1533 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1086 sky130_fd_sc_hd__o21ai_1_919/A1 la_data_out[56] vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1544 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1097 sky130_fd_sc_hd__inv_4_11/A wbs_adr_i[2] vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1555 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1566 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1577 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_280 sky130_fd_sc_hd__dfxtp_1_280/Q sky130_fd_sc_hd__dfxtp_1_2/CLK
+ sky130_fd_sc_hd__and2_0_256/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1588 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_291 sky130_fd_sc_hd__a22oi_1_0/B2 sky130_fd_sc_hd__dfxtp_1_2/CLK
+ sky130_fd_sc_hd__and2_0_267/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1599 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__mux2_4_1 sky130_fd_sc_hd__or2_1_10/B sky130_fd_sc_hd__mux2_8_1/S
+ sky130_fd_sc_hd__buf_6_16/X sky130_fd_sc_hd__mux2_4_1/A1 vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__mux2_4
Xsky130_fd_sc_hd__o22ai_1_0 sky130_fd_sc_hd__o22ai_1_0/A2 sky130_fd_sc_hd__o22ai_1_0/B1
+ sky130_fd_sc_hd__o22ai_1_0/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__o22ai_1_9/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_130 sky130_fd_sc_hd__fa_2_127/CIN sky130_fd_sc_hd__fa_2_131/A
+ sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__fa_2_130/B sky130_fd_sc_hd__xor2_1_182/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_141 sky130_fd_sc_hd__fa_2_140/CIN sky130_fd_sc_hd__or2_0_21/A
+ sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__fa_2_141/B sky130_fd_sc_hd__xor2_1_205/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_152 sky130_fd_sc_hd__fa_2_143/B sky130_fd_sc_hd__fa_2_158/CIN
+ sky130_fd_sc_hd__fa_2_152/A sky130_fd_sc_hd__fa_2_152/B sky130_fd_sc_hd__fa_2_152/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_163 sky130_fd_sc_hd__fa_2_158/A sky130_fd_sc_hd__fa_2_168/A
+ sky130_fd_sc_hd__fa_2_163/A sky130_fd_sc_hd__fa_2_163/B sky130_fd_sc_hd__xor2_1_248/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and3_4_2 sky130_fd_sc_hd__nor2_4_9/B sky130_fd_sc_hd__nor2_4_9/A
+ sky130_fd_sc_hd__and3_4_2/C sky130_fd_sc_hd__and3_4_2/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__fa_2_174 sky130_fd_sc_hd__fa_2_167/A sky130_fd_sc_hd__fa_2_175/B
+ sky130_fd_sc_hd__fa_2_174/A sky130_fd_sc_hd__fa_2_174/B sky130_fd_sc_hd__fa_2_174/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_185 sky130_fd_sc_hd__nor2_2_11/A sky130_fd_sc_hd__or2_0_29/B
+ sky130_fd_sc_hd__fa_2_185/A sky130_fd_sc_hd__fa_2_185/B sky130_fd_sc_hd__fa_2_185/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_196 sky130_fd_sc_hd__fa_2_189/A sky130_fd_sc_hd__fa_2_197/B
+ sky130_fd_sc_hd__fa_2_196/A sky130_fd_sc_hd__fa_2_196/B sky130_fd_sc_hd__fa_2_196/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o22ai_1_40 sky130_fd_sc_hd__nor2_1_27/A sky130_fd_sc_hd__o22ai_1_40/B1
+ sky130_fd_sc_hd__o22ai_1_40/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_51 sky130_fd_sc_hd__nor2_1_16/A sky130_fd_sc_hd__o22ai_1_51/B1
+ sky130_fd_sc_hd__o22ai_1_51/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_62 sky130_fd_sc_hd__nor2_1_5/A sky130_fd_sc_hd__o22ai_1_1/A2
+ sky130_fd_sc_hd__o22ai_1_62/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_180 vccd1 vssd1 sky130_fd_sc_hd__buf_2_180/X sky130_fd_sc_hd__inv_2_195/Y
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_73 sky130_fd_sc_hd__xnor2_1_253/Y sky130_fd_sc_hd__xnor2_1_224/Y
+ sky130_fd_sc_hd__fa_2_432/B sky130_fd_sc_hd__inv_2_65/Y sky130_fd_sc_hd__o22ai_1_99/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_191 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_3/D sky130_fd_sc_hd__dfxtp_1_4/Q
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_84 sky130_fd_sc_hd__xnor2_1_238/Y sky130_fd_sc_hd__xnor2_1_236/Y
+ sky130_fd_sc_hd__ha_2_14/B sky130_fd_sc_hd__inv_2_65/Y sky130_fd_sc_hd__o22ai_1_99/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_95 sky130_fd_sc_hd__xnor2_2_5/Y sky130_fd_sc_hd__xnor2_1_242/Y
+ sky130_fd_sc_hd__ha_2_13/A sky130_fd_sc_hd__xnor2_1_243/Y sky130_fd_sc_hd__o22ai_1_95/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_4_20 vccd1 vssd1 sky130_fd_sc_hd__buf_4_20/X sky130_fd_sc_hd__buf_4_20/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_31 vccd1 vssd1 sky130_fd_sc_hd__buf_4_31/X sky130_fd_sc_hd__buf_8_63/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_42 vccd1 vssd1 sky130_fd_sc_hd__buf_4_42/X sky130_fd_sc_hd__buf_4_42/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_12_102 sky130_fd_sc_hd__buf_4_34/X sky130_fd_sc_hd__buf_12_376/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_113 sky130_fd_sc_hd__buf_8_135/X sky130_fd_sc_hd__buf_12_425/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_124 sky130_fd_sc_hd__buf_8_133/X sky130_fd_sc_hd__buf_12_124/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_135 sky130_fd_sc_hd__buf_8_39/X sky130_fd_sc_hd__buf_12_384/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_146 sky130_fd_sc_hd__buf_12_26/X sky130_fd_sc_hd__buf_12_375/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_157 sky130_fd_sc_hd__buf_12_53/X sky130_fd_sc_hd__buf_12_303/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_80 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_8/A1 sky130_fd_sc_hd__clkbuf_1_80/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_168 sky130_fd_sc_hd__buf_12_42/X sky130_fd_sc_hd__buf_12_329/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_91 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_23/A1 sky130_fd_sc_hd__clkbuf_1_91/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_4_5 sky130_fd_sc_hd__nor2_2_5/B sky130_fd_sc_hd__buf_2_27/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_12_179 sky130_fd_sc_hd__buf_8_107/X sky130_fd_sc_hd__buf_12_179/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_302 sky130_fd_sc_hd__and2_0_246/A sky130_fd_sc_hd__a222oi_1_46/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_313 sky130_fd_sc_hd__o21ai_1_177/A2 sky130_fd_sc_hd__xnor2_1_6/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_324 sky130_fd_sc_hd__o21ai_1_207/A2 sky130_fd_sc_hd__xnor2_1_11/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_335 sky130_fd_sc_hd__o21ai_1_241/A2 sky130_fd_sc_hd__xnor2_1_17/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_346 sky130_fd_sc_hd__o21ai_1_261/A2 sky130_fd_sc_hd__xnor2_1_22/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_357 sky130_fd_sc_hd__nand2_1_227/A sky130_fd_sc_hd__nor2_1_69/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_368 sky130_fd_sc_hd__nand2_1_254/A sky130_fd_sc_hd__nor2_1_80/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_379 sky130_fd_sc_hd__nand2_1_268/A sky130_fd_sc_hd__nor2_1_87/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_2_9 sky130_fd_sc_hd__a21oi_2_9/B1 sky130_fd_sc_hd__or2_0_30/X
+ sky130_fd_sc_hd__xnor2_1_82/B sky130_fd_sc_hd__a21oi_2_9/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_2
Xsky130_fd_sc_hd__or2_0_60 sky130_fd_sc_hd__or2_0_60/A sky130_fd_sc_hd__or2_0_60/X
+ sky130_fd_sc_hd__or2_0_60/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__a31o_1_0 sky130_fd_sc_hd__nand3_1_5/B sky130_fd_sc_hd__nor2_2_1/B
+ sky130_fd_sc_hd__nand3_1_5/C sky130_fd_sc_hd__a31o_1_0/A3 sky130_fd_sc_hd__a31o_1_0/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__a31o_1
Xsky130_fd_sc_hd__or2_0_71 sky130_fd_sc_hd__or2_0_72/A sky130_fd_sc_hd__or2_0_71/X
+ sky130_fd_sc_hd__or2_0_71/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__clkinv_4_5 sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__clkinv_8_5/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__or2_0_82 sky130_fd_sc_hd__or2_0_82/A sky130_fd_sc_hd__or2_0_82/X
+ sky130_fd_sc_hd__or2_0_82/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_93 sky130_fd_sc_hd__or2_0_93/A sky130_fd_sc_hd__or2_0_93/X
+ sky130_fd_sc_hd__or2_0_93/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__buf_12_680 sky130_fd_sc_hd__mux2_2_34/X la_data_out[68] vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_320 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_331 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_342 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_353 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_364 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_375 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_386 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_270 sky130_fd_sc_hd__xor2_1_171/B sky130_fd_sc_hd__nand2_1_271/Y
+ sky130_fd_sc_hd__nand2_1_270/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_397 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_281 sky130_fd_sc_hd__xor2_1_186/B sky130_fd_sc_hd__nand2_1_282/Y
+ sky130_fd_sc_hd__nand2_1_281/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_880 sky130_fd_sc_hd__clkinv_1_880/Y sky130_fd_sc_hd__inv_4_16/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xor2_1_109 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__fa_2_74/A
+ sky130_fd_sc_hd__xor2_1_109/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_292 sky130_fd_sc_hd__nand2_1_292/Y sky130_fd_sc_hd__nor2_2_5/A
+ sky130_fd_sc_hd__nor2_2_5/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_891 sky130_fd_sc_hd__clkinv_1_891/Y sky130_fd_sc_hd__clkinv_4_88/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1330 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1341 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_80 sky130_fd_sc_hd__conb_1_80/LO sky130_fd_sc_hd__conb_1_80/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1352 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_91 sky130_fd_sc_hd__conb_1_91/LO sky130_fd_sc_hd__conb_1_91/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1363 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1374 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_805 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_9/X sky130_fd_sc_hd__nand2b_2_6/Y
+ sky130_fd_sc_hd__o21ai_1_805/B1 sky130_fd_sc_hd__xor2_1_578/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1385 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_816 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_597/A sky130_fd_sc_hd__nor2_1_200/Y
+ sky130_fd_sc_hd__nand2_1_613/Y sky130_fd_sc_hd__xnor2_1_169/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1396 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_827 vssd1 vccd1 sky130_fd_sc_hd__inv_2_49/Y sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_827/B1 sky130_fd_sc_hd__xor2_1_601/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_838 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_3/Y sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_838/B1 sky130_fd_sc_hd__xor2_1_611/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_849 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_9/X sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_849/B1 sky130_fd_sc_hd__xor2_1_623/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nand2b_2_6 sky130_fd_sc_hd__nor2_4_16/B sky130_fd_sc_hd__nand2b_2_6/Y
+ sky130_fd_sc_hd__nor2_4_16/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_2
Xsky130_fd_sc_hd__xor2_1_610 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__fa_2_405/B
+ sky130_fd_sc_hd__xor2_1_610/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_621 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__xor2_1_621/X
+ sky130_fd_sc_hd__xor2_1_621/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_632 sky130_fd_sc_hd__o21a_1_5/X sky130_fd_sc_hd__xor2_1_632/X
+ sky130_fd_sc_hd__xor2_1_632/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_643 sky130_fd_sc_hd__xor2_1_643/B sky130_fd_sc_hd__xor2_1_643/X
+ sky130_fd_sc_hd__xor2_1_643/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_654 sky130_fd_sc_hd__xor2_1_654/B sky130_fd_sc_hd__xor2_1_654/X
+ sky130_fd_sc_hd__xor2_1_654/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_665 sky130_fd_sc_hd__xor2_1_665/B sky130_fd_sc_hd__or2_0_91/B
+ sky130_fd_sc_hd__xor2_1_665/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_676 sky130_fd_sc_hd__xor2_1_676/B sky130_fd_sc_hd__xor2_1_676/X
+ sky130_fd_sc_hd__xor2_1_676/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_687 sky130_fd_sc_hd__xor2_1_687/B sky130_fd_sc_hd__xor2_1_687/X
+ sky130_fd_sc_hd__xor2_1_687/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkinv_1_19 la_data_out[108] sky130_fd_sc_hd__conb_1_123/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__fa_2_6 sky130_fd_sc_hd__xor3_1_8/A sky130_fd_sc_hd__fa_2_3/B sky130_fd_sc_hd__fa_2_6/A
+ sky130_fd_sc_hd__fa_2_6/B sky130_fd_sc_hd__fa_2_6/CIN vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a211o_1_12 vssd1 vccd1 sky130_fd_sc_hd__fa_2_262/B sky130_fd_sc_hd__dfxtp_1_75/Q
+ sky130_fd_sc_hd__nor2_1_16/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_12/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__a211o_1_23 vssd1 vccd1 sky130_fd_sc_hd__fa_2_206/A sky130_fd_sc_hd__dfxtp_1_86/Q
+ sky130_fd_sc_hd__nor2_1_27/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_23/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__clkinv_1_110 io_oeb[29] sky130_fd_sc_hd__conb_1_32/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_121 io_oeb[18] sky130_fd_sc_hd__conb_1_21/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_132 io_oeb[7] sky130_fd_sc_hd__conb_1_10/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_143 sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__nor2_2_1/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_154 sky130_fd_sc_hd__o22ai_1_33/B1 sky130_fd_sc_hd__dfxtp_1_187/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_165 sky130_fd_sc_hd__o21ai_1_6/A2 sky130_fd_sc_hd__dfxtp_1_121/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_176 sky130_fd_sc_hd__nor2_1_27/A sky130_fd_sc_hd__dfxtp_1_150/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_8 sky130_fd_sc_hd__buf_8_8/A sky130_fd_sc_hd__buf_8_8/X vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__clkinv_1_187 sky130_fd_sc_hd__o22ai_1_44/B1 sky130_fd_sc_hd__dfxtp_1_178/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_12 sky130_fd_sc_hd__inv_2_66/Y sky130_fd_sc_hd__xor2_1_664/X
+ sky130_fd_sc_hd__a22o_1_12/X sky130_fd_sc_hd__a22o_1_9/B2 sky130_fd_sc_hd__xor2_1_656/X
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_198 sky130_fd_sc_hd__o22ai_1_16/B1 sky130_fd_sc_hd__dfxtp_1_111/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_23 sky130_fd_sc_hd__buf_2_63/A sky130_fd_sc_hd__buf_2_98/X
+ sky130_fd_sc_hd__a22o_1_23/X sky130_fd_sc_hd__a22o_1_23/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_34 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__buf_2_109/X
+ sky130_fd_sc_hd__a22o_1_34/X sky130_fd_sc_hd__a22o_1_34/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_45 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__buf_2_120/X
+ sky130_fd_sc_hd__a22o_1_45/X sky130_fd_sc_hd__a22o_1_45/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_56 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__buf_2_47/A
+ sky130_fd_sc_hd__a22o_1_56/X sky130_fd_sc_hd__ha_2_27/SUM sky130_fd_sc_hd__a22o_1_71/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_67 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__a22o_1_67/A2
+ sky130_fd_sc_hd__a22o_1_67/X sky130_fd_sc_hd__ha_2_36/SUM sky130_fd_sc_hd__a22o_1_71/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_78 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__a22o_1_78/A2
+ sky130_fd_sc_hd__a22o_1_78/X sky130_fd_sc_hd__ha_2_24/SUM sky130_fd_sc_hd__nor2_1_269/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_2_2 sky130_fd_sc_hd__clkinv_2_2/Y sky130_fd_sc_hd__clkinv_2_2/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__nor2_1_270 sky130_fd_sc_hd__nor2_4_0/B sky130_fd_sc_hd__o31ai_1_1/A1
+ sky130_fd_sc_hd__nor2_4_0/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_281 wbs_adr_i[2] sky130_fd_sc_hd__a21o_2_1/B1 wbs_adr_i[3]
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_12_150 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_161 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_172 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_183 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_13 sky130_fd_sc_hd__nand2_1_13/Y sky130_fd_sc_hd__nand2_1_13/B
+ sky130_fd_sc_hd__nand2_1_13/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_194 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_24 sky130_fd_sc_hd__nand2_8_3/B sky130_fd_sc_hd__nand2_1_8/B
+ sky130_fd_sc_hd__mux2_2_38/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_35 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__nand2_1_8/B
+ sky130_fd_sc_hd__mux2_2_49/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_240 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_4/B sky130_fd_sc_hd__xnor2_1_240/Y
+ la_data_out[71] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_46 sky130_fd_sc_hd__nand2_1_46/Y sky130_fd_sc_hd__nand2_1_7/B
+ la_data_out[68] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_251 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_5/B sky130_fd_sc_hd__xnor2_1_251/Y
+ sky130_fd_sc_hd__or2_0_84/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_57 sky130_fd_sc_hd__nand2_1_57/Y sky130_fd_sc_hd__nand2_1_57/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_262 vssd1 vccd1 la_data_out[81] sky130_fd_sc_hd__xnor2_1_262/Y
+ sky130_fd_sc_hd__or2_0_80/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_68 sky130_fd_sc_hd__nand2_1_68/Y sky130_fd_sc_hd__nand2_1_68/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_273 vssd1 vccd1 sky130_fd_sc_hd__or2_0_82/B sky130_fd_sc_hd__xnor2_1_273/Y
+ sky130_fd_sc_hd__or2_0_79/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_79 sky130_fd_sc_hd__nand2_1_79/Y sky130_fd_sc_hd__nand2_1_79/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_284 vssd1 vccd1 la_data_out[81] sky130_fd_sc_hd__xnor2_1_284/Y
+ sky130_fd_sc_hd__or2_0_79/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_295 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_295/B sky130_fd_sc_hd__xnor2_1_295/Y
+ sky130_fd_sc_hd__xnor2_1_295/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_1160 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1171 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_602 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_399/B sky130_fd_sc_hd__nor2_1_154/Y
+ sky130_fd_sc_hd__nand2_1_457/Y sky130_fd_sc_hd__xnor2_1_113/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1182 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_613 vssd1 vccd1 sky130_fd_sc_hd__inv_2_28/Y sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_613/B1 sky130_fd_sc_hd__xor2_1_405/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1193 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_624 vssd1 vccd1 sky130_fd_sc_hd__buf_2_10/X sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_624/B1 sky130_fd_sc_hd__xor2_1_416/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_635 vssd1 vccd1 sky130_fd_sc_hd__inv_2_47/Y sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_635/B1 sky130_fd_sc_hd__xor2_1_587/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_646 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_679/A2 sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_646/B1 sky130_fd_sc_hd__xor2_1_433/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_657 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_780/A2 sky130_fd_sc_hd__nand2b_1_16/Y
+ sky130_fd_sc_hd__o21ai_1_657/B1 sky130_fd_sc_hd__xor2_1_442/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_668 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_733/A2 sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__o21ai_1_668/B1 sky130_fd_sc_hd__xor2_1_451/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_679 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_679/A2 sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_679/B1 sky130_fd_sc_hd__xor2_1_460/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fah_1_0 sky130_fd_sc_hd__or2_0_11/A sky130_fd_sc_hd__fah_1_0/B sky130_fd_sc_hd__fah_1_0/A
+ sky130_fd_sc_hd__nor2_1_43/B sky130_fd_sc_hd__fah_1_0/CI vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__fah_1
Xsky130_fd_sc_hd__xor2_1_440 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__fa_2_290/A
+ sky130_fd_sc_hd__xor2_1_440/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_451 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__fa_2_292/B
+ sky130_fd_sc_hd__xor2_1_451/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_462 sky130_fd_sc_hd__fa_2_357/A sky130_fd_sc_hd__xor2_1_462/X
+ sky130_fd_sc_hd__xor2_1_462/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_473 sky130_fd_sc_hd__fa_2_338/A sky130_fd_sc_hd__fa_2_312/B
+ sky130_fd_sc_hd__xor2_1_473/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_484 sky130_fd_sc_hd__fa_2_338/A sky130_fd_sc_hd__xor2_1_484/X
+ sky130_fd_sc_hd__xor2_1_484/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_495 sky130_fd_sc_hd__fa_2_338/A sky130_fd_sc_hd__fa_2_327/B
+ sky130_fd_sc_hd__xor2_1_495/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a222oi_1_504 vccd1 vssd1 sky130_fd_sc_hd__and3_4_18/X sky130_fd_sc_hd__or2_0_72/A
+ sky130_fd_sc_hd__or2_0_71/B sky130_fd_sc_hd__nor2_2_32/Y sky130_fd_sc_hd__buf_2_29/X
+ sky130_fd_sc_hd__o21ai_1_800/B1 sky130_fd_sc_hd__nor2b_2_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_515 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__buf_2_21/X
+ sky130_fd_sc_hd__nor2_1_87/A sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__o21ai_1_635/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__dfxtp_4_2 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_4_2/D sky130_fd_sc_hd__clkinv_4_4/Y
+ sky130_fd_sc_hd__or2_0_51/A vssd1 vccd1 sky130_fd_sc_hd__dfxtp_4
Xsky130_fd_sc_hd__a222oi_1_526 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__buf_4_7/A
+ sky130_fd_sc_hd__buf_4_0/A sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__buf_2_27/X
+ sky130_fd_sc_hd__o21ai_1_829/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_537 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__buf_2_25/A
+ sky130_fd_sc_hd__inv_6_0/Y sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__buf_8_0/A
+ sky130_fd_sc_hd__o21ai_1_847/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_548 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_422/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_454/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_745/A sky130_fd_sc_hd__dfxtp_1_390/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_559 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_411/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_443/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_756/A sky130_fd_sc_hd__dfxtp_1_379/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nor2b_1_104 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_104/Y
+ sky130_fd_sc_hd__nor2b_1_104/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_115 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_115/Y
+ sky130_fd_sc_hd__nor2b_1_115/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_126 sky130_fd_sc_hd__clkinv_4_45/Y sky130_fd_sc_hd__nor2b_1_126/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_137 sky130_fd_sc_hd__clkinv_4_56/Y sky130_fd_sc_hd__nor2b_1_137/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_148 sky130_fd_sc_hd__clkinv_4_67/Y sky130_fd_sc_hd__nor2b_1_148/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__fah_1_17 sky130_fd_sc_hd__nor2_1_253/A sky130_fd_sc_hd__fah_1_17/B
+ sky130_fd_sc_hd__fah_1_17/A sky130_fd_sc_hd__or2_1_12/B sky130_fd_sc_hd__fah_1_17/CI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__fah_1
Xsky130_fd_sc_hd__buf_6_5 vccd1 vssd1 sky130_fd_sc_hd__buf_6_5/X sky130_fd_sc_hd__buf_6_5/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__clkinv_2_40 sky130_fd_sc_hd__inv_2_166/A sky130_fd_sc_hd__clkinv_2_40/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_51 sky130_fd_sc_hd__buf_2_46/A sky130_fd_sc_hd__inv_2_199/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__or2_1_0 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__or2_1_0/X sky130_fd_sc_hd__or2_1_0/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_1
Xsky130_fd_sc_hd__sdlclkp_4_3 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_8_1/Y
+ sky130_fd_sc_hd__dfxtp_1_45/CLK sky130_fd_sc_hd__o21ai_1_0/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_6 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_6/Y
+ sky130_fd_sc_hd__nor2_1_6/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__dfxtp_1_109 sky130_fd_sc_hd__dfxtp_1_109/Q sky130_fd_sc_hd__dfxtp_1_99/CLK
+ sky130_fd_sc_hd__and2_0_176/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_410 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_476/A2 sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_410/B1 sky130_fd_sc_hd__xor2_1_221/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_421 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_421/A2 sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_421/B1 sky130_fd_sc_hd__xor2_1_230/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_432 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_472/A2 sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_432/B1 sky130_fd_sc_hd__xor2_1_239/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_443 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_7/X sky130_fd_sc_hd__nand2_1_352/Y
+ sky130_fd_sc_hd__a21oi_1_76/Y sky130_fd_sc_hd__xnor2_1_74/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_454 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_454/A2 sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_454/B1 sky130_fd_sc_hd__xor2_1_258/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_465 vssd1 vccd1 sky130_fd_sc_hd__inv_2_34/Y sky130_fd_sc_hd__nand2b_1_14/Y
+ sky130_fd_sc_hd__o21ai_1_465/B1 sky130_fd_sc_hd__xor2_1_268/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_476 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_476/A2 sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_476/B1 sky130_fd_sc_hd__xor2_1_278/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_3_3 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__o21ai_1_487 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_7/X sky130_fd_sc_hd__nand2_1_374/Y
+ sky130_fd_sc_hd__a21oi_1_80/Y sky130_fd_sc_hd__xnor2_1_83/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_498 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_125/Y sky130_fd_sc_hd__nor2_1_123/A
+ sky130_fd_sc_hd__nor2_1_122/Y sky130_fd_sc_hd__o21ai_1_498/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_908 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_919 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_803 sky130_fd_sc_hd__nand2_1_803/Y sky130_fd_sc_hd__or2_0_102/A
+ sky130_fd_sc_hd__or2_0_102/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_814 sky130_fd_sc_hd__xnor2_1_296/A sky130_fd_sc_hd__nand2_1_815/Y
+ sky130_fd_sc_hd__or2_0_105/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_825 sky130_fd_sc_hd__nand2_1_825/Y sky130_fd_sc_hd__nor2_1_262/A
+ sky130_fd_sc_hd__nor2_1_262/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_836 sky130_fd_sc_hd__xor2_1_687/B sky130_fd_sc_hd__nand2_1_837/Y
+ sky130_fd_sc_hd__nand2_1_836/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_847 sky130_fd_sc_hd__inv_2_151/A la_data_out[36] la_data_out[47]
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_858 sky130_fd_sc_hd__a21o_2_0/B1 sky130_fd_sc_hd__o21ai_1_915/Y
+ sky130_fd_sc_hd__nand2_1_858/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o21ai_1_14 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_19/B1 sky130_fd_sc_hd__inv_2_53/A
+ sky130_fd_sc_hd__o21ai_1_14/B1 sky130_fd_sc_hd__fa_2_90/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_25 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_8/B1 sky130_fd_sc_hd__nor2_4_4/B
+ sky130_fd_sc_hd__o21ai_1_25/B1 sky130_fd_sc_hd__fa_2_133/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_36 vssd1 vccd1 sky130_fd_sc_hd__inv_2_62/Y sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__o21ai_1_36/B1 sky130_fd_sc_hd__and2_0_4/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_47 vssd1 vccd1 sky130_fd_sc_hd__inv_2_63/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_91/Y sky130_fd_sc_hd__o21ai_1_47/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_270 sky130_fd_sc_hd__xor2_1_362/B sky130_fd_sc_hd__xor2_1_270/X
+ sky130_fd_sc_hd__xor2_1_270/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__o21ai_1_58 vssd1 vccd1 sky130_fd_sc_hd__inv_2_60/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_96/Y sky130_fd_sc_hd__o21ai_1_58/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_281 sky130_fd_sc_hd__fa_2_217/A sky130_fd_sc_hd__fa_2_191/B
+ sky130_fd_sc_hd__xor2_1_281/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__o21ai_1_69 vssd1 vccd1 sky130_fd_sc_hd__inv_2_56/Y sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__o21ai_1_69/B1 sky130_fd_sc_hd__o21ai_1_69/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_292 sky130_fd_sc_hd__xor2_1_383/B sky130_fd_sc_hd__fa_2_199/A
+ sky130_fd_sc_hd__xor2_1_292/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_230 vssd1 vccd1 sky130_fd_sc_hd__buf_8_124/A sky130_fd_sc_hd__buf_8_40/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_301 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__buf_4_3/X sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__o21ai_1_513/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_241 vssd1 vccd1 sky130_fd_sc_hd__buf_8_114/A sky130_fd_sc_hd__buf_8_69/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_312 vccd1 vssd1 sky130_fd_sc_hd__and3_4_11/X sky130_fd_sc_hd__and2_0_38/A
+ sky130_fd_sc_hd__and2_0_49/A sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__and2_0_45/A
+ sky130_fd_sc_hd__o21ai_1_527/B1 sky130_fd_sc_hd__and2b_4_8/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_252 vssd1 vccd1 sky130_fd_sc_hd__buf_8_146/A sky130_fd_sc_hd__clkbuf_1_51/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_323 vccd1 vssd1 sky130_fd_sc_hd__and3_4_17/X sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__buf_4_7/X sky130_fd_sc_hd__nor2_2_20/Y sky130_fd_sc_hd__buf_4_0/X
+ sky130_fd_sc_hd__o21ai_1_541/B1 sky130_fd_sc_hd__nor2b_2_4/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_263 vssd1 vccd1 sky130_fd_sc_hd__buf_12_42/A sky130_fd_sc_hd__buf_2_53/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_334 vccd1 vssd1 sky130_fd_sc_hd__and3_4_10/X sky130_fd_sc_hd__buf_4_7/X
+ sky130_fd_sc_hd__buf_4_0/X sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__buf_2_23/X
+ sky130_fd_sc_hd__o21ai_1_555/B1 sky130_fd_sc_hd__and2b_4_7/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_274 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_15/A1 sky130_fd_sc_hd__clkbuf_1_274/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_345 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__buf_2_19/X
+ sky130_fd_sc_hd__buf_6_5/X sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__o21ai_1_572/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_285 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_286/A sky130_fd_sc_hd__buf_8_100/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_356 vccd1 vssd1 sky130_fd_sc_hd__and3_4_10/X sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__inv_6_0/Y sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__o21ai_1_588/B1 sky130_fd_sc_hd__and2b_4_7/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_296 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_296/X sky130_fd_sc_hd__clkbuf_1_296/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_367 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__buf_4_0/X
+ sky130_fd_sc_hd__buf_2_23/X sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__buf_2_31/X
+ sky130_fd_sc_hd__o21ai_1_608/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_378 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__or2_0_52/B
+ sky130_fd_sc_hd__or2_0_53/A sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__o21ai_1_627/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_389 vccd1 vssd1 sky130_fd_sc_hd__and3_4_26/X sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__nor2_2_10/B sky130_fd_sc_hd__nor2_2_31/Y sky130_fd_sc_hd__buf_6_4/X
+ sky130_fd_sc_hd__o21ai_1_652/B1 sky130_fd_sc_hd__nor2b_1_12/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__buf_4_2 vccd1 vssd1 sky130_fd_sc_hd__buf_4_2/X sky130_fd_sc_hd__buf_4_2/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__and2_0_250 vccd1 vssd1 sky130_fd_sc_hd__and2_0_250/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__o21ai_1_37/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_261 vccd1 vssd1 sky130_fd_sc_hd__and2_0_261/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__and2_0_261/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_272 vccd1 vssd1 sky130_fd_sc_hd__and2_0_272/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__xor2_1_642/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__a21oi_2_13 sky130_fd_sc_hd__a21oi_2_13/B1 sky130_fd_sc_hd__or2_1_5/X
+ sky130_fd_sc_hd__xnor2_1_149/B sky130_fd_sc_hd__xor2_1_509/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_2
Xsky130_fd_sc_hd__and2_0_283 vccd1 vssd1 sky130_fd_sc_hd__and2_0_283/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__xor2_1_638/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_294 vccd1 vssd1 sky130_fd_sc_hd__and2_0_294/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_15/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_12_509 sky130_fd_sc_hd__buf_12_509/A sky130_fd_sc_hd__buf_12_509/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__sdlclkp_2_0 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_8_3/Y
+ sky130_fd_sc_hd__dfxtp_1_89/CLK sky130_fd_sc_hd__o21ai_2_0/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__inv_4_2 sky130_fd_sc_hd__inv_4_2/Y sky130_fd_sc_hd__inv_4_2/A vccd1
+ vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__clkinv_1_709 sky130_fd_sc_hd__nor2b_1_88/A sky130_fd_sc_hd__fa_2_460/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__or2_0_107 sky130_fd_sc_hd__or2_0_107/A sky130_fd_sc_hd__or2_0_107/X
+ sky130_fd_sc_hd__or2_0_107/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__o21ai_1_240 vssd1 vccd1 sky130_fd_sc_hd__inv_2_14/Y sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__o21ai_1_240/B1 sky130_fd_sc_hd__xor2_1_64/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_251 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_251/A2 sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__o21ai_1_251/B1 sky130_fd_sc_hd__xor2_1_74/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_262 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_2/X sky130_fd_sc_hd__or2_0_5/B
+ sky130_fd_sc_hd__o21a_1_0/A2 sky130_fd_sc_hd__xnor2_1_22/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_273 vssd1 vccd1 sky130_fd_sc_hd__inv_2_15/Y sky130_fd_sc_hd__nand2b_1_6/Y
+ sky130_fd_sc_hd__o21ai_1_273/B1 sky130_fd_sc_hd__xor2_1_94/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_284 vssd1 vccd1 sky130_fd_sc_hd__inv_2_20/Y sky130_fd_sc_hd__nand2b_2_0/Y
+ sky130_fd_sc_hd__o21ai_1_284/B1 sky130_fd_sc_hd__xor2_1_105/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_295 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_295/A2 sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__o21ai_1_295/B1 sky130_fd_sc_hd__xor2_1_116/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_705 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_716 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_600 sky130_fd_sc_hd__xor2_2_2/A sky130_fd_sc_hd__nand2_1_601/Y
+ sky130_fd_sc_hd__nand2_1_600/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_727 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_611 sky130_fd_sc_hd__nand2_1_611/Y sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__buf_2_21/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_738 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_622 sky130_fd_sc_hd__nand2_1_622/Y sky130_fd_sc_hd__nor2_1_206/A
+ sky130_fd_sc_hd__nor2_1_206/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_749 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_633 sky130_fd_sc_hd__xnor2_1_127/B sky130_fd_sc_hd__nand2_1_634/Y
+ sky130_fd_sc_hd__nand2_1_633/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_644 sky130_fd_sc_hd__xnor2_1_181/A sky130_fd_sc_hd__nand2_1_645/Y
+ sky130_fd_sc_hd__nand2_1_644/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_655 sky130_fd_sc_hd__nand2_1_655/Y sky130_fd_sc_hd__nor2_1_219/A
+ sky130_fd_sc_hd__xor2_1_633/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_666 sky130_fd_sc_hd__xnor2_1_189/A sky130_fd_sc_hd__nand2_1_667/Y
+ sky130_fd_sc_hd__or2_0_74/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_2_2 sky130_fd_sc_hd__nor2_2_8/A sky130_fd_sc_hd__and3_4_8/B
+ sky130_fd_sc_hd__nor2b_2_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_2
Xsky130_fd_sc_hd__nand2_1_677 sky130_fd_sc_hd__nand2_1_677/Y sky130_fd_sc_hd__mux2_2_8/X
+ sky130_fd_sc_hd__mux2_2_39/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_688 sky130_fd_sc_hd__xor2_1_646/B sky130_fd_sc_hd__nand2_1_689/Y
+ sky130_fd_sc_hd__nand2_1_688/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_699 sky130_fd_sc_hd__nand2_1_699/Y sky130_fd_sc_hd__or2_1_10/A
+ sky130_fd_sc_hd__or2_1_10/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_1704 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1715 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_14 sky130_fd_sc_hd__inv_2_14/A sky130_fd_sc_hd__inv_2_14/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1726 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_25 sky130_fd_sc_hd__inv_2_25/A sky130_fd_sc_hd__xor2_2_0/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1737 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_36 sky130_fd_sc_hd__inv_2_36/A sky130_fd_sc_hd__inv_2_36/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_440 sky130_fd_sc_hd__dfxtp_1_440/Q sky130_fd_sc_hd__dfxtp_1_446/CLK
+ sky130_fd_sc_hd__nor2b_1_107/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1748 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_47 sky130_fd_sc_hd__inv_2_47/A sky130_fd_sc_hd__inv_2_47/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_451 sky130_fd_sc_hd__dfxtp_1_451/Q sky130_fd_sc_hd__dfxtp_1_451/CLK
+ sky130_fd_sc_hd__nor2b_1_96/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1759 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_58 sky130_fd_sc_hd__inv_2_58/A sky130_fd_sc_hd__inv_2_58/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_462 sky130_fd_sc_hd__xnor2_1_306/B sky130_fd_sc_hd__dfxtp_1_515/CLK
+ sky130_fd_sc_hd__and2_0_362/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_69 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_473 sky130_fd_sc_hd__dfxtp_1_473/Q sky130_fd_sc_hd__dfxtp_1_479/CLK
+ sky130_fd_sc_hd__and2_0_381/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_484 sky130_fd_sc_hd__buf_8_75/A sky130_fd_sc_hd__dfxtp_1_489/CLK
+ sky130_fd_sc_hd__and2_0_363/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_2_4 sky130_fd_sc_hd__nand2_2_4/Y sky130_fd_sc_hd__nand2_2_4/A
+ sky130_fd_sc_hd__nand2_2_4/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__dfxtp_1_495 la_data_out[44] sky130_fd_sc_hd__dfxtp_1_498/CLK sky130_fd_sc_hd__and2_0_376/X
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2b_1_10 sky130_fd_sc_hd__nand2b_1_10/Y sky130_fd_sc_hd__xnor2_1_71/Y
+ sky130_fd_sc_hd__xnor2_1_68/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__nand2b_1_21 sky130_fd_sc_hd__nand2b_1_21/Y sky130_fd_sc_hd__and3_4_25/C
+ sky130_fd_sc_hd__and3_4_25/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a222oi_1_120 vccd1 vssd1 sky130_fd_sc_hd__and3_4_6/X sky130_fd_sc_hd__buf_4_6/X
+ sky130_fd_sc_hd__buf_4_1/X sky130_fd_sc_hd__nor2_1_72/Y sky130_fd_sc_hd__nor2_2_5/A
+ sky130_fd_sc_hd__o21ai_1_258/B1 sky130_fd_sc_hd__nor2b_1_6/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2b_1_32 sky130_fd_sc_hd__buf_2_143/A sky130_fd_sc_hd__nand2_2_14/A
+ sky130_fd_sc_hd__dfxtp_1_0/Q vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a222oi_1_131 vccd1 vssd1 sky130_fd_sc_hd__and3_4_7/X sky130_fd_sc_hd__buf_4_1/X
+ sky130_fd_sc_hd__nor2_2_5/A sky130_fd_sc_hd__nor2_2_7/Y sky130_fd_sc_hd__nor2_2_5/B
+ sky130_fd_sc_hd__o21ai_1_272/B1 sky130_fd_sc_hd__nor2b_2_1/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_142 vccd1 vssd1 sky130_fd_sc_hd__and3_4_8/X sky130_fd_sc_hd__nor2_2_5/B
+ sky130_fd_sc_hd__nor2_2_4/B sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__buf_2_4/X
+ sky130_fd_sc_hd__o21ai_1_287/B1 sky130_fd_sc_hd__nor2b_2_2/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_153 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__buf_4_3/X sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__o21ai_1_299/B1 sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_301 sky130_fd_sc_hd__fa_2_294/B sky130_fd_sc_hd__fa_2_304/A
+ sky130_fd_sc_hd__fa_2_301/A sky130_fd_sc_hd__fa_2_301/B sky130_fd_sc_hd__fa_2_301/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_164 vccd1 vssd1 sky130_fd_sc_hd__and3_4_1/X sky130_fd_sc_hd__nor2_2_5/A
+ sky130_fd_sc_hd__nor2_2_5/B sky130_fd_sc_hd__nor2_2_9/Y sky130_fd_sc_hd__nor2_2_4/B
+ sky130_fd_sc_hd__o21ai_1_315/B1 sky130_fd_sc_hd__and2b_4_3/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_312 sky130_fd_sc_hd__fa_2_305/A sky130_fd_sc_hd__fa_2_311/B
+ sky130_fd_sc_hd__fa_2_312/A sky130_fd_sc_hd__fa_2_312/B sky130_fd_sc_hd__fa_2_312/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_175 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__buf_6_1/X sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__o21ai_1_330/B1 sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_323 sky130_fd_sc_hd__fa_2_317/B sky130_fd_sc_hd__fa_2_325/CIN
+ sky130_fd_sc_hd__fa_2_323/A sky130_fd_sc_hd__fa_2_323/B sky130_fd_sc_hd__fa_2_323/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_186 vccd1 vssd1 sky130_fd_sc_hd__and3_4_2/X sky130_fd_sc_hd__and2_0_25/A
+ sky130_fd_sc_hd__nor2_2_5/A sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__nor2_2_5/B
+ sky130_fd_sc_hd__o21ai_1_345/B1 sky130_fd_sc_hd__and2b_4_4/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_334 sky130_fd_sc_hd__fa_2_329/CIN sky130_fd_sc_hd__fa_2_341/A
+ sky130_fd_sc_hd__fa_2_334/A sky130_fd_sc_hd__fa_2_334/B sky130_fd_sc_hd__fa_2_339/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_197 vccd1 vssd1 sky130_fd_sc_hd__and3_4_2/X sky130_fd_sc_hd__buf_2_32/X
+ sky130_fd_sc_hd__buf_8_0/X sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__buf_4_6/X
+ sky130_fd_sc_hd__o21ai_1_362/B1 sky130_fd_sc_hd__and2b_4_4/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_345 sky130_fd_sc_hd__fa_2_341/B sky130_fd_sc_hd__fa_2_348/CIN
+ sky130_fd_sc_hd__fa_2_345/A sky130_fd_sc_hd__fa_2_345/B sky130_fd_sc_hd__fa_2_345/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_356 sky130_fd_sc_hd__fa_2_352/CIN sky130_fd_sc_hd__fa_2_362/A
+ sky130_fd_sc_hd__fa_2_356/A sky130_fd_sc_hd__fa_2_356/B sky130_fd_sc_hd__fa_2_361/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_367 sky130_fd_sc_hd__fa_2_356/B sky130_fd_sc_hd__fa_2_367/SUM
+ sky130_fd_sc_hd__fa_2_367/A sky130_fd_sc_hd__fa_2_367/B sky130_fd_sc_hd__xor2_1_539/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_378 sky130_fd_sc_hd__fa_2_374/B sky130_fd_sc_hd__fah_1_7/CI
+ sky130_fd_sc_hd__fa_2_378/A sky130_fd_sc_hd__fa_2_378/B sky130_fd_sc_hd__fa_2_378/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_19 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_4_1/Y
+ sky130_fd_sc_hd__dfxtp_1_177/CLK sky130_fd_sc_hd__o21ai_2_1/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_389 sky130_fd_sc_hd__fa_2_383/CIN sky130_fd_sc_hd__fa_2_391/A
+ sky130_fd_sc_hd__fa_2_389/A sky130_fd_sc_hd__fa_2_389/B sky130_fd_sc_hd__xor2_1_574/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_8_50 sky130_fd_sc_hd__clkinv_8_50/Y sky130_fd_sc_hd__clkinv_8_76/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_61 sky130_fd_sc_hd__clkinv_8_61/Y sky130_fd_sc_hd__clkinv_8_61/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_72 sky130_fd_sc_hd__clkinv_8_73/A sky130_fd_sc_hd__clkinv_8_72/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_83 sky130_fd_sc_hd__clkinv_8_83/Y sky130_fd_sc_hd__clkinv_8_83/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_70 sky130_fd_sc_hd__buf_8_15/X sky130_fd_sc_hd__buf_12_70/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_81 sky130_fd_sc_hd__buf_12_81/A sky130_fd_sc_hd__buf_12_81/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_92 sky130_fd_sc_hd__buf_8_146/X sky130_fd_sc_hd__buf_12_92/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_19 sky130_fd_sc_hd__nor2_4_0/Y sky130_fd_sc_hd__nor2_2_0/Y
+ sky130_fd_sc_hd__dfxtp_1_331/Q sky130_fd_sc_hd__nor2_1_239/A sky130_fd_sc_hd__nand2_2_4/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_306 sky130_fd_sc_hd__buf_12_83/X sky130_fd_sc_hd__buf_12_507/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_317 sky130_fd_sc_hd__buf_12_317/A sky130_fd_sc_hd__buf_12_500/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_328 sky130_fd_sc_hd__buf_12_8/X sky130_fd_sc_hd__buf_12_580/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_339 sky130_fd_sc_hd__buf_12_339/A sky130_fd_sc_hd__buf_12_608/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_209 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__nor2b_2_4/Y sky130_fd_sc_hd__nor2_2_20/Y sky130_fd_sc_hd__a22oi_1_209/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_506 sky130_fd_sc_hd__xnor2_1_66/A sky130_fd_sc_hd__nand2_1_483/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_517 sky130_fd_sc_hd__xor2_1_425/B sky130_fd_sc_hd__a21oi_1_104/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_528 sky130_fd_sc_hd__nor2_1_168/A sky130_fd_sc_hd__nand2_1_532/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_539 sky130_fd_sc_hd__o21ai_1_709/A2 sky130_fd_sc_hd__xnor2_1_142/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_20 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_20/Y
+ sky130_fd_sc_hd__nor2_1_20/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_31 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_31/Y
+ sky130_fd_sc_hd__nor2_1_31/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_42 sky130_fd_sc_hd__nor2_1_42/B sky130_fd_sc_hd__nor2_1_42/Y
+ sky130_fd_sc_hd__nor2_1_42/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_53 sky130_fd_sc_hd__nor2_1_53/B sky130_fd_sc_hd__nor2_1_53/Y
+ sky130_fd_sc_hd__nor2_1_53/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_64 sky130_fd_sc_hd__nor2_1_67/A sky130_fd_sc_hd__nor2_1_64/Y
+ sky130_fd_sc_hd__nor2_1_64/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_19 sky130_fd_sc_hd__buf_8_98/A sky130_fd_sc_hd__inv_2_144/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_75 sky130_fd_sc_hd__nor2_2_10/Y sky130_fd_sc_hd__nor2_1_75/Y
+ sky130_fd_sc_hd__nor2_1_77/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_86 sky130_fd_sc_hd__nor2_1_86/B sky130_fd_sc_hd__nor2_1_86/Y
+ sky130_fd_sc_hd__nor2_1_86/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_97 sky130_fd_sc_hd__nor2_1_97/B sky130_fd_sc_hd__nor2_1_97/Y
+ sky130_fd_sc_hd__nor2_1_97/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_12_502 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_513 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_524 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_535 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_546 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_430 sky130_fd_sc_hd__xnor2_1_104/A sky130_fd_sc_hd__nand2_1_431/Y
+ sky130_fd_sc_hd__nand2_1_430/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_557 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_441 sky130_fd_sc_hd__xor2_1_384/B sky130_fd_sc_hd__nand2_1_442/Y
+ sky130_fd_sc_hd__nand2_1_441/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_568 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_452 sky130_fd_sc_hd__xnor2_1_64/B sky130_fd_sc_hd__nand2_1_453/Y
+ sky130_fd_sc_hd__nand2_1_452/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_579 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_463 sky130_fd_sc_hd__nand2_1_463/Y sky130_fd_sc_hd__buf_4_0/X
+ sky130_fd_sc_hd__buf_2_23/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_474 sky130_fd_sc_hd__nand2_1_474/Y sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__buf_4_7/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_485 sky130_fd_sc_hd__nand2_1_485/Y sky130_fd_sc_hd__a211o_1_2/X
+ sky130_fd_sc_hd__xor2_1_420/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_496 sky130_fd_sc_hd__nand2_1_496/Y sky130_fd_sc_hd__nor2_1_186/Y
+ sky130_fd_sc_hd__or2_0_72/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_10 sky130_fd_sc_hd__and3_4_14/C sky130_fd_sc_hd__nor2b_1_10/Y
+ sky130_fd_sc_hd__and3_4_14/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_21 sky130_fd_sc_hd__or2_0_84/A sky130_fd_sc_hd__or2_0_97/A
+ sky130_fd_sc_hd__xnor2_2_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_32 sky130_fd_sc_hd__fa_2_418/A sky130_fd_sc_hd__fa_2_467/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_43 sky130_fd_sc_hd__mux2_2_20/X sky130_fd_sc_hd__nor2b_1_43/Y
+ sky130_fd_sc_hd__buf_2_214/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1010 sky130_fd_sc_hd__clkinv_1_1011/A sky130_fd_sc_hd__inv_4_1/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_54 sky130_fd_sc_hd__mux2_2_37/X sky130_fd_sc_hd__fa_2_478/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1021 sky130_fd_sc_hd__buf_6_20/A sky130_fd_sc_hd__inv_2_158/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_65 sky130_fd_sc_hd__or2_0_79/B sky130_fd_sc_hd__nor2b_1_65/Y
+ sky130_fd_sc_hd__mux2_4_5/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1032 sky130_fd_sc_hd__buf_8_149/A sky130_fd_sc_hd__inv_2_161/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_76 sky130_fd_sc_hd__or2_0_81/A sky130_fd_sc_hd__fa_2_489/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1043 sky130_fd_sc_hd__clkinv_1_1044/A sky130_fd_sc_hd__clkinv_1_926/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1501 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_87 la_data_out[67] sky130_fd_sc_hd__ha_2_18/A sky130_fd_sc_hd__mux2_4_5/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1054 sky130_fd_sc_hd__inv_2_187/A sky130_fd_sc_hd__clkbuf_1_271/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1512 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_98 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_98/Y
+ sky130_fd_sc_hd__nor2b_1_98/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1065 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__buf_8_157/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_6 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_6/B sky130_fd_sc_hd__xnor2_1_6/Y
+ sky130_fd_sc_hd__xnor2_1_6/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_1523 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1076 sky130_fd_sc_hd__a22o_1_62/B2 la_data_out[39] vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1534 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1087 sky130_fd_sc_hd__nand2_1_861/B sky130_fd_sc_hd__ha_2_54/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1545 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1098 sky130_fd_sc_hd__o21ai_1_926/A2 wbs_adr_i[4] vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1556 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1567 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_270 sky130_fd_sc_hd__fa_2_56/A sky130_fd_sc_hd__dfxtp_1_275/CLK
+ sky130_fd_sc_hd__and2_0_97/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1578 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_281 sky130_fd_sc_hd__dfxtp_1_281/Q sky130_fd_sc_hd__dfxtp_1_2/CLK
+ sky130_fd_sc_hd__and2_0_257/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1589 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_292 sky130_fd_sc_hd__dfxtp_1_292/Q sky130_fd_sc_hd__clkinv_8_6/Y
+ sky130_fd_sc_hd__and2_0_268/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__mux2_4_2 sky130_fd_sc_hd__mux2_4_2/X sky130_fd_sc_hd__mux2_8_1/S
+ sky130_fd_sc_hd__buf_4_14/X sky130_fd_sc_hd__mux2_4_2/A1 vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__mux2_4
Xsky130_fd_sc_hd__o22ai_1_1 sky130_fd_sc_hd__o22ai_1_1/A2 sky130_fd_sc_hd__o22ai_1_1/B1
+ sky130_fd_sc_hd__o22ai_1_1/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__o22ai_1_9/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_120 sky130_fd_sc_hd__fa_2_117/A sky130_fd_sc_hd__fa_2_123/A
+ sky130_fd_sc_hd__fa_2_120/A sky130_fd_sc_hd__fa_2_120/B sky130_fd_sc_hd__fa_2_120/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_131 sky130_fd_sc_hd__fa_2_129/A sky130_fd_sc_hd__fa_2_132/CIN
+ sky130_fd_sc_hd__fa_2_131/A sky130_fd_sc_hd__fa_2_131/B sky130_fd_sc_hd__fa_2_131/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_142 sky130_fd_sc_hd__xor2_1_213/B sky130_fd_sc_hd__or2_0_27/B
+ sky130_fd_sc_hd__fa_2_142/A sky130_fd_sc_hd__fa_2_142/B sky130_fd_sc_hd__fa_2_147/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_153 sky130_fd_sc_hd__fa_2_143/A sky130_fd_sc_hd__fa_2_156/CIN
+ sky130_fd_sc_hd__fa_2_153/A sky130_fd_sc_hd__fa_2_153/B sky130_fd_sc_hd__xor2_1_240/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_164 sky130_fd_sc_hd__fa_2_153/A sky130_fd_sc_hd__fa_2_163/B
+ sky130_fd_sc_hd__fa_2_164/A sky130_fd_sc_hd__fa_2_164/B sky130_fd_sc_hd__xor2_1_249/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and3_4_3 sky130_fd_sc_hd__and3_4_3/A sky130_fd_sc_hd__and3_4_3/B
+ sky130_fd_sc_hd__and3_4_3/C sky130_fd_sc_hd__and3_4_3/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__fa_2_175 sky130_fd_sc_hd__fa_2_160/B sky130_fd_sc_hd__fa_2_177/CIN
+ sky130_fd_sc_hd__fa_2_175/A sky130_fd_sc_hd__fa_2_175/B sky130_fd_sc_hd__fa_2_176/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_186 sky130_fd_sc_hd__fa_2_183/CIN sky130_fd_sc_hd__fa_2_193/A
+ sky130_fd_sc_hd__fa_2_186/A sky130_fd_sc_hd__fa_2_186/B sky130_fd_sc_hd__fa_2_190/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_197 sky130_fd_sc_hd__fa_2_193/B sky130_fd_sc_hd__fa_2_201/CIN
+ sky130_fd_sc_hd__fa_2_197/A sky130_fd_sc_hd__fa_2_197/B sky130_fd_sc_hd__fa_2_197/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o22ai_1_30 sky130_fd_sc_hd__o22ai_1_35/B1 sky130_fd_sc_hd__o21ai_1_5/A2
+ sky130_fd_sc_hd__o22ai_1_30/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__inv_4_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_41 sky130_fd_sc_hd__nor2_1_26/A sky130_fd_sc_hd__o22ai_1_41/B1
+ sky130_fd_sc_hd__o22ai_1_41/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_52 sky130_fd_sc_hd__nor2_1_15/A sky130_fd_sc_hd__o22ai_1_52/B1
+ sky130_fd_sc_hd__o22ai_1_52/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_170 vccd1 vssd1 la_data_out[52] sky130_fd_sc_hd__ha_2_36/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_63 sky130_fd_sc_hd__nor2_1_6/A sky130_fd_sc_hd__o22ai_1_2/A2
+ sky130_fd_sc_hd__o22ai_1_63/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_181 vccd1 vssd1 sky130_fd_sc_hd__buf_2_181/X sky130_fd_sc_hd__inv_2_196/Y
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_74 sky130_fd_sc_hd__xnor2_1_224/Y sky130_fd_sc_hd__xnor2_1_233/Y
+ sky130_fd_sc_hd__ha_2_12/B sky130_fd_sc_hd__inv_2_65/Y sky130_fd_sc_hd__o22ai_1_99/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_192 vccd1 vssd1 sky130_fd_sc_hd__buf_2_192/X sky130_fd_sc_hd__buf_2_192/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_85 sky130_fd_sc_hd__xnor2_2_6/Y sky130_fd_sc_hd__xnor2_1_234/Y
+ sky130_fd_sc_hd__ha_2_14/A sky130_fd_sc_hd__xnor2_1_237/Y sky130_fd_sc_hd__o22ai_1_98/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_96 sky130_fd_sc_hd__xnor2_2_4/Y sky130_fd_sc_hd__xnor2_1_252/Y
+ sky130_fd_sc_hd__o22ai_1_96/Y sky130_fd_sc_hd__xnor2_1_244/Y sky130_fd_sc_hd__o22ai_1_96/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_4_10 vccd1 vssd1 sky130_fd_sc_hd__buf_4_10/X sky130_fd_sc_hd__buf_4_10/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_21 vccd1 vssd1 sky130_fd_sc_hd__buf_4_21/X sky130_fd_sc_hd__buf_4_21/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_32 vccd1 vssd1 sky130_fd_sc_hd__buf_4_32/X sky130_fd_sc_hd__buf_8_18/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_12_103 sky130_fd_sc_hd__buf_8_109/X sky130_fd_sc_hd__buf_12_298/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_114 sky130_fd_sc_hd__buf_8_104/X sky130_fd_sc_hd__buf_12_359/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_125 sky130_fd_sc_hd__buf_8_52/X sky130_fd_sc_hd__buf_12_432/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_136 sky130_fd_sc_hd__buf_12_40/X sky130_fd_sc_hd__buf_12_305/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_147 sky130_fd_sc_hd__buf_8_137/X sky130_fd_sc_hd__buf_12_450/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_70 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_29/A1 sky130_fd_sc_hd__clkbuf_1_70/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_158 sky130_fd_sc_hd__buf_12_12/X sky130_fd_sc_hd__buf_12_158/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_81 vssd1 vccd1 sky130_fd_sc_hd__mux2_4_3/A1 sky130_fd_sc_hd__clkbuf_1_81/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_169 sky130_fd_sc_hd__buf_12_27/X sky130_fd_sc_hd__buf_12_332/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_92 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_45/A1 sky130_fd_sc_hd__clkbuf_1_92/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_4_6 sky130_fd_sc_hd__nor2_2_4/B sky130_fd_sc_hd__buf_2_31/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_1_303 sky130_fd_sc_hd__nand3_1_3/C sky130_fd_sc_hd__ha_2_5/COUT
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_314 sky130_fd_sc_hd__nor2_1_45/B sky130_fd_sc_hd__nand2_1_172/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_325 sky130_fd_sc_hd__o21ai_1_209/A2 sky130_fd_sc_hd__o21ai_1_221/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_336 sky130_fd_sc_hd__a21oi_1_44/B1 sky130_fd_sc_hd__nor2_1_59/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_347 sky130_fd_sc_hd__nor2_1_63/B sky130_fd_sc_hd__nand2_1_216/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_358 sky130_fd_sc_hd__o21ai_1_300/B1 sky130_fd_sc_hd__nand2_1_229/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_369 sky130_fd_sc_hd__a21oi_1_54/B1 sky130_fd_sc_hd__nand2_1_264/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_200 la_data_out[56] sky130_fd_sc_hd__ha_2_58/COUT sky130_fd_sc_hd__a21oi_1_200/Y
+ sky130_fd_sc_hd__o21ai_1_922/A2 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__or2_0_50 sky130_fd_sc_hd__or2_0_50/A sky130_fd_sc_hd__or2_0_50/X
+ sky130_fd_sc_hd__or2_0_50/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_61 sky130_fd_sc_hd__or2_0_61/A sky130_fd_sc_hd__or2_0_61/X
+ sky130_fd_sc_hd__or2_0_61/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_72 sky130_fd_sc_hd__or2_0_72/A sky130_fd_sc_hd__or2_0_72/X
+ sky130_fd_sc_hd__or2_0_72/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__clkinv_4_6 sky130_fd_sc_hd__clkinv_4_6/A sky130_fd_sc_hd__clkinv_4_6/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__or2_0_83 sky130_fd_sc_hd__or2_0_83/A sky130_fd_sc_hd__or2_0_83/X
+ la_data_out[67] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_94 sky130_fd_sc_hd__or2_0_94/A sky130_fd_sc_hd__or2_0_94/X
+ sky130_fd_sc_hd__or2_0_94/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__buf_12_670 sky130_fd_sc_hd__buf_12_670/A sky130_fd_sc_hd__buf_12_670/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_681 sky130_fd_sc_hd__mux2_2_55/X sky130_fd_sc_hd__or2_0_84/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_310 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_321 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_332 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_343 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_354 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_365 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_376 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_260 sky130_fd_sc_hd__nand2_1_260/Y sky130_fd_sc_hd__nor2_1_83/A
+ sky130_fd_sc_hd__nor2_1_83/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_387 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_271 sky130_fd_sc_hd__nand2_1_271/Y sky130_fd_sc_hd__nor2_1_88/A
+ sky130_fd_sc_hd__nor2_1_88/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_398 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_870 sky130_fd_sc_hd__clkinv_1_870/Y sky130_fd_sc_hd__clkinv_4_83/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_282 sky130_fd_sc_hd__nand2_1_282/Y sky130_fd_sc_hd__buf_2_4/X
+ sky130_fd_sc_hd__nor2_2_4/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_881 sky130_fd_sc_hd__clkinv_1_881/Y sky130_fd_sc_hd__clkinv_4_86/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_293 sky130_fd_sc_hd__nand2_1_293/Y sky130_fd_sc_hd__nand2_1_303/Y
+ sky130_fd_sc_hd__nand2_1_297/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_892 sky130_fd_sc_hd__clkinv_1_894/A sky130_fd_sc_hd__buf_2_45/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1320 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1331 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_70 sky130_fd_sc_hd__conb_1_70/LO sky130_fd_sc_hd__conb_1_70/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1342 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_81 sky130_fd_sc_hd__conb_1_81/LO sky130_fd_sc_hd__conb_1_81/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1353 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_92 sky130_fd_sc_hd__conb_1_92/LO sky130_fd_sc_hd__conb_1_92/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1364 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1375 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_806 vssd1 vccd1 sky130_fd_sc_hd__inv_2_49/Y sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__o21ai_1_806/B1 sky130_fd_sc_hd__xor2_1_581/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1386 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_817 vssd1 vccd1 sky130_fd_sc_hd__inv_2_45/Y sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_817/B1 sky130_fd_sc_hd__xor2_1_591/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1397 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_828 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_602/A sky130_fd_sc_hd__nor2_1_203/Y
+ sky130_fd_sc_hd__nand2_1_618/Y sky130_fd_sc_hd__o21ai_1_828/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_839 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_616/B sky130_fd_sc_hd__nor2_1_211/Y
+ sky130_fd_sc_hd__nand2_1_632/Y sky130_fd_sc_hd__o21ai_1_839/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nand2b_2_7 sky130_fd_sc_hd__nor2_4_17/B sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__nor2_4_17/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_2
Xsky130_fd_sc_hd__xor2_1_600 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__fa_2_400/A
+ sky130_fd_sc_hd__xor2_1_600/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_611 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__fa_2_405/A
+ sky130_fd_sc_hd__xor2_1_611/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_622 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__nor2_4_17/B
+ sky130_fd_sc_hd__xor2_1_622/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_633 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__xor2_1_633/X
+ sky130_fd_sc_hd__xor2_1_633/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_644 sky130_fd_sc_hd__xor2_1_644/B sky130_fd_sc_hd__xor2_1_644/X
+ sky130_fd_sc_hd__xor2_1_644/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_655 sky130_fd_sc_hd__xor2_1_655/B sky130_fd_sc_hd__xor2_1_655/X
+ sky130_fd_sc_hd__xor2_1_655/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_666 sky130_fd_sc_hd__xor2_1_666/B sky130_fd_sc_hd__or2_0_92/B
+ sky130_fd_sc_hd__xor2_1_666/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_677 sky130_fd_sc_hd__xor2_1_677/B sky130_fd_sc_hd__xor2_1_677/X
+ sky130_fd_sc_hd__xor2_1_677/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_688 sky130_fd_sc_hd__xor2_1_688/B sky130_fd_sc_hd__xor2_1_688/X
+ sky130_fd_sc_hd__xor2_1_688/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__fa_2_7 sky130_fd_sc_hd__xor3_1_7/B sky130_fd_sc_hd__fa_2_8/CIN sky130_fd_sc_hd__fa_2_7/A
+ sky130_fd_sc_hd__fa_2_7/B sky130_fd_sc_hd__fa_2_7/CIN vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a211o_1_13 vssd1 vccd1 sky130_fd_sc_hd__fa_2_258/A sky130_fd_sc_hd__dfxtp_1_76/Q
+ sky130_fd_sc_hd__nor2_1_17/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_13/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__a211o_1_24 vssd1 vccd1 sky130_fd_sc_hd__fa_2_198/B sky130_fd_sc_hd__dfxtp_1_87/Q
+ sky130_fd_sc_hd__nor2_1_28/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_24/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__clkinv_1_100 io_out[1] sky130_fd_sc_hd__conb_1_42/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_111 io_oeb[28] sky130_fd_sc_hd__conb_1_31/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_122 io_oeb[17] sky130_fd_sc_hd__conb_1_20/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_133 io_oeb[6] sky130_fd_sc_hd__conb_1_9/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_144 sky130_fd_sc_hd__a22oi_1_8/A1 sky130_fd_sc_hd__nor2_1_0/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_155 sky130_fd_sc_hd__nor2_1_32/A sky130_fd_sc_hd__dfxtp_1_155/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_166 sky130_fd_sc_hd__o22ai_1_37/B1 sky130_fd_sc_hd__dfxtp_1_184/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_177 sky130_fd_sc_hd__o22ai_1_23/B1 sky130_fd_sc_hd__dfxtp_1_118/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_9 sky130_fd_sc_hd__inv_4_9/Y sky130_fd_sc_hd__buf_8_9/X vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__a22o_1_13 sky130_fd_sc_hd__inv_2_66/Y sky130_fd_sc_hd__or2_0_88/B
+ sky130_fd_sc_hd__a22o_1_13/X sky130_fd_sc_hd__nor2_1_233/Y sky130_fd_sc_hd__a22o_1_13/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_188 sky130_fd_sc_hd__nor2_1_23/A sky130_fd_sc_hd__dfxtp_1_146/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_199 sky130_fd_sc_hd__o22ai_1_48/B1 sky130_fd_sc_hd__dfxtp_1_174/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_24 sky130_fd_sc_hd__buf_2_63/A sky130_fd_sc_hd__buf_2_99/X
+ sky130_fd_sc_hd__a22o_1_24/X sky130_fd_sc_hd__a22o_1_24/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_35 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__buf_2_110/X
+ sky130_fd_sc_hd__a22o_1_35/X sky130_fd_sc_hd__a22o_1_35/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_46 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__buf_2_121/X
+ sky130_fd_sc_hd__a22o_1_46/X sky130_fd_sc_hd__a22o_1_46/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__o21ai_1_0 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_2/Y sky130_fd_sc_hd__o21ai_2_1/A2
+ sky130_fd_sc_hd__o21ai_2_0/B1 sky130_fd_sc_hd__o21ai_1_0/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a22o_1_57 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__and2_0_356/A
+ sky130_fd_sc_hd__a22o_1_57/X sky130_fd_sc_hd__ha_2_28/SUM sky130_fd_sc_hd__a22o_1_71/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_68 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__buf_2_41/A
+ sky130_fd_sc_hd__a22o_1_68/X sky130_fd_sc_hd__ha_2_37/SUM sky130_fd_sc_hd__a22o_1_71/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_79 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__a22o_1_79/A2
+ sky130_fd_sc_hd__a22o_1_79/X sky130_fd_sc_hd__ha_2_25/SUM sky130_fd_sc_hd__nor2_1_269/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_2_3 sky130_fd_sc_hd__nor2_4_3/A sky130_fd_sc_hd__ha_2_8/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__nor2_1_260 sky130_fd_sc_hd__nor2_1_260/B sky130_fd_sc_hd__nor2_1_260/Y
+ sky130_fd_sc_hd__nor2_1_260/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_271 sky130_fd_sc_hd__nor2_2_0/B sky130_fd_sc_hd__nor2_1_271/Y
+ sky130_fd_sc_hd__nor2_4_0/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_282 sky130_fd_sc_hd__a21o_2_4/A2 sky130_fd_sc_hd__a21o_2_4/B1
+ wbs_adr_i[9] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_12_140 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_151 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_162 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_173 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_184 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_14 sky130_fd_sc_hd__nand2_1_14/Y sky130_fd_sc_hd__nand2_1_14/B
+ sky130_fd_sc_hd__nand2_1_14/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_195 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_25 sky130_fd_sc_hd__nand2_8_3/A sky130_fd_sc_hd__nand2_1_7/B
+ sky130_fd_sc_hd__mux2_2_24/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_230 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_5/B sky130_fd_sc_hd__xnor2_1_230/Y
+ sky130_fd_sc_hd__buf_4_41/X vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_36 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__nand2_1_7/B
+ la_data_out[72] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_241 vssd1 vccd1 la_data_out[77] sky130_fd_sc_hd__xnor2_1_241/Y
+ sky130_fd_sc_hd__or2_1_10/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_47 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__nand2_1_8/B
+ sky130_fd_sc_hd__or2_0_83/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_252 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_5/B sky130_fd_sc_hd__xnor2_1_252/Y
+ la_data_out[67] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_58 sky130_fd_sc_hd__nand2_1_58/Y sky130_fd_sc_hd__nand2_1_58/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_263 vssd1 vccd1 la_data_out[79] sky130_fd_sc_hd__xnor2_1_263/Y
+ sky130_fd_sc_hd__mux2_2_31/X vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_69 sky130_fd_sc_hd__nand2_1_69/Y sky130_fd_sc_hd__nand2_1_69/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_274 vssd1 vccd1 la_data_out[77] sky130_fd_sc_hd__xnor2_1_274/Y
+ sky130_fd_sc_hd__or2_0_78/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_285 vssd1 vccd1 la_data_out[85] sky130_fd_sc_hd__xnor2_1_285/Y
+ sky130_fd_sc_hd__or2_1_10/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_296 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_296/B sky130_fd_sc_hd__xnor2_1_296/Y
+ sky130_fd_sc_hd__xnor2_1_296/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_1150 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1161 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1172 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_603 vssd1 vccd1 sky130_fd_sc_hd__buf_2_10/X sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_603/B1 sky130_fd_sc_hd__xor2_1_394/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1183 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_614 vssd1 vccd1 sky130_fd_sc_hd__nand2_2_12/Y sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__a22oi_1_210/Y sky130_fd_sc_hd__xor2_1_406/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1194 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_625 vssd1 vccd1 sky130_fd_sc_hd__inv_2_27/Y sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__nand2_1_332/Y sky130_fd_sc_hd__xor2_1_417/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_636 vssd1 vccd1 sky130_fd_sc_hd__xor2_2_2/X sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_636/B1 sky130_fd_sc_hd__xor2_1_583/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_647 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_713/A2 sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__o21ai_1_647/B1 sky130_fd_sc_hd__xor2_1_434/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_658 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_658/A2 sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_658/B1 sky130_fd_sc_hd__xor2_1_443/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_669 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_709/A2 sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_669/B1 sky130_fd_sc_hd__xor2_1_452/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fah_1_1 sky130_fd_sc_hd__fah_1_1/COUT sky130_fd_sc_hd__fah_1_1/B
+ sky130_fd_sc_hd__fah_1_1/A sky130_fd_sc_hd__fa_2_115/A sky130_fd_sc_hd__fah_1_1/CI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__fah_1
Xsky130_fd_sc_hd__xor2_1_430 sky130_fd_sc_hd__fa_2_379/A sky130_fd_sc_hd__xor3_1_23/A
+ sky130_fd_sc_hd__xor2_1_430/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_441 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__xor2_1_441/X
+ sky130_fd_sc_hd__xor2_1_441/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_452 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__fa_2_292/A
+ sky130_fd_sc_hd__xor2_1_452/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_463 sky130_fd_sc_hd__fa_2_338/A sky130_fd_sc_hd__fa_2_304/B
+ sky130_fd_sc_hd__xor2_1_463/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_474 sky130_fd_sc_hd__fa_2_310/A sky130_fd_sc_hd__xor2_1_474/X
+ sky130_fd_sc_hd__xor2_1_474/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_485 sky130_fd_sc_hd__fa_2_357/A sky130_fd_sc_hd__fa_2_321/A
+ sky130_fd_sc_hd__xor2_1_485/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_496 sky130_fd_sc_hd__fah_1_14/A sky130_fd_sc_hd__fa_2_330/A
+ sky130_fd_sc_hd__xor2_1_496/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a222oi_1_505 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__buf_2_20/X
+ sky130_fd_sc_hd__buf_2_21/X sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__o21ai_1_802/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_516 vccd1 vssd1 sky130_fd_sc_hd__and3_4_21/X sky130_fd_sc_hd__buf_2_26/X
+ sky130_fd_sc_hd__buf_2_24/X sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__buf_2_27/X
+ sky130_fd_sc_hd__o21ai_1_813/B1 sky130_fd_sc_hd__and2b_4_12/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__dfxtp_4_3 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_4_3/D sky130_fd_sc_hd__dfxtp_4_3/CLK
+ sky130_fd_sc_hd__or2_0_70/A vssd1 vccd1 sky130_fd_sc_hd__dfxtp_4
Xsky130_fd_sc_hd__a222oi_1_527 vccd1 vssd1 sky130_fd_sc_hd__and3_4_21/X sky130_fd_sc_hd__buf_2_14/A
+ sky130_fd_sc_hd__buf_2_29/X sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__buf_2_30/X
+ sky130_fd_sc_hd__o21ai_1_830/B1 sky130_fd_sc_hd__and2b_4_12/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_538 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__buf_4_6/X
+ sky130_fd_sc_hd__buf_4_1/X sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__buf_4_0/A
+ sky130_fd_sc_hd__o21ai_1_849/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_549 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_421/Q sky130_fd_sc_hd__inv_2_68/Y
+ sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__dfxtp_1_453/Q sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__clkinv_1_746/A sky130_fd_sc_hd__dfxtp_1_389/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nor2b_1_105 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_105/Y
+ sky130_fd_sc_hd__nor2b_1_105/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_116 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_116/Y
+ sky130_fd_sc_hd__nor2b_1_116/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_127 sky130_fd_sc_hd__clkinv_4_46/Y sky130_fd_sc_hd__nor2b_1_127/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_138 sky130_fd_sc_hd__clkinv_4_57/Y sky130_fd_sc_hd__nor2b_1_138/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_149 sky130_fd_sc_hd__clkinv_4_68/Y sky130_fd_sc_hd__nor2b_1_149/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__fah_1_18 sky130_fd_sc_hd__fa_2_447/B sky130_fd_sc_hd__fah_1_18/B
+ sky130_fd_sc_hd__fah_1_18/A sky130_fd_sc_hd__fah_1_17/CI sky130_fd_sc_hd__fah_1_18/CI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__fah_1
Xsky130_fd_sc_hd__buf_6_6 vccd1 vssd1 sky130_fd_sc_hd__buf_6_6/X sky130_fd_sc_hd__buf_6_6/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__clkinv_2_30 sky130_fd_sc_hd__clkinv_2_30/Y sky130_fd_sc_hd__clkinv_2_30/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_41 sky130_fd_sc_hd__inv_2_167/A sky130_fd_sc_hd__inv_8_0/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_52 sky130_fd_sc_hd__inv_2_200/A wbs_dat_i[2] vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__or2_1_1 sky130_fd_sc_hd__or2_1_1/A sky130_fd_sc_hd__or2_1_1/X sky130_fd_sc_hd__or2_1_1/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_1
Xsky130_fd_sc_hd__sdlclkp_4_4 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_4_0/Y
+ sky130_fd_sc_hd__dfxtp_1_62/CLK sky130_fd_sc_hd__o21ai_1_0/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_7 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_7/Y
+ sky130_fd_sc_hd__nor2_1_7/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__o21ai_1_400 vssd1 vccd1 sky130_fd_sc_hd__inv_2_38/Y sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_400/B1 sky130_fd_sc_hd__xor2_1_370/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_411 vssd1 vccd1 sky130_fd_sc_hd__inv_2_39/Y sky130_fd_sc_hd__nand2b_1_9/Y
+ sky130_fd_sc_hd__o21ai_1_411/B1 sky130_fd_sc_hd__xor2_1_222/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_422 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_7/X sky130_fd_sc_hd__nand2_1_340/Y
+ sky130_fd_sc_hd__a21oi_1_73/Y sky130_fd_sc_hd__xnor2_1_70/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_433 vssd1 vccd1 sky130_fd_sc_hd__inv_2_37/Y sky130_fd_sc_hd__nand2b_2_3/Y
+ sky130_fd_sc_hd__o21ai_1_433/B1 sky130_fd_sc_hd__xor2_1_240/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_444 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_444/A2 sky130_fd_sc_hd__nor2_1_116/Y
+ sky130_fd_sc_hd__nand2_1_360/Y sky130_fd_sc_hd__o21ai_1_444/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_455 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_7/X sky130_fd_sc_hd__nand2_1_357/Y
+ sky130_fd_sc_hd__a21oi_1_77/Y sky130_fd_sc_hd__xnor2_1_76/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_466 vssd1 vccd1 sky130_fd_sc_hd__inv_2_38/Y sky130_fd_sc_hd__nand2b_1_9/Y
+ sky130_fd_sc_hd__o21ai_1_466/B1 sky130_fd_sc_hd__xor2_1_269/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_477 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_7/X sky130_fd_sc_hd__nand2_1_368/Y
+ sky130_fd_sc_hd__a21oi_1_79/Y sky130_fd_sc_hd__xnor2_1_80/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_3_4 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__o21ai_1_488 vssd1 vccd1 sky130_fd_sc_hd__inv_2_40/Y sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_488/B1 sky130_fd_sc_hd__xor2_1_288/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_499 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_0/Y sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_499/B1 sky130_fd_sc_hd__xor2_1_299/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_909 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_804 sky130_fd_sc_hd__xor2_1_679/B sky130_fd_sc_hd__nand2_1_805/Y
+ sky130_fd_sc_hd__nand2_1_804/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_815 sky130_fd_sc_hd__nand2_1_815/Y sky130_fd_sc_hd__or2_0_105/A
+ sky130_fd_sc_hd__or2_0_105/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_826 sky130_fd_sc_hd__xnor2_1_299/A sky130_fd_sc_hd__nand2_1_827/Y
+ sky130_fd_sc_hd__or2_0_108/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_837 sky130_fd_sc_hd__nand2_1_837/Y sky130_fd_sc_hd__nor2_1_265/A
+ sky130_fd_sc_hd__nor2_1_265/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_848 sky130_fd_sc_hd__nand2_1_848/Y la_data_out[35] sky130_fd_sc_hd__nand2_1_848/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_859 sky130_fd_sc_hd__nand2_1_859/Y sky130_fd_sc_hd__nand2_1_859/B
+ la_data_out[43] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o21ai_1_15 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_18/B1 sky130_fd_sc_hd__inv_2_53/A
+ sky130_fd_sc_hd__o21ai_1_15/B1 sky130_fd_sc_hd__fa_2_97/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_26 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_7/B1 sky130_fd_sc_hd__nor2_4_4/B
+ sky130_fd_sc_hd__o21ai_1_26/B1 sky130_fd_sc_hd__fa_2_135/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_37 vssd1 vccd1 sky130_fd_sc_hd__inv_2_62/Y sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_37/B1 sky130_fd_sc_hd__o21ai_1_37/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_260 sky130_fd_sc_hd__fa_2_198/A sky130_fd_sc_hd__fa_2_172/B
+ sky130_fd_sc_hd__xor2_1_260/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__o21ai_1_48 vssd1 vccd1 sky130_fd_sc_hd__inv_2_63/Y sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_48/B1 sky130_fd_sc_hd__o21ai_1_48/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_271 sky130_fd_sc_hd__fa_2_198/A sky130_fd_sc_hd__xor2_1_271/X
+ sky130_fd_sc_hd__xor2_1_271/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__o21ai_1_59 vssd1 vccd1 sky130_fd_sc_hd__inv_2_60/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_97/Y sky130_fd_sc_hd__o21ai_1_59/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_282 sky130_fd_sc_hd__fa_2_198/A sky130_fd_sc_hd__fa_2_187/B
+ sky130_fd_sc_hd__xor2_1_282/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_293 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__xor2_1_293/X
+ sky130_fd_sc_hd__xor2_1_293/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_220 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_220/X sky130_fd_sc_hd__clkinv_1_907/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_231 vssd1 vccd1 sky130_fd_sc_hd__buf_12_57/A sky130_fd_sc_hd__clkbuf_4_30/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_302 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__buf_4_4/X sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__o21ai_1_514/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_242 vssd1 vccd1 sky130_fd_sc_hd__buf_12_54/A sky130_fd_sc_hd__clkbuf_4_25/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_313 vccd1 vssd1 sky130_fd_sc_hd__and3_4_15/X sky130_fd_sc_hd__or2_0_52/B
+ sky130_fd_sc_hd__or2_0_53/A sky130_fd_sc_hd__nor2_1_130/Y sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__o21ai_1_528/B1 sky130_fd_sc_hd__nor2b_1_11/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_253 vssd1 vccd1 sky130_fd_sc_hd__buf_12_53/A sky130_fd_sc_hd__clkbuf_1_57/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_2_0 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__dfxtp_2_0/CLK
+ sky130_fd_sc_hd__dfxtp_2_4/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_2
Xsky130_fd_sc_hd__a222oi_1_324 vccd1 vssd1 sky130_fd_sc_hd__and3_4_10/X sky130_fd_sc_hd__buf_2_23/X
+ sky130_fd_sc_hd__buf_2_31/X sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__buf_2_19/X
+ sky130_fd_sc_hd__o21ai_1_542/B1 sky130_fd_sc_hd__and2b_4_7/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_264 vssd1 vccd1 sky130_fd_sc_hd__buf_12_44/A sky130_fd_sc_hd__buf_8_20/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_335 vccd1 vssd1 sky130_fd_sc_hd__and3_4_17/X sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__buf_8_0/X sky130_fd_sc_hd__nor2_2_20/Y sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__o21ai_1_556/B1 sky130_fd_sc_hd__nor2b_2_4/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_275 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_275/X sky130_fd_sc_hd__clkbuf_1_59/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_346 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__and2_0_38/A
+ sky130_fd_sc_hd__and2_0_49/A sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__and2_0_45/A
+ sky130_fd_sc_hd__o21ai_1_400/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_286 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_286/X sky130_fd_sc_hd__clkbuf_1_286/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_357 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__buf_2_19/X
+ sky130_fd_sc_hd__buf_6_5/X sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__o21ai_1_590/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_297 vssd1 vccd1 sky130_fd_sc_hd__bufinv_16_0/A sky130_fd_sc_hd__clkbuf_1_297/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_368 vccd1 vssd1 sky130_fd_sc_hd__and3_4_11/X sky130_fd_sc_hd__or2_0_52/B
+ sky130_fd_sc_hd__or2_0_53/A sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__o21ai_1_610/B1 sky130_fd_sc_hd__and2b_4_8/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_379 vccd1 vssd1 sky130_fd_sc_hd__and3_4_20/X sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__buf_4_5/X sky130_fd_sc_hd__nor2_4_16/Y sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__o21ai_1_639/B1 sky130_fd_sc_hd__and2b_4_11/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__buf_4_3 vccd1 vssd1 sky130_fd_sc_hd__buf_4_3/X sky130_fd_sc_hd__buf_4_3/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__and2_0_240 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_58/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_50/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_251 vccd1 vssd1 sky130_fd_sc_hd__and2_0_251/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_251/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_262 vccd1 vssd1 sky130_fd_sc_hd__and2_0_262/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__xor2_1_647/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_273 vccd1 vssd1 sky130_fd_sc_hd__and2_0_273/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__and2_0_273/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_284 vccd1 vssd1 sky130_fd_sc_hd__and2_0_284/X sky130_fd_sc_hd__and2_0_284/B
+ sky130_fd_sc_hd__or2_0_84/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__a21oi_2_14 sky130_fd_sc_hd__a21oi_2_14/B1 sky130_fd_sc_hd__or2_1_8/X
+ sky130_fd_sc_hd__o21ai_2_12/Y sky130_fd_sc_hd__xor2_1_447/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_2
Xsky130_fd_sc_hd__and2_0_295 vccd1 vssd1 sky130_fd_sc_hd__and2_0_295/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_16/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__sdlclkp_2_1 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_2_7/Y
+ sky130_fd_sc_hd__dfxtp_1_65/CLK sky130_fd_sc_hd__o21ai_2_0/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__inv_4_3 sky130_fd_sc_hd__inv_4_3/Y sky130_fd_sc_hd__inv_4_3/A vccd1
+ vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__or2_0_108 sky130_fd_sc_hd__or2_0_108/A sky130_fd_sc_hd__or2_0_108/X
+ sky130_fd_sc_hd__or2_0_108/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__o21ai_1_230 vssd1 vccd1 sky130_fd_sc_hd__inv_2_18/Y sky130_fd_sc_hd__nand2b_1_6/Y
+ sky130_fd_sc_hd__a222oi_1_98/Y sky130_fd_sc_hd__xor2_1_55/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_241 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_241/A2 sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__o21ai_1_241/B1 sky130_fd_sc_hd__xor2_1_65/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_252 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_2/X sky130_fd_sc_hd__nand2_1_203/Y
+ sky130_fd_sc_hd__a21oi_1_45/Y sky130_fd_sc_hd__xnor2_1_20/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_263 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_66/Y sky130_fd_sc_hd__nor2_1_64/A
+ sky130_fd_sc_hd__nor2_1_63/Y sky130_fd_sc_hd__o21ai_1_263/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_274 vssd1 vccd1 sky130_fd_sc_hd__nand2_4_4/Y sky130_fd_sc_hd__nand2b_1_5/Y
+ sky130_fd_sc_hd__a22oi_1_194/Y sky130_fd_sc_hd__xor2_1_95/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_285 vssd1 vccd1 sky130_fd_sc_hd__inv_2_21/Y sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__o21ai_1_285/B1 sky130_fd_sc_hd__xor2_1_106/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_296 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_2/X sky130_fd_sc_hd__nand2_1_224/Y
+ sky130_fd_sc_hd__a21oi_1_48/Y sky130_fd_sc_hd__xnor2_1_29/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_706 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_717 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_601 sky130_fd_sc_hd__nand2_1_601/Y sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__nor2_2_10/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_728 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_612 sky130_fd_sc_hd__xor2_1_597/B sky130_fd_sc_hd__nand2_1_613/Y
+ sky130_fd_sc_hd__nand2_1_612/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_739 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_623 sky130_fd_sc_hd__xnor2_2_3/B sky130_fd_sc_hd__nand2_1_624/Y
+ sky130_fd_sc_hd__nand2_1_623/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_634 sky130_fd_sc_hd__nand2_1_634/Y sky130_fd_sc_hd__buf_2_24/X
+ sky130_fd_sc_hd__buf_2_27/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_645 sky130_fd_sc_hd__nand2_1_645/Y sky130_fd_sc_hd__buf_2_30/X
+ sky130_fd_sc_hd__buf_2_26/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_656 sky130_fd_sc_hd__xnor2_1_129/A sky130_fd_sc_hd__nand2_1_657/Y
+ sky130_fd_sc_hd__or2_0_71/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_667 sky130_fd_sc_hd__nand2_1_667/Y sky130_fd_sc_hd__or2_0_74/A
+ sky130_fd_sc_hd__or2_0_74/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_2_3 sky130_fd_sc_hd__nor2_2_19/A sky130_fd_sc_hd__nor2b_2_3/A
+ sky130_fd_sc_hd__nor2b_2_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_2
Xsky130_fd_sc_hd__nand2_1_678 sky130_fd_sc_hd__xnor2_1_192/A sky130_fd_sc_hd__nand2_1_679/Y
+ sky130_fd_sc_hd__or2_1_11/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_689 sky130_fd_sc_hd__nand2_1_689/Y sky130_fd_sc_hd__mux2_2_24/X
+ sky130_fd_sc_hd__mux2_2_38/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_1705 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1716 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_15 sky130_fd_sc_hd__inv_2_15/A sky130_fd_sc_hd__inv_2_15/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__decap_12_1727 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_26 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__inv_2_26/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_430 sky130_fd_sc_hd__dfxtp_1_430/Q sky130_fd_sc_hd__clkinv_4_9/Y
+ sky130_fd_sc_hd__nor2b_1_117/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1738 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_37 sky130_fd_sc_hd__inv_2_37/A sky130_fd_sc_hd__inv_2_37/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_441 sky130_fd_sc_hd__dfxtp_1_441/Q sky130_fd_sc_hd__dfxtp_1_446/CLK
+ sky130_fd_sc_hd__nor2b_1_106/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1749 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_48 sky130_fd_sc_hd__inv_2_48/A sky130_fd_sc_hd__inv_2_48/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_452 sky130_fd_sc_hd__dfxtp_1_452/Q sky130_fd_sc_hd__dfxtp_1_459/CLK
+ sky130_fd_sc_hd__nor2b_1_95/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_59 sky130_fd_sc_hd__inv_2_59/A sky130_fd_sc_hd__inv_2_59/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_463 sky130_fd_sc_hd__ha_2_48/B sky130_fd_sc_hd__dfxtp_1_520/CLK
+ sky130_fd_sc_hd__and2_0_361/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_474 sky130_fd_sc_hd__ha_2_24/A sky130_fd_sc_hd__dfxtp_1_479/CLK
+ sky130_fd_sc_hd__and2_0_382/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_485 sky130_fd_sc_hd__ha_2_36/A sky130_fd_sc_hd__dfxtp_1_489/CLK
+ sky130_fd_sc_hd__and2_0_377/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_2_5 sky130_fd_sc_hd__nand2_2_5/Y sky130_fd_sc_hd__nand2_2_5/A
+ sky130_fd_sc_hd__nand2_2_5/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__dfxtp_1_496 la_data_out[45] sky130_fd_sc_hd__dfxtp_1_498/CLK sky130_fd_sc_hd__and2_0_365/X
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2b_1_11 sky130_fd_sc_hd__nand2b_1_11/Y sky130_fd_sc_hd__and3_1_1/C
+ sky130_fd_sc_hd__and3_1_1/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a222oi_1_110 vccd1 vssd1 sky130_fd_sc_hd__and3_4_5/X sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__buf_8_0/X sky130_fd_sc_hd__nor2_1_68/Y sky130_fd_sc_hd__buf_4_6/X
+ sky130_fd_sc_hd__o21ai_1_245/B1 sky130_fd_sc_hd__nor2b_1_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2b_1_22 sky130_fd_sc_hd__o22ai_1_78/A1 sky130_fd_sc_hd__or2_0_84/A
+ la_data_out[85] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a222oi_1_121 vccd1 vssd1 sky130_fd_sc_hd__and3_4_7/X sky130_fd_sc_hd__nor2_2_5/B
+ sky130_fd_sc_hd__nor2_2_4/B sky130_fd_sc_hd__nor2_2_7/Y sky130_fd_sc_hd__buf_2_4/X
+ sky130_fd_sc_hd__o21ai_1_259/B1 sky130_fd_sc_hd__nor2b_2_1/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2b_1_33 sky130_fd_sc_hd__nand2b_1_33/Y sky130_fd_sc_hd__ha_2_50/SUM
+ la_data_out[44] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a222oi_1_132 vccd1 vssd1 sky130_fd_sc_hd__and3_4_6/X sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__buf_8_0/X sky130_fd_sc_hd__nor2_1_72/Y sky130_fd_sc_hd__buf_4_6/X
+ sky130_fd_sc_hd__o21ai_1_273/B1 sky130_fd_sc_hd__nor2b_1_6/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_143 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__nor2_1_73/B sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__o21ai_1_288/B1 sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_154 vccd1 vssd1 sky130_fd_sc_hd__and3_4_8/X sky130_fd_sc_hd__and2_0_25/A
+ sky130_fd_sc_hd__nor2_2_5/A sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__nor2_2_5/B
+ sky130_fd_sc_hd__o21ai_1_301/B1 sky130_fd_sc_hd__nor2b_2_2/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_302 sky130_fd_sc_hd__fa_2_298/B sky130_fd_sc_hd__fa_2_308/B
+ sky130_fd_sc_hd__fa_2_302/A sky130_fd_sc_hd__fa_2_302/B sky130_fd_sc_hd__xor2_1_458/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_165 vccd1 vssd1 sky130_fd_sc_hd__and3_4_2/X sky130_fd_sc_hd__buf_2_4/A
+ sky130_fd_sc_hd__buf_6_5/X sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__o21ai_1_316/B1 sky130_fd_sc_hd__and2b_4_4/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_313 sky130_fd_sc_hd__fa_2_306/A sky130_fd_sc_hd__fa_2_314/B
+ sky130_fd_sc_hd__fa_2_313/A sky130_fd_sc_hd__fa_2_313/B sky130_fd_sc_hd__xor2_1_477/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_176 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__nor2_2_10/B sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__buf_6_4/X
+ sky130_fd_sc_hd__o21ai_1_331/B1 sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_324 sky130_fd_sc_hd__fa_2_317/A sky130_fd_sc_hd__fa_2_325/A
+ sky130_fd_sc_hd__fa_2_324/A sky130_fd_sc_hd__fa_2_324/B sky130_fd_sc_hd__fa_2_324/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_187 vccd1 vssd1 sky130_fd_sc_hd__and3_4_1/X sky130_fd_sc_hd__buf_2_32/X
+ sky130_fd_sc_hd__buf_8_0/X sky130_fd_sc_hd__nor2_2_9/Y sky130_fd_sc_hd__buf_4_6/X
+ sky130_fd_sc_hd__o21ai_1_346/B1 sky130_fd_sc_hd__and2b_4_3/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_335 sky130_fd_sc_hd__fa_2_328/CIN sky130_fd_sc_hd__fa_2_334/A
+ sky130_fd_sc_hd__fa_2_335/A sky130_fd_sc_hd__fa_2_335/B sky130_fd_sc_hd__xor2_1_506/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_198 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__nor2_2_4/B
+ sky130_fd_sc_hd__buf_2_4/A sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__o21ai_1_364/B1 sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_346 sky130_fd_sc_hd__fa_2_340/CIN sky130_fd_sc_hd__fa_2_343/B
+ sky130_fd_sc_hd__fa_2_346/A sky130_fd_sc_hd__fa_2_346/B sky130_fd_sc_hd__xor2_1_516/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_357 sky130_fd_sc_hd__fa_2_354/CIN sky130_fd_sc_hd__fa_2_360/A
+ sky130_fd_sc_hd__fa_2_357/A sky130_fd_sc_hd__fa_2_357/B sky130_fd_sc_hd__xor2_1_529/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_368 sky130_fd_sc_hd__nor2_2_26/A sky130_fd_sc_hd__or2_1_4/B
+ sky130_fd_sc_hd__fa_2_368/A sky130_fd_sc_hd__fa_2_368/B sky130_fd_sc_hd__fa_2_368/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_379 sky130_fd_sc_hd__fa_2_372/CIN sky130_fd_sc_hd__fa_2_376/A
+ sky130_fd_sc_hd__fa_2_379/A sky130_fd_sc_hd__fa_2_379/B sky130_fd_sc_hd__xor2_1_556/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_8_40 sky130_fd_sc_hd__clkinv_8_40/Y sky130_fd_sc_hd__clkinv_8_40/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_51 sky130_fd_sc_hd__clkinv_8_69/A sky130_fd_sc_hd__clkinv_8_90/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_62 sky130_fd_sc_hd__clkinv_8_63/A sky130_fd_sc_hd__clkinv_8_62/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_73 sky130_fd_sc_hd__clkinv_8_73/Y sky130_fd_sc_hd__clkinv_8_73/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_84 sky130_fd_sc_hd__clkinv_8_85/A sky130_fd_sc_hd__clkinv_8_84/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_60 sky130_fd_sc_hd__inv_2_180/Y sky130_fd_sc_hd__buf_12_60/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_71 sky130_fd_sc_hd__buf_8_59/X sky130_fd_sc_hd__buf_12_71/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_82 sky130_fd_sc_hd__buf_8_145/X sky130_fd_sc_hd__buf_12_82/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_93 sky130_fd_sc_hd__buf_8_71/X sky130_fd_sc_hd__buf_12_93/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_2_0 vccd1 vssd1 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__buf_2_0/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_12_307 sky130_fd_sc_hd__buf_12_307/A sky130_fd_sc_hd__buf_12_307/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_318 sky130_fd_sc_hd__buf_12_318/A sky130_fd_sc_hd__buf_12_639/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_329 sky130_fd_sc_hd__buf_12_329/A sky130_fd_sc_hd__buf_12_529/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__inv_2_0 sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__inv_2_0/Y vccd1
+ vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__clkinv_1_507 sky130_fd_sc_hd__nand2_1_484/A sky130_fd_sc_hd__nor2_1_162/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_518 sky130_fd_sc_hd__clkinv_1_518/Y sky130_fd_sc_hd__nand2_1_512/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_529 sky130_fd_sc_hd__a21oi_2_14/B1 sky130_fd_sc_hd__nand2_1_523/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_10 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_10/Y
+ sky130_fd_sc_hd__nor2_1_10/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_21 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_21/Y
+ sky130_fd_sc_hd__nor2_1_21/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_32 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_32/Y
+ sky130_fd_sc_hd__nor2_1_32/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_43 sky130_fd_sc_hd__nor2_1_43/B sky130_fd_sc_hd__nor2_1_43/Y
+ sky130_fd_sc_hd__nor2_1_43/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_54 sky130_fd_sc_hd__nor2_1_57/B sky130_fd_sc_hd__nor2_1_54/Y
+ sky130_fd_sc_hd__nor2_1_54/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_65 sky130_fd_sc_hd__nor2_1_65/B sky130_fd_sc_hd__nor2_1_65/Y
+ sky130_fd_sc_hd__nor2_1_65/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_76 sky130_fd_sc_hd__nor2_1_76/B sky130_fd_sc_hd__nor2_1_76/Y
+ sky130_fd_sc_hd__nor2_2_10/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_87 sky130_fd_sc_hd__buf_6_1/X sky130_fd_sc_hd__nor2_1_87/Y
+ sky130_fd_sc_hd__nor2_1_87/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_98 sky130_fd_sc_hd__nor2_1_98/B sky130_fd_sc_hd__nor2_1_98/Y
+ sky130_fd_sc_hd__nor2_1_98/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_12_503 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_514 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_525 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_536 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_420 sky130_fd_sc_hd__nand2_1_420/Y sky130_fd_sc_hd__or2_1_0/A
+ sky130_fd_sc_hd__or2_1_0/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_547 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_431 sky130_fd_sc_hd__nand2_1_431/Y sky130_fd_sc_hd__nor2_1_142/A
+ sky130_fd_sc_hd__nor2_1_142/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_558 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_442 sky130_fd_sc_hd__nand2_1_442/Y sky130_fd_sc_hd__nor2_1_147/A
+ sky130_fd_sc_hd__nor2_1_147/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_569 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_453 sky130_fd_sc_hd__nand2_1_453/Y sky130_fd_sc_hd__buf_2_19/X
+ sky130_fd_sc_hd__buf_2_31/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_464 sky130_fd_sc_hd__nand2_1_464/Y sky130_fd_sc_hd__nand2_1_474/Y
+ sky130_fd_sc_hd__nand2_1_468/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_475 sky130_fd_sc_hd__xnor2_1_120/A sky130_fd_sc_hd__nand2_1_476/Y
+ sky130_fd_sc_hd__or2_0_50/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_486 sky130_fd_sc_hd__xnor2_1_67/A sky130_fd_sc_hd__nand2_1_487/Y
+ sky130_fd_sc_hd__or2_0_53/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_497 sky130_fd_sc_hd__nand2_1_497/Y sky130_fd_sc_hd__nor2_2_31/Y
+ sky130_fd_sc_hd__or2_0_72/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_11 sky130_fd_sc_hd__and3_4_15/C sky130_fd_sc_hd__nor2b_1_11/Y
+ sky130_fd_sc_hd__and3_4_15/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_22 sky130_fd_sc_hd__or2_0_84/A sky130_fd_sc_hd__fa_2_443/A
+ sky130_fd_sc_hd__xnor2_2_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_33 sky130_fd_sc_hd__mux2_2_9/X sky130_fd_sc_hd__nor2b_1_33/Y
+ sky130_fd_sc_hd__buf_2_214/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1000 sky130_fd_sc_hd__clkinv_1_1000/Y sky130_fd_sc_hd__clkinv_1_999/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_44 sky130_fd_sc_hd__or2_0_75/A sky130_fd_sc_hd__fa_2_473/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1011 sky130_fd_sc_hd__clkinv_1_1011/Y sky130_fd_sc_hd__clkinv_1_1011/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_55 sky130_fd_sc_hd__mux2_2_18/X sky130_fd_sc_hd__nor2b_1_55/Y
+ sky130_fd_sc_hd__buf_2_214/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1022 sky130_fd_sc_hd__buf_8_33/A sky130_fd_sc_hd__clkinv_1_1022/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_66 sky130_fd_sc_hd__mux2_2_46/X sky130_fd_sc_hd__fa_2_484/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1033 sky130_fd_sc_hd__clkinv_1_1034/A sky130_fd_sc_hd__buf_8_30/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_77 la_data_out[71] sky130_fd_sc_hd__nor2b_1_77/Y sky130_fd_sc_hd__mux2_4_5/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1044 sky130_fd_sc_hd__buf_8_20/A sky130_fd_sc_hd__clkinv_1_1044/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1502 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_88 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_88/Y
+ sky130_fd_sc_hd__nor2b_1_88/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1055 sky130_fd_sc_hd__inv_2_188/A sky130_fd_sc_hd__clkbuf_1_214/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1513 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_99 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_99/Y
+ sky130_fd_sc_hd__nor2b_1_99/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1066 sky130_fd_sc_hd__bufinv_8_2/A sky130_fd_sc_hd__buf_8_116/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_7 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_7/B sky130_fd_sc_hd__xnor2_1_7/Y
+ sky130_fd_sc_hd__xnor2_1_7/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_1524 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1077 sky130_fd_sc_hd__a22o_1_71/B2 la_data_out[48] vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1535 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1088 sky130_fd_sc_hd__o21ai_1_922/A2 sky130_fd_sc_hd__ha_2_58/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1546 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1099 sky130_fd_sc_hd__nor2b_1_125/B_N sky130_fd_sc_hd__nor4_1_1/D
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1557 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_260 sky130_fd_sc_hd__xor2_1_149/A sky130_fd_sc_hd__dfxtp_1_266/CLK
+ sky130_fd_sc_hd__and2_0_86/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1568 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_271 sky130_fd_sc_hd__xnor2_1_14/B sky130_fd_sc_hd__dfxtp_1_275/CLK
+ sky130_fd_sc_hd__and2_0_96/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1579 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_282 sky130_fd_sc_hd__dfxtp_1_282/Q sky130_fd_sc_hd__dfxtp_1_2/CLK
+ sky130_fd_sc_hd__and2_0_258/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_293 sky130_fd_sc_hd__dfxtp_1_293/Q sky130_fd_sc_hd__clkinv_8_6/Y
+ sky130_fd_sc_hd__and2_0_269/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__mux2_4_3 sky130_fd_sc_hd__or2_0_80/B sky130_fd_sc_hd__mux2_8_1/S
+ sky130_fd_sc_hd__buf_6_15/X sky130_fd_sc_hd__mux2_4_3/A1 vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__mux2_4
Xsky130_fd_sc_hd__o22ai_1_2 sky130_fd_sc_hd__o22ai_1_2/A2 sky130_fd_sc_hd__o22ai_1_2/B1
+ sky130_fd_sc_hd__o22ai_1_2/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__o22ai_1_9/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_110 sky130_fd_sc_hd__fa_2_104/CIN sky130_fd_sc_hd__fa_2_112/A
+ sky130_fd_sc_hd__fa_2_110/A sky130_fd_sc_hd__fa_2_110/B sky130_fd_sc_hd__xor2_1_148/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_121 sky130_fd_sc_hd__fa_2_119/B sky130_fd_sc_hd__fa_2_123/CIN
+ sky130_fd_sc_hd__fa_2_121/A sky130_fd_sc_hd__fa_2_121/B sky130_fd_sc_hd__xor2_1_165/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_132 sky130_fd_sc_hd__nor2_1_91/A sky130_fd_sc_hd__nor2_1_94/B
+ sky130_fd_sc_hd__fa_2_132/A sky130_fd_sc_hd__fa_2_132/B sky130_fd_sc_hd__fa_2_132/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_143 sky130_fd_sc_hd__xor3_1_11/C sky130_fd_sc_hd__fa_2_147/CIN
+ sky130_fd_sc_hd__fa_2_143/A sky130_fd_sc_hd__fa_2_143/B sky130_fd_sc_hd__fa_2_150/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_154 sky130_fd_sc_hd__fa_2_148/CIN sky130_fd_sc_hd__fa_2_151/B
+ sky130_fd_sc_hd__fa_2_154/A sky130_fd_sc_hd__fa_2_154/B sky130_fd_sc_hd__xor2_1_236/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_165 sky130_fd_sc_hd__fa_2_156/B sky130_fd_sc_hd__fa_2_166/B
+ sky130_fd_sc_hd__fa_2_165/A sky130_fd_sc_hd__fa_2_165/B sky130_fd_sc_hd__xor2_1_253/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and3_4_4 sky130_fd_sc_hd__and3_4_4/A sky130_fd_sc_hd__and3_4_4/B
+ sky130_fd_sc_hd__and3_4_4/C sky130_fd_sc_hd__and3_4_4/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__fa_2_176 sky130_fd_sc_hd__fa_2_160/A sky130_fd_sc_hd__fa_2_176/SUM
+ sky130_fd_sc_hd__fa_2_176/A sky130_fd_sc_hd__fa_2_176/B sky130_fd_sc_hd__fa_2_176/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_187 sky130_fd_sc_hd__fa_2_179/B sky130_fd_sc_hd__fa_2_191/A
+ sky130_fd_sc_hd__fa_2_187/A sky130_fd_sc_hd__fa_2_187/B sky130_fd_sc_hd__fa_2_187/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_198 sky130_fd_sc_hd__fa_2_187/CIN sky130_fd_sc_hd__fa_2_200/A
+ sky130_fd_sc_hd__fa_2_198/A sky130_fd_sc_hd__fa_2_198/B sky130_fd_sc_hd__xor2_1_290/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o22ai_1_20 sky130_fd_sc_hd__o22ai_1_43/B1 sky130_fd_sc_hd__o22ai_1_20/B1
+ sky130_fd_sc_hd__o22ai_1_20/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__inv_4_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_31 sky130_fd_sc_hd__o22ai_1_39/B1 sky130_fd_sc_hd__o21ai_1_9/A2
+ sky130_fd_sc_hd__o22ai_1_31/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__inv_4_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_42 sky130_fd_sc_hd__nor2_1_25/A sky130_fd_sc_hd__o22ai_1_42/B1
+ sky130_fd_sc_hd__o22ai_1_42/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_160 vccd1 vssd1 sky130_fd_sc_hd__buf_6_24/A sky130_fd_sc_hd__inv_2_126/Y
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_53 sky130_fd_sc_hd__nor2_1_14/A sky130_fd_sc_hd__o22ai_1_53/B1
+ sky130_fd_sc_hd__o22ai_1_53/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_171 vccd1 vssd1 la_data_out[51] sky130_fd_sc_hd__buf_8_75/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_64 sky130_fd_sc_hd__xnor2_2_6/Y sky130_fd_sc_hd__xnor2_1_223/Y
+ sky130_fd_sc_hd__o22ai_1_64/Y sky130_fd_sc_hd__xnor2_1_256/Y sky130_fd_sc_hd__o22ai_1_98/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_182 vccd1 vssd1 sky130_fd_sc_hd__buf_2_182/X sky130_fd_sc_hd__inv_2_197/Y
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_75 sky130_fd_sc_hd__nor2b_1_20/A sky130_fd_sc_hd__xnor2_1_225/Y
+ sky130_fd_sc_hd__ha_2_12/A sky130_fd_sc_hd__xnor2_1_226/Y sky130_fd_sc_hd__o22ai_1_78/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_193 vccd1 vssd1 sky130_fd_sc_hd__buf_2_193/X sky130_fd_sc_hd__buf_2_193/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_86 sky130_fd_sc_hd__xnor2_2_6/Y sky130_fd_sc_hd__o22ai_1_86/B1
+ sky130_fd_sc_hd__o22ai_1_86/Y sky130_fd_sc_hd__o22ai_1_86/A1 sky130_fd_sc_hd__o22ai_1_98/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_97 sky130_fd_sc_hd__xnor2_1_245/Y sky130_fd_sc_hd__xnor2_1_248/Y
+ sky130_fd_sc_hd__fa_2_445/B sky130_fd_sc_hd__inv_2_65/Y sky130_fd_sc_hd__o22ai_1_99/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_4_11 vccd1 vssd1 sky130_fd_sc_hd__buf_4_11/X sky130_fd_sc_hd__buf_4_11/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_22 vccd1 vssd1 sky130_fd_sc_hd__buf_4_22/X sky130_fd_sc_hd__buf_4_22/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_33 vccd1 vssd1 sky130_fd_sc_hd__buf_4_33/X sky130_fd_sc_hd__buf_8_17/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_12_104 sky130_fd_sc_hd__buf_8_30/X sky130_fd_sc_hd__buf_12_275/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_115 sky130_fd_sc_hd__buf_8_53/X sky130_fd_sc_hd__buf_12_115/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_126 sky130_fd_sc_hd__buf_8_60/X sky130_fd_sc_hd__buf_12_391/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_137 sky130_fd_sc_hd__buf_12_17/X sky130_fd_sc_hd__buf_12_137/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_60 vssd1 vccd1 sky130_fd_sc_hd__buf_8_25/A sky130_fd_sc_hd__clkbuf_1_60/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_148 sky130_fd_sc_hd__buf_12_20/X sky130_fd_sc_hd__buf_12_295/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_71 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_30/A1 sky130_fd_sc_hd__clkbuf_1_71/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_159 sky130_fd_sc_hd__buf_12_50/X sky130_fd_sc_hd__buf_12_307/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_82 vssd1 vccd1 sky130_fd_sc_hd__mux2_4_2/A1 sky130_fd_sc_hd__clkbuf_1_82/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_93 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_19/A1 sky130_fd_sc_hd__clkbuf_1_93/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_4_7 sky130_fd_sc_hd__clkbuf_4_7/X sky130_fd_sc_hd__clkbuf_4_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_1_304 sky130_fd_sc_hd__nand3_1_4/C sky130_fd_sc_hd__ha_2_4/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_315 sky130_fd_sc_hd__o21ai_1_186/A2 sky130_fd_sc_hd__xnor2_1_7/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_326 sky130_fd_sc_hd__nor2_1_51/B sky130_fd_sc_hd__nor2_1_54/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_337 sky130_fd_sc_hd__nor2_1_59/B sky130_fd_sc_hd__nand2_1_205/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_348 sky130_fd_sc_hd__a21oi_2_3/B1 sky130_fd_sc_hd__nand2_1_213/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_359 sky130_fd_sc_hd__nor2_1_67/B sky130_fd_sc_hd__nor2_1_70/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_201 la_data_out[54] sky130_fd_sc_hd__o21ai_1_923/Y sky130_fd_sc_hd__nor4b_1_0/D_N
+ sky130_fd_sc_hd__o21ai_1_923/A2 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__or2_0_40 sky130_fd_sc_hd__or2_0_60/A sky130_fd_sc_hd__or2_0_40/X
+ sky130_fd_sc_hd__or2_0_60/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_51 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__or2_0_51/X
+ sky130_fd_sc_hd__or2_0_51/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_62 sky130_fd_sc_hd__or2_0_62/A sky130_fd_sc_hd__or2_0_62/X
+ sky130_fd_sc_hd__or2_0_62/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_73 sky130_fd_sc_hd__or2_0_73/A sky130_fd_sc_hd__or2_0_73/X
+ sky130_fd_sc_hd__or2_0_73/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__clkinv_4_7 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkinv_4_7/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__or2_0_84 sky130_fd_sc_hd__or2_0_84/A sky130_fd_sc_hd__or2_0_84/X
+ sky130_fd_sc_hd__or2_0_84/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_95 sky130_fd_sc_hd__or2_0_95/A sky130_fd_sc_hd__or2_0_95/X
+ sky130_fd_sc_hd__or2_0_95/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__clkinv_4_120 sky130_fd_sc_hd__clkinv_8_76/Y sky130_fd_sc_hd__clkinv_8_77/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_12_660 sky130_fd_sc_hd__buf_12_660/A sky130_fd_sc_hd__buf_12_660/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_671 sky130_fd_sc_hd__buf_12_671/A sky130_fd_sc_hd__buf_12_671/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_300 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_682 sky130_fd_sc_hd__mux2_2_32/X la_data_out[72] vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_311 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_322 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_333 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_344 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_355 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_366 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_250 sky130_fd_sc_hd__nand2_1_250/Y sky130_fd_sc_hd__nand2_1_264/Y
+ sky130_fd_sc_hd__nand2_1_258/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_377 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_261 sky130_fd_sc_hd__nand2_1_261/Y sky130_fd_sc_hd__nand2_1_274/Y
+ sky130_fd_sc_hd__nand2_1_269/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_388 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_860 sky130_fd_sc_hd__clkinv_1_860/Y sky130_fd_sc_hd__inv_2_196/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_272 sky130_fd_sc_hd__nand2_1_272/Y sky130_fd_sc_hd__nand2_1_282/Y
+ sky130_fd_sc_hd__nand2_1_278/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_399 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_871 sky130_fd_sc_hd__clkinv_1_871/Y sky130_fd_sc_hd__clkinv_4_83/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_283 sky130_fd_sc_hd__nand2_1_283/Y sky130_fd_sc_hd__nand2_1_292/Y
+ sky130_fd_sc_hd__nand2_1_288/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_882 sky130_fd_sc_hd__clkinv_1_882/Y sky130_fd_sc_hd__clkinv_4_86/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_294 sky130_fd_sc_hd__xnor2_1_54/B sky130_fd_sc_hd__nand2_1_295/Y
+ sky130_fd_sc_hd__or2_0_16/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_893 sky130_fd_sc_hd__clkinv_1_893/Y sky130_fd_sc_hd__inv_2_102/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1310 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1321 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_60 sky130_fd_sc_hd__conb_1_60/LO sky130_fd_sc_hd__conb_1_60/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1332 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_71 sky130_fd_sc_hd__conb_1_71/LO sky130_fd_sc_hd__conb_1_71/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1343 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_82 sky130_fd_sc_hd__conb_1_82/LO sky130_fd_sc_hd__conb_1_82/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1354 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_93 sky130_fd_sc_hd__conb_1_93/LO sky130_fd_sc_hd__conb_1_93/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1365 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1376 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_807 vssd1 vccd1 sky130_fd_sc_hd__inv_2_43/Y sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_807/B1 sky130_fd_sc_hd__xor2_1_582/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1387 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_818 vssd1 vccd1 sky130_fd_sc_hd__inv_2_52/Y sky130_fd_sc_hd__nand2_1_609/Y
+ sky130_fd_sc_hd__a21oi_1_128/Y sky130_fd_sc_hd__xnor2_1_170/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1398 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_829 vssd1 vccd1 sky130_fd_sc_hd__buf_2_12/X sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_829/B1 sky130_fd_sc_hd__xor2_1_603/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__mux2_2_0 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_0/A1 sky130_fd_sc_hd__buf_6_22/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2b_2_8 sky130_fd_sc_hd__nor2_4_18/B sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__nor2_4_18/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_2
Xsky130_fd_sc_hd__xor2_1_601 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__fah_1_10/A
+ sky130_fd_sc_hd__xor2_1_601/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_612 sky130_fd_sc_hd__xor2_1_612/B sky130_fd_sc_hd__xor2_1_612/X
+ sky130_fd_sc_hd__xor2_1_612/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_623 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__or2_0_62/A
+ sky130_fd_sc_hd__xor2_1_623/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_634 sky130_fd_sc_hd__o21a_1_5/A1 sky130_fd_sc_hd__xor2_1_634/X
+ sky130_fd_sc_hd__xor2_1_634/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_645 sky130_fd_sc_hd__xor2_1_645/B sky130_fd_sc_hd__xor2_1_645/X
+ sky130_fd_sc_hd__xor2_1_645/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_656 sky130_fd_sc_hd__xor2_1_656/B sky130_fd_sc_hd__xor2_1_656/X
+ sky130_fd_sc_hd__xor2_1_656/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_667 sky130_fd_sc_hd__xnor2_2_4/A sky130_fd_sc_hd__xor2_1_667/X
+ sky130_fd_sc_hd__xnor2_2_5/B vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_678 sky130_fd_sc_hd__xor2_1_678/B sky130_fd_sc_hd__xor2_1_678/X
+ sky130_fd_sc_hd__xor2_1_678/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_689 sky130_fd_sc_hd__buf_2_175/A sky130_fd_sc_hd__xor2_1_689/X
+ sky130_fd_sc_hd__xor2_1_689/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__fa_2_8 sky130_fd_sc_hd__xor3_1_6/B sky130_fd_sc_hd__fa_2_8/SUM sky130_fd_sc_hd__fa_2_8/A
+ sky130_fd_sc_hd__fa_2_8/B sky130_fd_sc_hd__fa_2_8/CIN vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a211o_1_14 vssd1 vccd1 sky130_fd_sc_hd__fa_2_253/A sky130_fd_sc_hd__dfxtp_1_77/Q
+ sky130_fd_sc_hd__nor2_1_18/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_14/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__a211o_1_25 vssd1 vccd1 sky130_fd_sc_hd__fa_2_187/A sky130_fd_sc_hd__dfxtp_1_88/Q
+ sky130_fd_sc_hd__nor2_1_29/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_25/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__clkinv_1_101 io_out[0] sky130_fd_sc_hd__conb_1_41/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_112 io_oeb[27] sky130_fd_sc_hd__conb_1_30/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_123 io_oeb[16] sky130_fd_sc_hd__conb_1_19/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_134 io_oeb[5] sky130_fd_sc_hd__conb_1_8/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_145 sky130_fd_sc_hd__clkinv_4_33/A sky130_fd_sc_hd__buf_2_203/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_156 sky130_fd_sc_hd__o21ai_1_3/A2 sky130_fd_sc_hd__dfxtp_1_123/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_167 sky130_fd_sc_hd__nor2_1_29/A sky130_fd_sc_hd__dfxtp_1_152/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_178 sky130_fd_sc_hd__o22ai_1_41/B1 sky130_fd_sc_hd__dfxtp_1_181/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_14 sky130_fd_sc_hd__inv_2_66/Y sky130_fd_sc_hd__or2_0_89/B
+ sky130_fd_sc_hd__a22o_1_14/X sky130_fd_sc_hd__nor2_1_233/Y sky130_fd_sc_hd__a22o_1_14/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_189 sky130_fd_sc_hd__o22ai_1_19/B1 sky130_fd_sc_hd__dfxtp_1_114/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_25 sky130_fd_sc_hd__buf_2_63/A sky130_fd_sc_hd__buf_2_100/X
+ sky130_fd_sc_hd__a22o_1_25/X sky130_fd_sc_hd__a22o_1_25/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_36 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__buf_2_111/X
+ sky130_fd_sc_hd__a22o_1_36/X sky130_fd_sc_hd__a22o_1_36/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_47 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__buf_2_122/X
+ sky130_fd_sc_hd__a22o_1_47/X sky130_fd_sc_hd__a22o_1_47/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__o21ai_1_1 vssd1 vccd1 sky130_fd_sc_hd__o21ai_2_1/A2 sky130_fd_sc_hd__a21oi_1_0/Y
+ sky130_fd_sc_hd__buf_2_16/A sky130_fd_sc_hd__o21ai_1_1/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a22o_1_58 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__buf_2_48/A
+ sky130_fd_sc_hd__a22o_1_58/X sky130_fd_sc_hd__ha_2_29/SUM sky130_fd_sc_hd__a22o_1_71/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_69 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__buf_2_43/A
+ sky130_fd_sc_hd__a22o_1_69/X sky130_fd_sc_hd__ha_2_38/SUM sky130_fd_sc_hd__a22o_1_71/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__bufbuf_16_0 sky130_fd_sc_hd__clkbuf_1_35/X sky130_fd_sc_hd__buf_6_59/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__bufbuf_16
Xsky130_fd_sc_hd__edfxbp_1_0 vccd1 vssd1 sky130_fd_sc_hd__edfxbp_1_0/CLK sky130_fd_sc_hd__nor2_1_273/A
+ sky130_fd_sc_hd__o21ai_1_910/Y sky130_fd_sc_hd__edfxbp_1_0/D sky130_fd_sc_hd__edfxbp_1_0/Q
+ vssd1 vccd1 sky130_fd_sc_hd__edfxbp_1
Xsky130_fd_sc_hd__nor2_1_250 sky130_fd_sc_hd__nor2_1_251/Y sky130_fd_sc_hd__nor2_1_250/Y
+ sky130_fd_sc_hd__nor2_1_252/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_2_4 sky130_fd_sc_hd__clkinv_2_5/A sky130_fd_sc_hd__clkinv_8_3/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__nor2_1_261 sky130_fd_sc_hd__nor2_1_261/B sky130_fd_sc_hd__nor2_1_261/Y
+ sky130_fd_sc_hd__nor2_1_261/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_272 sky130_fd_sc_hd__nor2_1_278/B sky130_fd_sc_hd__nand3_1_5/B
+ sky130_fd_sc_hd__nor2_2_0/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_283 sky130_fd_sc_hd__a21o_2_3/A2 sky130_fd_sc_hd__a21o_2_3/B1
+ wbs_adr_i[7] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_490 sky130_fd_sc_hd__buf_12_490/A sky130_fd_sc_hd__buf_12_582/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_130 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_141 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_152 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_163 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_174 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_185 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_15 sky130_fd_sc_hd__nand2_1_15/Y sky130_fd_sc_hd__nand2_1_15/B
+ sky130_fd_sc_hd__nand2_1_15/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_220 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_5/B sky130_fd_sc_hd__xnor2_1_220/Y
+ la_data_out[72] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_196 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_26 sky130_fd_sc_hd__buf_6_1/A sky130_fd_sc_hd__nand2_1_27/Y
+ sky130_fd_sc_hd__nand2_1_28/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_231 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_4/B sky130_fd_sc_hd__xnor2_1_231/Y
+ la_data_out[72] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_37 sky130_fd_sc_hd__buf_4_7/A sky130_fd_sc_hd__nand2_1_38/Y
+ sky130_fd_sc_hd__nand2_1_39/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_242 vssd1 vccd1 sky130_fd_sc_hd__or2_1_10/A sky130_fd_sc_hd__xnor2_1_242/Y
+ sky130_fd_sc_hd__or2_0_84/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_48 sky130_fd_sc_hd__nor2_2_1/A sky130_fd_sc_hd__nor2_4_0/B
+ sky130_fd_sc_hd__nor2_2_0/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_690 sky130_fd_sc_hd__xor2_1_664/A sky130_fd_sc_hd__o21ai_1_889/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_253 vssd1 vccd1 la_data_out[77] sky130_fd_sc_hd__xnor2_1_253/Y
+ sky130_fd_sc_hd__mux2_2_31/X vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_59 sky130_fd_sc_hd__nand2_1_59/Y sky130_fd_sc_hd__nand2_1_59/B
+ sky130_fd_sc_hd__nor2_4_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_264 vssd1 vccd1 la_data_out[68] sky130_fd_sc_hd__xnor2_1_264/Y
+ sky130_fd_sc_hd__or2_0_79/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_275 vssd1 vccd1 la_data_out[81] sky130_fd_sc_hd__xnor2_1_275/Y
+ sky130_fd_sc_hd__mux2_2_31/X vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_286 vssd1 vccd1 sky130_fd_sc_hd__or2_0_82/B sky130_fd_sc_hd__xnor2_1_286/Y
+ sky130_fd_sc_hd__or2_0_78/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_297 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_297/B sky130_fd_sc_hd__xnor2_1_297/Y
+ sky130_fd_sc_hd__xnor2_1_297/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_1140 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1151 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1162 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1173 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_604 vssd1 vccd1 sky130_fd_sc_hd__inv_2_27/Y sky130_fd_sc_hd__nand2b_2_3/Y
+ sky130_fd_sc_hd__nand2_1_329/Y sky130_fd_sc_hd__xor2_1_395/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1184 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_615 vssd1 vccd1 sky130_fd_sc_hd__buf_2_10/X sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_615/B1 sky130_fd_sc_hd__xor2_1_407/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1195 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_626 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_162/Y sky130_fd_sc_hd__o21a_1_3/X
+ sky130_fd_sc_hd__nand2_1_485/Y sky130_fd_sc_hd__xnor2_1_123/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_637 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_3/Y sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__o21ai_1_637/B1 sky130_fd_sc_hd__xor2_1_579/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_648 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_771/A2 sky130_fd_sc_hd__nand2b_1_16/Y
+ sky130_fd_sc_hd__o21ai_1_648/B1 sky130_fd_sc_hd__xor2_1_435/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_659 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_10/X sky130_fd_sc_hd__nand2_1_513/Y
+ sky130_fd_sc_hd__a21oi_1_108/Y sky130_fd_sc_hd__xnor2_1_133/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fah_1_2 sky130_fd_sc_hd__or2_0_37/A sky130_fd_sc_hd__fah_1_2/B sky130_fd_sc_hd__fah_1_2/A
+ sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__fah_1_2/CI vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__fah_1
Xsky130_fd_sc_hd__xor2_1_420 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__xor2_1_420/X
+ sky130_fd_sc_hd__xor2_1_420/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_90 vssd1 vccd1 sky130_fd_sc_hd__fa_2_239/A sky130_fd_sc_hd__and3_4_14/C
+ sky130_fd_sc_hd__xnor2_1_90/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_431 sky130_fd_sc_hd__fa_2_357/A sky130_fd_sc_hd__xor3_1_28/C
+ sky130_fd_sc_hd__xor2_1_431/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_442 sky130_fd_sc_hd__fah_1_14/A sky130_fd_sc_hd__fa_2_284/B
+ sky130_fd_sc_hd__xor2_1_442/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_453 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__xor2_1_453/X
+ sky130_fd_sc_hd__xor2_1_453/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_464 sky130_fd_sc_hd__fa_2_310/A sky130_fd_sc_hd__fa_2_301/B
+ sky130_fd_sc_hd__xor2_1_464/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_475 sky130_fd_sc_hd__fa_2_310/A sky130_fd_sc_hd__and3_1_2/B
+ sky130_fd_sc_hd__xor2_1_475/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_486 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__fa_2_322/A
+ sky130_fd_sc_hd__xor2_1_486/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_497 sky130_fd_sc_hd__xor2_1_548/B sky130_fd_sc_hd__xor2_1_497/X
+ sky130_fd_sc_hd__xor2_1_497/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a222oi_1_506 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__nor2_2_10/B sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__buf_6_4/X
+ sky130_fd_sc_hd__o21ai_1_803/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_517 vccd1 vssd1 sky130_fd_sc_hd__and3_4_20/X sky130_fd_sc_hd__or2_0_71/B
+ sky130_fd_sc_hd__buf_2_29/X sky130_fd_sc_hd__nor2_4_16/Y sky130_fd_sc_hd__buf_2_30/X
+ sky130_fd_sc_hd__o21ai_1_814/B1 sky130_fd_sc_hd__and2b_4_11/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_528 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__buf_2_31/X
+ sky130_fd_sc_hd__buf_2_4/A sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__buf_2_20/X
+ sky130_fd_sc_hd__o21ai_1_832/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_539 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__or2_0_52/B
+ sky130_fd_sc_hd__buf_2_25/A sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__o21ai_1_851/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nor2b_1_106 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_106/Y
+ sky130_fd_sc_hd__nor2b_1_106/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_117 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_117/Y
+ sky130_fd_sc_hd__nor2b_1_117/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_128 sky130_fd_sc_hd__clkinv_4_47/Y sky130_fd_sc_hd__nor2b_1_128/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_139 sky130_fd_sc_hd__clkinv_4_58/Y sky130_fd_sc_hd__nor2b_1_139/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__buf_6_7 vccd1 vssd1 sky130_fd_sc_hd__buf_6_7/X sky130_fd_sc_hd__buf_6_7/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__clkinv_2_20 sky130_fd_sc_hd__inv_2_112/A sky130_fd_sc_hd__inv_4_10/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_31 sky130_fd_sc_hd__clkinv_2_32/A sky130_fd_sc_hd__nand2_1_845/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_42 sky130_fd_sc_hd__inv_2_168/A sky130_fd_sc_hd__buf_8_99/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__and2_0_400 vccd1 vssd1 sky130_fd_sc_hd__and2_0_400/X sky130_fd_sc_hd__and2_0_401/B
+ sky130_fd_sc_hd__and2_0_400/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_2_53 la_data_out[94] sky130_fd_sc_hd__inv_2_153/A vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__inv_2_200 sky130_fd_sc_hd__inv_2_200/A sky130_fd_sc_hd__buf_6_6/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__or2_1_2 sky130_fd_sc_hd__or2_1_2/A sky130_fd_sc_hd__or2_1_2/X sky130_fd_sc_hd__or2_1_2/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_1
Xsky130_fd_sc_hd__sdlclkp_4_5 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_4_1/Y
+ sky130_fd_sc_hd__dfxtp_1_81/CLK sky130_fd_sc_hd__o21ai_2_0/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_8 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_8/Y
+ sky130_fd_sc_hd__nor2_1_8/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_190 sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__xnor2_1_125/Y sky130_fd_sc_hd__xnor2_1_62/Y sky130_fd_sc_hd__a22oi_1_190/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__o21ai_1_401 vssd1 vccd1 sky130_fd_sc_hd__a21oi_1_100/Y sky130_fd_sc_hd__nand2_1_455/Y
+ sky130_fd_sc_hd__a21oi_1_95/Y sky130_fd_sc_hd__inv_2_42/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_412 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_412/A2 sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_412/B1 sky130_fd_sc_hd__xor2_1_223/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_423 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_444/A2 sky130_fd_sc_hd__nor2_1_108/A
+ sky130_fd_sc_hd__a21oi_1_74/Y sky130_fd_sc_hd__o21ai_1_423/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_434 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_434/A2 sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_434/B1 sky130_fd_sc_hd__xor2_1_241/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_445 vssd1 vccd1 sky130_fd_sc_hd__inv_2_39/Y sky130_fd_sc_hd__nand2b_2_3/Y
+ sky130_fd_sc_hd__o21ai_1_445/B1 sky130_fd_sc_hd__xor2_1_248/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_456 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_119/Y sky130_fd_sc_hd__nor2_1_115/A
+ sky130_fd_sc_hd__nor2_1_114/Y sky130_fd_sc_hd__o21ai_1_456/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_467 vssd1 vccd1 sky130_fd_sc_hd__inv_2_30/Y sky130_fd_sc_hd__nand2b_1_8/Y
+ sky130_fd_sc_hd__o21ai_1_467/B1 sky130_fd_sc_hd__xor2_1_270/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_478 vssd1 vccd1 sky130_fd_sc_hd__inv_2_39/Y sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_478/B1 sky130_fd_sc_hd__xor2_1_279/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_489 vssd1 vccd1 sky130_fd_sc_hd__buf_2_10/X sky130_fd_sc_hd__nand2b_1_13/Y
+ sky130_fd_sc_hd__o21ai_1_489/B1 sky130_fd_sc_hd__xor2_1_289/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2_4_10 sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__and3_4_3/B
+ sky130_fd_sc_hd__and3_4_3/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__nand2_1_805 sky130_fd_sc_hd__nand2_1_805/Y sky130_fd_sc_hd__nor2_1_257/A
+ sky130_fd_sc_hd__nor2_1_257/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_816 sky130_fd_sc_hd__xor2_1_682/B sky130_fd_sc_hd__nand2_1_817/Y
+ sky130_fd_sc_hd__nand2_1_816/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_827 sky130_fd_sc_hd__nand2_1_827/Y sky130_fd_sc_hd__or2_0_108/A
+ sky130_fd_sc_hd__or2_0_108/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_838 sky130_fd_sc_hd__xnor2_1_302/B sky130_fd_sc_hd__nand2_1_839/Y
+ sky130_fd_sc_hd__or2_0_111/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_849 sky130_fd_sc_hd__nand2_1_849/Y sky130_fd_sc_hd__nor2_2_1/B
+ sky130_fd_sc_hd__a22o_1_71/B1 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o21ai_1_16 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_17/B1 sky130_fd_sc_hd__inv_2_53/A
+ sky130_fd_sc_hd__o21ai_1_16/B1 sky130_fd_sc_hd__fa_2_102/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_27 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_6/B1 sky130_fd_sc_hd__nor2_4_4/B
+ sky130_fd_sc_hd__o21ai_1_27/B1 sky130_fd_sc_hd__fa_2_137/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_250 sky130_fd_sc_hd__fa_2_198/A sky130_fd_sc_hd__fa_2_164/B
+ sky130_fd_sc_hd__xor2_1_250/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__o21ai_1_38 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_41/A2 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_86/Y sky130_fd_sc_hd__and2_0_13/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_261 sky130_fd_sc_hd__fa_2_170/A sky130_fd_sc_hd__xor2_1_261/X
+ sky130_fd_sc_hd__xor2_1_261/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__o21ai_1_49 vssd1 vccd1 sky130_fd_sc_hd__inv_2_63/Y sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__o21ai_1_49/B1 sky130_fd_sc_hd__o21ai_1_49/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_272 sky130_fd_sc_hd__fa_2_217/A sky130_fd_sc_hd__fa_2_181/A
+ sky130_fd_sc_hd__xor2_1_272/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_283 sky130_fd_sc_hd__xor2_1_383/B sky130_fd_sc_hd__fa_2_190/A
+ sky130_fd_sc_hd__xor2_1_283/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_294 sky130_fd_sc_hd__fa_2_239/A sky130_fd_sc_hd__fa_2_195/B
+ sky130_fd_sc_hd__xor2_1_294/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_210 vssd1 vccd1 sky130_fd_sc_hd__buf_8_22/A sky130_fd_sc_hd__inv_2_81/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_221 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2_33/A sky130_fd_sc_hd__nand2_2_6/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_232 vssd1 vccd1 sky130_fd_sc_hd__buf_8_130/A sky130_fd_sc_hd__buf_6_17/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_303 vccd1 vssd1 sky130_fd_sc_hd__and3_4_15/X sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__inv_6_0/Y sky130_fd_sc_hd__nor2_1_130/Y sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__o21ai_1_517/B1 sky130_fd_sc_hd__nor2b_1_11/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_243 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_16_0/A sky130_fd_sc_hd__clkbuf_4_27/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_314 vccd1 vssd1 sky130_fd_sc_hd__and3_4_16/X sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__buf_6_2/X sky130_fd_sc_hd__nor2_2_19/Y sky130_fd_sc_hd__buf_4_7/X
+ sky130_fd_sc_hd__o21ai_1_529/B1 sky130_fd_sc_hd__nor2b_2_3/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_254 vssd1 vccd1 sky130_fd_sc_hd__buf_8_123/A sky130_fd_sc_hd__clkbuf_1_254/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_2_1 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__dfxtp_2_1/CLK
+ sky130_fd_sc_hd__dfxtp_2_1/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_2
Xsky130_fd_sc_hd__a222oi_1_325 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__nor2_1_73/B sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__o21ai_1_543/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_265 vssd1 vccd1 sky130_fd_sc_hd__buf_8_10/A sky130_fd_sc_hd__clkbuf_1_326/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_336 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__and2_0_38/A sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__and2_0_49/A
+ sky130_fd_sc_hd__o21ai_1_558/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_276 vssd1 vccd1 sky130_fd_sc_hd__buf_8_142/A sky130_fd_sc_hd__clkbuf_1_55/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_347 vccd1 vssd1 sky130_fd_sc_hd__and3_4_17/X sky130_fd_sc_hd__or2_0_52/B
+ sky130_fd_sc_hd__or2_0_53/A sky130_fd_sc_hd__nor2_2_20/Y sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__o21ai_1_574/B1 sky130_fd_sc_hd__nor2b_2_4/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_287 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_288/A sky130_fd_sc_hd__buf_8_28/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_358 vccd1 vssd1 sky130_fd_sc_hd__and3_4_10/X sky130_fd_sc_hd__or2_0_52/B
+ sky130_fd_sc_hd__or2_0_53/A sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__o21ai_1_592/B1 sky130_fd_sc_hd__and2b_4_7/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_298 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_299/A sky130_fd_sc_hd__buf_8_63/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_369 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__buf_6_2/X sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__buf_4_7/X
+ sky130_fd_sc_hd__o21ai_1_611/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__buf_4_4 vccd1 vssd1 sky130_fd_sc_hd__buf_4_4/X sky130_fd_sc_hd__buf_4_4/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__and2_0_230 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_88/D sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__o21ai_1_58/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_241 vccd1 vssd1 sky130_fd_sc_hd__and2_0_241/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_241/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_252 vccd1 vssd1 sky130_fd_sc_hd__and2_0_252/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__and2_0_284/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_263 vccd1 vssd1 sky130_fd_sc_hd__and2_0_263/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__and2_0_263/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_274 vccd1 vssd1 sky130_fd_sc_hd__and2_0_274/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__xor2_1_641/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__a21oi_2_15 sky130_fd_sc_hd__a21oi_2_15/B1 sky130_fd_sc_hd__or2_1_7/X
+ sky130_fd_sc_hd__o21ai_2_13/Y sky130_fd_sc_hd__xor2_1_468/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_2
Xsky130_fd_sc_hd__and2_0_285 vccd1 vssd1 sky130_fd_sc_hd__and2_0_285/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_6/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_296 vccd1 vssd1 sky130_fd_sc_hd__and2_0_296/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_17/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__sdlclkp_2_2 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_8_1/Y
+ sky130_fd_sc_hd__dfxtp_1_78/CLK sky130_fd_sc_hd__o21ai_2_0/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__inv_4_4 sky130_fd_sc_hd__inv_4_4/Y sky130_fd_sc_hd__inv_4_4/A vccd1
+ vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__or2_0_109 sky130_fd_sc_hd__or2_0_109/A sky130_fd_sc_hd__or2_0_109/X
+ sky130_fd_sc_hd__or2_0_109/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__o21ai_1_220 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_2/X sky130_fd_sc_hd__nand2_1_186/Y
+ sky130_fd_sc_hd__a21oi_1_42/Y sky130_fd_sc_hd__xnor2_1_13/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_231 vssd1 vccd1 sky130_fd_sc_hd__inv_2_13/Y sky130_fd_sc_hd__nand2b_1_1/Y
+ sky130_fd_sc_hd__a222oi_1_99/Y sky130_fd_sc_hd__xor2_1_56/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_242 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_2/X sky130_fd_sc_hd__nand2_1_197/Y
+ sky130_fd_sc_hd__a21oi_1_44/Y sky130_fd_sc_hd__xnor2_1_17/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_253 vssd1 vccd1 sky130_fd_sc_hd__inv_2_24/Y sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__o21ai_1_253/B1 sky130_fd_sc_hd__xor2_1_75/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_264 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_0/Y sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__o21ai_1_264/B1 sky130_fd_sc_hd__xor2_1_86/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_275 vssd1 vccd1 sky130_fd_sc_hd__inv_2_12/Y sky130_fd_sc_hd__nand2b_2_0/Y
+ sky130_fd_sc_hd__o21ai_1_275/B1 sky130_fd_sc_hd__xor2_1_96/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_286 vssd1 vccd1 sky130_fd_sc_hd__buf_2_1/X sky130_fd_sc_hd__nand2b_1_7/Y
+ sky130_fd_sc_hd__o21ai_1_286/B1 sky130_fd_sc_hd__xor2_1_107/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_297 vssd1 vccd1 sky130_fd_sc_hd__inv_2_22/Y sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__o21ai_1_297/B1 sky130_fd_sc_hd__xor2_1_118/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_707 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_718 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_602 sky130_fd_sc_hd__xnor2_1_166/A sky130_fd_sc_hd__nand2_1_602/B
+ sky130_fd_sc_hd__nand2_1_602/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_729 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_613 sky130_fd_sc_hd__nand2_1_613/Y sky130_fd_sc_hd__nor2_1_200/A
+ sky130_fd_sc_hd__nor2_1_200/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_624 sky130_fd_sc_hd__nand2_1_624/Y sky130_fd_sc_hd__buf_2_4/A
+ sky130_fd_sc_hd__buf_2_15/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_635 sky130_fd_sc_hd__nand2_1_635/Y sky130_fd_sc_hd__nand2_1_645/Y
+ sky130_fd_sc_hd__nand2_1_639/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_646 sky130_fd_sc_hd__xnor2_1_182/A sky130_fd_sc_hd__nand2_1_647/Y
+ sky130_fd_sc_hd__or2_0_68/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_657 sky130_fd_sc_hd__nand2_1_657/Y sky130_fd_sc_hd__or2_0_72/A
+ sky130_fd_sc_hd__or2_0_71/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_668 sky130_fd_sc_hd__xor2_1_641/B sky130_fd_sc_hd__nand2_1_669/Y
+ sky130_fd_sc_hd__nand2_1_668/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_2_4 sky130_fd_sc_hd__nor2_2_20/A sky130_fd_sc_hd__nor2b_2_4/A
+ sky130_fd_sc_hd__nor2b_2_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_2
Xsky130_fd_sc_hd__nand2_1_679 sky130_fd_sc_hd__nand2_1_679/Y sky130_fd_sc_hd__or2_1_11/A
+ sky130_fd_sc_hd__or2_1_11/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_1706 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1717 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_16 sky130_fd_sc_hd__inv_2_16/A sky130_fd_sc_hd__inv_2_16/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_420 sky130_fd_sc_hd__dfxtp_1_420/Q sky130_fd_sc_hd__dfxtp_1_427/CLK
+ sky130_fd_sc_hd__nor2b_1_95/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1728 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_27 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__inv_2_27/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_431 sky130_fd_sc_hd__dfxtp_1_431/Q sky130_fd_sc_hd__clkinv_4_9/Y
+ sky130_fd_sc_hd__nor2b_1_116/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1739 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_38 sky130_fd_sc_hd__inv_2_38/A sky130_fd_sc_hd__inv_2_38/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_442 sky130_fd_sc_hd__dfxtp_1_442/Q sky130_fd_sc_hd__dfxtp_1_446/CLK
+ sky130_fd_sc_hd__nor2b_1_105/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_49 sky130_fd_sc_hd__inv_2_49/A sky130_fd_sc_hd__inv_2_49/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_453 sky130_fd_sc_hd__dfxtp_1_453/Q sky130_fd_sc_hd__dfxtp_1_459/CLK
+ sky130_fd_sc_hd__nor2b_1_94/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_464 sky130_fd_sc_hd__ha_2_48/A sky130_fd_sc_hd__dfxtp_1_515/CLK
+ sky130_fd_sc_hd__and2_0_354/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_475 sky130_fd_sc_hd__ha_2_23/A sky130_fd_sc_hd__dfxtp_1_480/CLK
+ sky130_fd_sc_hd__and2_0_386/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_486 sky130_fd_sc_hd__ha_2_35/A sky130_fd_sc_hd__dfxtp_1_489/CLK
+ sky130_fd_sc_hd__and2_0_374/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_2_6 sky130_fd_sc_hd__nand2_2_6/Y sky130_fd_sc_hd__nand2_2_6/A
+ sky130_fd_sc_hd__nand2_2_6/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__dfxtp_1_497 la_data_out[46] sky130_fd_sc_hd__dfxtp_1_498/CLK sky130_fd_sc_hd__and2_0_373/X
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a222oi_1_100 vccd1 vssd1 sky130_fd_sc_hd__and3_4_7/X sky130_fd_sc_hd__buf_2_4/X
+ sky130_fd_sc_hd__buf_6_5/X sky130_fd_sc_hd__nor2_2_7/Y sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__o21ai_1_232/B1 sky130_fd_sc_hd__nor2b_2_1/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2b_1_12 sky130_fd_sc_hd__nand2b_1_12/Y sky130_fd_sc_hd__and3_4_13/C
+ sky130_fd_sc_hd__and3_4_13/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a222oi_1_111 vccd1 vssd1 sky130_fd_sc_hd__and3_4_8/X sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__nor2_1_87/A sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__o21ai_1_247/B1 sky130_fd_sc_hd__nor2b_2_2/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2b_1_23 sky130_fd_sc_hd__o22ai_1_86/A1 sky130_fd_sc_hd__or2_0_84/A
+ la_data_out[79] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a222oi_1_122 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__buf_4_2/X sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__o21ai_1_260/B1 sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2b_1_34 sky130_fd_sc_hd__nand2b_1_34/Y sky130_fd_sc_hd__ha_2_57/SUM
+ la_data_out[53] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a222oi_1_133 vccd1 vssd1 sky130_fd_sc_hd__and3_4_1/X sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__nor2_1_87/A sky130_fd_sc_hd__nor2_2_9/Y sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__o21ai_1_275/B1 sky130_fd_sc_hd__and2b_4_3/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_144 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__buf_6_4/X
+ sky130_fd_sc_hd__buf_6_0/X sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__o21ai_1_289/B1 sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_155 vccd1 vssd1 sky130_fd_sc_hd__and3_4_7/X sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__buf_8_0/X sky130_fd_sc_hd__nor2_2_7/Y sky130_fd_sc_hd__buf_4_6/X
+ sky130_fd_sc_hd__o21ai_1_302/B1 sky130_fd_sc_hd__nor2b_2_1/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_303 sky130_fd_sc_hd__fa_2_298/A sky130_fd_sc_hd__fa_2_308/A
+ sky130_fd_sc_hd__fa_2_303/A sky130_fd_sc_hd__fa_2_303/B sky130_fd_sc_hd__xor2_1_461/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_166 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__nor2_1_85/B sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__nor2_2_10/B
+ sky130_fd_sc_hd__o21ai_1_317/B1 sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_314 sky130_fd_sc_hd__fa_2_307/A sky130_fd_sc_hd__fa_2_315/B
+ sky130_fd_sc_hd__fa_2_314/A sky130_fd_sc_hd__fa_2_314/B sky130_fd_sc_hd__fa_2_314/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_177 vccd1 vssd1 sky130_fd_sc_hd__and3_4_1/X sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__and2_0_25/A sky130_fd_sc_hd__nor2_2_9/Y sky130_fd_sc_hd__nor2_2_5/A
+ sky130_fd_sc_hd__o21ai_1_333/B1 sky130_fd_sc_hd__and2b_4_3/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_325 sky130_fd_sc_hd__nor2_2_21/A sky130_fd_sc_hd__or2_1_7/B
+ sky130_fd_sc_hd__fa_2_325/A sky130_fd_sc_hd__fa_2_325/B sky130_fd_sc_hd__fa_2_325/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_188 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__buf_6_1/X sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__o21ai_1_349/B1 sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_336 sky130_fd_sc_hd__fa_2_329/A sky130_fd_sc_hd__fa_2_337/B
+ sky130_fd_sc_hd__fa_2_336/A sky130_fd_sc_hd__fa_2_336/B sky130_fd_sc_hd__fa_2_336/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_199 vccd1 vssd1 sky130_fd_sc_hd__and3_4_2/X sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__buf_2_32/X sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__o21ai_1_368/B1 sky130_fd_sc_hd__and2b_4_4/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_347 sky130_fd_sc_hd__fa_2_334/B sky130_fd_sc_hd__fa_2_342/B
+ sky130_fd_sc_hd__fa_2_347/A sky130_fd_sc_hd__fa_2_347/B sky130_fd_sc_hd__xor2_1_512/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_358 sky130_fd_sc_hd__fa_2_352/A sky130_fd_sc_hd__fa_2_359/B
+ sky130_fd_sc_hd__fa_2_358/A sky130_fd_sc_hd__fa_2_358/B sky130_fd_sc_hd__xor2_1_527/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_369 sky130_fd_sc_hd__fa_2_366/CIN sky130_fd_sc_hd__fa_2_374/A
+ sky130_fd_sc_hd__fa_2_369/A sky130_fd_sc_hd__fa_2_369/B sky130_fd_sc_hd__xor2_1_546/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_8_30 sky130_fd_sc_hd__clkinv_8_30/Y sky130_fd_sc_hd__clkinv_8_30/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_41 sky130_fd_sc_hd__clkinv_8_42/A sky130_fd_sc_hd__clkinv_8_41/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_52 sky130_fd_sc_hd__clkinv_8_53/A sky130_fd_sc_hd__clkinv_8_69/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_63 sky130_fd_sc_hd__clkinv_8_4/A sky130_fd_sc_hd__clkinv_8_63/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_74 sky130_fd_sc_hd__dfxtp_1_0/CLK sky130_fd_sc_hd__clkinv_8_74/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_85 sky130_fd_sc_hd__clkinv_8_86/A sky130_fd_sc_hd__clkinv_8_85/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_50 sky130_fd_sc_hd__buf_12_50/A sky130_fd_sc_hd__buf_12_50/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_61 sky130_fd_sc_hd__buf_12_61/A sky130_fd_sc_hd__buf_12_61/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_72 sky130_fd_sc_hd__buf_4_29/X sky130_fd_sc_hd__buf_12_72/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_83 sky130_fd_sc_hd__buf_12_83/A sky130_fd_sc_hd__buf_12_83/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_94 sky130_fd_sc_hd__buf_8_27/X sky130_fd_sc_hd__buf_12_94/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_2_1 vccd1 vssd1 sky130_fd_sc_hd__buf_2_1/X sky130_fd_sc_hd__buf_2_1/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_12_308 sky130_fd_sc_hd__buf_12_86/X sky130_fd_sc_hd__buf_12_493/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_319 sky130_fd_sc_hd__buf_12_70/X sky130_fd_sc_hd__buf_12_666/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__inv_2_1 sky130_fd_sc_hd__inv_2_1/A sky130_fd_sc_hd__inv_2_1/Y vccd1
+ vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__clkinv_1_508 sky130_fd_sc_hd__clkinv_1_508/Y sky130_fd_sc_hd__nand2_1_491/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_519 sky130_fd_sc_hd__o21ai_1_649/A2 sky130_fd_sc_hd__xnor2_1_131/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_11 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_11/Y
+ sky130_fd_sc_hd__nor2_1_11/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_22 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_22/Y
+ sky130_fd_sc_hd__nor2_1_22/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_33 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_33/Y
+ sky130_fd_sc_hd__nor2_1_33/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_44 sky130_fd_sc_hd__nor2_1_44/B sky130_fd_sc_hd__nor2_1_44/Y
+ sky130_fd_sc_hd__nor2_1_99/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_55 sky130_fd_sc_hd__or2_0_42/B sky130_fd_sc_hd__nor2_1_55/Y
+ sky130_fd_sc_hd__or2_0_58/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_66 sky130_fd_sc_hd__nor2_1_66/B sky130_fd_sc_hd__nor2_1_66/Y
+ sky130_fd_sc_hd__nor2_1_66/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_77 sky130_fd_sc_hd__buf_6_4/X sky130_fd_sc_hd__nor2_1_77/Y
+ sky130_fd_sc_hd__buf_6_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_88 sky130_fd_sc_hd__nor2_1_88/B sky130_fd_sc_hd__nor2_1_88/Y
+ sky130_fd_sc_hd__nor2_1_88/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_99 sky130_fd_sc_hd__buf_4_1/X sky130_fd_sc_hd__nor2_1_99/Y
+ sky130_fd_sc_hd__nor2_2_5/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_12_504 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_515 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_526 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_410 sky130_fd_sc_hd__nand2_1_410/Y sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__nor2_1_73/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_537 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_421 sky130_fd_sc_hd__nand2_1_421/Y sky130_fd_sc_hd__nand2_1_435/Y
+ sky130_fd_sc_hd__nand2_1_429/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_548 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_432 sky130_fd_sc_hd__nand2_1_432/Y sky130_fd_sc_hd__nand2_1_445/Y
+ sky130_fd_sc_hd__nand2_1_440/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_559 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_443 sky130_fd_sc_hd__nand2_1_443/Y sky130_fd_sc_hd__nand2_1_453/Y
+ sky130_fd_sc_hd__nand2_1_449/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_454 sky130_fd_sc_hd__nand2_1_454/Y sky130_fd_sc_hd__nand2_1_463/Y
+ sky130_fd_sc_hd__nand2_1_459/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_465 sky130_fd_sc_hd__xnor2_1_117/B sky130_fd_sc_hd__nand2_1_466/Y
+ sky130_fd_sc_hd__or2_0_43/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_476 sky130_fd_sc_hd__nand2_1_476/Y sky130_fd_sc_hd__or2_0_50/A
+ sky130_fd_sc_hd__or2_0_50/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_487 sky130_fd_sc_hd__nand2_1_487/Y sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__inv_6_0/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_498 sky130_fd_sc_hd__nand2_1_498/Y sky130_fd_sc_hd__nor2_4_16/Y
+ sky130_fd_sc_hd__or2_0_72/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_12 sky130_fd_sc_hd__nor2_2_31/A sky130_fd_sc_hd__nor2b_1_12/Y
+ sky130_fd_sc_hd__and3_4_26/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_23 sky130_fd_sc_hd__or2_0_84/A sky130_fd_sc_hd__fa_2_445/A
+ sky130_fd_sc_hd__xnor2_2_5/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_34 sky130_fd_sc_hd__fa_2_419/B sky130_fd_sc_hd__fa_2_468/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1001 sky130_fd_sc_hd__clkinv_2_36/A sky130_fd_sc_hd__inv_4_3/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_45 sky130_fd_sc_hd__or2_0_75/B sky130_fd_sc_hd__nor2b_1_45/Y
+ sky130_fd_sc_hd__buf_2_214/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1012 sky130_fd_sc_hd__clkinv_1_1013/A sky130_fd_sc_hd__inv_4_0/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_56 sky130_fd_sc_hd__or2_0_77/A sky130_fd_sc_hd__fa_2_479/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1023 sky130_fd_sc_hd__inv_2_159/A sky130_fd_sc_hd__buf_8_36/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_67 sky130_fd_sc_hd__mux2_2_31/X sky130_fd_sc_hd__nor2b_1_67/Y
+ sky130_fd_sc_hd__mux2_4_5/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1034 sky130_fd_sc_hd__buf_12_5/A sky130_fd_sc_hd__clkinv_1_1034/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_78 sky130_fd_sc_hd__xnor2_2_4/A sky130_fd_sc_hd__fa_2_490/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1045 sky130_fd_sc_hd__inv_2_178/A sky130_fd_sc_hd__inv_2_86/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1503 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2b_1_89 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_89/Y
+ sky130_fd_sc_hd__nor2b_1_89/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1056 sky130_fd_sc_hd__inv_16_1/A sky130_fd_sc_hd__buf_8_55/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1514 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1067 sky130_fd_sc_hd__bufinv_16_1/A sky130_fd_sc_hd__buf_6_74/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_8 vssd1 vccd1 sky130_fd_sc_hd__fa_2_28/A sky130_fd_sc_hd__xnor2_1_8/Y
+ sky130_fd_sc_hd__xnor2_1_8/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_1525 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1078 sky130_fd_sc_hd__maj3_1_1/B la_data_out[41] vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1536 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1089 sky130_fd_sc_hd__o21ai_1_923/A2 sky130_fd_sc_hd__ha_2_60/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1547 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_250 sky130_fd_sc_hd__xor2_1_206/A sky130_fd_sc_hd__clkinv_4_6/Y
+ sky130_fd_sc_hd__and2_0_22/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1558 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_261 sky130_fd_sc_hd__fa_2_110/A sky130_fd_sc_hd__dfxtp_1_264/CLK
+ sky130_fd_sc_hd__and2_0_36/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1569 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_272 sky130_fd_sc_hd__xor2_1_49/A sky130_fd_sc_hd__dfxtp_1_275/CLK
+ sky130_fd_sc_hd__and2_0_94/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_283 sky130_fd_sc_hd__dfxtp_1_283/Q sky130_fd_sc_hd__dfxtp_1_2/CLK
+ sky130_fd_sc_hd__and2_0_259/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_294 sky130_fd_sc_hd__dfxtp_1_294/Q sky130_fd_sc_hd__clkinv_8_6/Y
+ sky130_fd_sc_hd__and2_0_270/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__mux2_4_4 sky130_fd_sc_hd__mux2_4_4/X sky130_fd_sc_hd__mux2_4_4/S
+ sky130_fd_sc_hd__buf_4_25/X sky130_fd_sc_hd__mux2_4_4/A1 vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__mux2_4
Xsky130_fd_sc_hd__o22ai_1_3 sky130_fd_sc_hd__o22ai_1_3/A2 sky130_fd_sc_hd__o22ai_1_3/B1
+ sky130_fd_sc_hd__o22ai_1_3/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__o22ai_1_9/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_100 sky130_fd_sc_hd__fa_2_96/A sky130_fd_sc_hd__fa_2_101/B
+ sky130_fd_sc_hd__fa_2_100/A sky130_fd_sc_hd__fa_2_100/B sky130_fd_sc_hd__xor2_1_137/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_111 sky130_fd_sc_hd__fa_2_108/B sky130_fd_sc_hd__fah_1_0/CI
+ sky130_fd_sc_hd__fa_2_111/A sky130_fd_sc_hd__fa_2_111/B sky130_fd_sc_hd__fah_1_1/COUT
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_122 sky130_fd_sc_hd__fa_2_118/CIN sky130_fd_sc_hd__fa_2_120/A
+ sky130_fd_sc_hd__fa_2_122/A sky130_fd_sc_hd__fa_2_122/B sky130_fd_sc_hd__xor2_1_169/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_133 sky130_fd_sc_hd__fa_2_131/CIN sky130_fd_sc_hd__fa_2_134/B
+ sky130_fd_sc_hd__fa_2_133/A sky130_fd_sc_hd__fa_2_133/B sky130_fd_sc_hd__xor2_1_189/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_144 sky130_fd_sc_hd__xor3_1_12/C sky130_fd_sc_hd__fa_2_146/CIN
+ sky130_fd_sc_hd__fa_2_144/A sky130_fd_sc_hd__fa_2_144/B sky130_fd_sc_hd__xor2_1_228/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_155 sky130_fd_sc_hd__fa_2_146/A sky130_fd_sc_hd__fa_2_156/A
+ sky130_fd_sc_hd__fa_2_155/A sky130_fd_sc_hd__fa_2_155/B sky130_fd_sc_hd__xor2_1_242/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_166 sky130_fd_sc_hd__fa_2_157/A sky130_fd_sc_hd__fa_2_167/B
+ sky130_fd_sc_hd__fa_2_166/A sky130_fd_sc_hd__fa_2_166/B sky130_fd_sc_hd__fa_2_166/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and3_4_5 sky130_fd_sc_hd__and3_4_5/A sky130_fd_sc_hd__and3_4_5/B
+ sky130_fd_sc_hd__and3_4_5/C sky130_fd_sc_hd__and3_4_5/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__fa_2_177 sky130_fd_sc_hd__or2_0_28/A sky130_fd_sc_hd__nor2_2_11/B
+ sky130_fd_sc_hd__fa_2_177/A sky130_fd_sc_hd__fa_2_177/B sky130_fd_sc_hd__fa_2_177/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_188 sky130_fd_sc_hd__fa_2_183/A sky130_fd_sc_hd__fa_2_189/B
+ sky130_fd_sc_hd__fa_2_188/A sky130_fd_sc_hd__fa_2_188/B sky130_fd_sc_hd__fa_2_188/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_199 sky130_fd_sc_hd__fa_2_186/B sky130_fd_sc_hd__fa_2_199/SUM
+ sky130_fd_sc_hd__fa_2_199/A sky130_fd_sc_hd__fa_2_199/B sky130_fd_sc_hd__xor2_1_288/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o22ai_1_10 sky130_fd_sc_hd__o22ai_1_53/B1 sky130_fd_sc_hd__o22ai_1_10/B1
+ sky130_fd_sc_hd__o22ai_1_10/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__o22ai_1_9/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_21 sky130_fd_sc_hd__o22ai_1_42/B1 sky130_fd_sc_hd__o22ai_1_21/B1
+ sky130_fd_sc_hd__o22ai_1_21/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__inv_4_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_32 sky130_fd_sc_hd__nor2_1_33/A sky130_fd_sc_hd__o22ai_1_32/B1
+ sky130_fd_sc_hd__o22ai_1_32/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_150 vccd1 vssd1 sky130_fd_sc_hd__buf_2_150/X sky130_fd_sc_hd__buf_2_150/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_43 sky130_fd_sc_hd__nor2_1_24/A sky130_fd_sc_hd__o22ai_1_43/B1
+ sky130_fd_sc_hd__o22ai_1_43/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_161 vccd1 vssd1 sky130_fd_sc_hd__buf_8_101/A sky130_fd_sc_hd__buf_2_161/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_54 sky130_fd_sc_hd__nor2_1_13/A sky130_fd_sc_hd__o22ai_1_9/A2
+ sky130_fd_sc_hd__o22ai_1_54/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_172 vccd1 vssd1 sky130_fd_sc_hd__ha_2_30/A la_data_out[42]
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_65 sky130_fd_sc_hd__nor2b_1_20/A sky130_fd_sc_hd__xnor2_1_222/Y
+ sky130_fd_sc_hd__fa_2_426/B sky130_fd_sc_hd__xnor2_1_255/Y sky130_fd_sc_hd__o22ai_1_78/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_183 vccd1 vssd1 sky130_fd_sc_hd__buf_2_183/X sky130_fd_sc_hd__inv_2_198/Y
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_76 sky130_fd_sc_hd__xnor2_2_6/Y sky130_fd_sc_hd__xnor2_1_231/Y
+ sky130_fd_sc_hd__fa_2_435/A sky130_fd_sc_hd__xnor2_1_227/Y sky130_fd_sc_hd__o22ai_1_98/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_194 vccd1 vssd1 la_data_out[83] sky130_fd_sc_hd__buf_2_207/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_87 sky130_fd_sc_hd__xnor2_1_235/Y sky130_fd_sc_hd__or2_0_84/A
+ sky130_fd_sc_hd__or2_0_98/A sky130_fd_sc_hd__inv_2_65/Y sky130_fd_sc_hd__o22ai_1_99/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_98 sky130_fd_sc_hd__xnor2_2_6/Y sky130_fd_sc_hd__xnor2_1_250/Y
+ sky130_fd_sc_hd__fa_2_446/A sky130_fd_sc_hd__xnor2_1_246/Y sky130_fd_sc_hd__o22ai_1_98/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_4_12 vccd1 vssd1 sky130_fd_sc_hd__buf_4_12/X sky130_fd_sc_hd__buf_4_12/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_23 vccd1 vssd1 sky130_fd_sc_hd__buf_4_23/X sky130_fd_sc_hd__buf_4_23/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_34 vccd1 vssd1 sky130_fd_sc_hd__buf_4_34/X sky130_fd_sc_hd__buf_4_34/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_12_105 sky130_fd_sc_hd__buf_8_148/X sky130_fd_sc_hd__buf_12_297/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_116 sky130_fd_sc_hd__buf_8_64/X sky130_fd_sc_hd__buf_12_434/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_127 sky130_fd_sc_hd__buf_8_42/X sky130_fd_sc_hd__buf_12_127/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_50 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_50/X sky130_fd_sc_hd__clkbuf_1_52/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_138 sky130_fd_sc_hd__buf_12_18/X sky130_fd_sc_hd__buf_12_324/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_61 vssd1 vccd1 sky130_fd_sc_hd__buf_12_50/A sky130_fd_sc_hd__buf_2_61/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_149 sky130_fd_sc_hd__buf_8_51/X sky130_fd_sc_hd__buf_12_348/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_72 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_9/A1 sky130_fd_sc_hd__clkbuf_1_72/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_83 vssd1 vccd1 sky130_fd_sc_hd__mux2_4_1/A1 sky130_fd_sc_hd__clkbuf_1_83/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_94 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_40/A1 sky130_fd_sc_hd__clkbuf_1_94/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_4_8 sky130_fd_sc_hd__clkbuf_4_8/X sky130_fd_sc_hd__clkbuf_4_8/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_1_305 sky130_fd_sc_hd__nand3_1_4/A sky130_fd_sc_hd__ha_2_3/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_316 sky130_fd_sc_hd__nor2_1_45/A sky130_fd_sc_hd__nand2_1_178/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_327 sky130_fd_sc_hd__nand2_1_184/A sky130_fd_sc_hd__nor2_1_52/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_338 sky130_fd_sc_hd__nand2_1_197/B sky130_fd_sc_hd__nor2_1_57/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_349 sky130_fd_sc_hd__nor2_1_63/A sky130_fd_sc_hd__nand2_1_221/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__or2_0_30 sky130_fd_sc_hd__or2_0_30/A sky130_fd_sc_hd__or2_0_30/X
+ sky130_fd_sc_hd__or2_0_30/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_41 sky130_fd_sc_hd__or2_0_66/A sky130_fd_sc_hd__or2_0_41/X
+ sky130_fd_sc_hd__or2_0_60/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_52 sky130_fd_sc_hd__or2_0_53/A sky130_fd_sc_hd__or2_0_52/X
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_63 sky130_fd_sc_hd__buf_4_3/X sky130_fd_sc_hd__or2_0_63/X
+ sky130_fd_sc_hd__buf_4_2/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_74 sky130_fd_sc_hd__or2_0_74/A sky130_fd_sc_hd__or2_0_74/X
+ sky130_fd_sc_hd__or2_0_74/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__clkinv_4_8 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkinv_4_8/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__or2_0_85 sky130_fd_sc_hd__or2_0_85/A sky130_fd_sc_hd__or2_0_85/X
+ sky130_fd_sc_hd__or2_0_85/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_96 sky130_fd_sc_hd__or2_0_96/A sky130_fd_sc_hd__or2_0_96/X
+ sky130_fd_sc_hd__or2_0_96/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__clkinv_4_110 sky130_fd_sc_hd__clkinv_4_110/A sky130_fd_sc_hd__clkinv_4_114/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_12_650 sky130_fd_sc_hd__buf_12_650/A sky130_fd_sc_hd__buf_12_650/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_4_121 sky130_fd_sc_hd__clkinv_8_83/Y sky130_fd_sc_hd__clkinv_8_84/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_12_661 sky130_fd_sc_hd__buf_12_661/A sky130_fd_sc_hd__buf_12_661/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_672 sky130_fd_sc_hd__buf_12_672/A sky130_fd_sc_hd__buf_12_672/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_301 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_312 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_323 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_334 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_345 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_356 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_240 sky130_fd_sc_hd__nand2_1_240/Y sky130_fd_sc_hd__nand2_1_253/Y
+ sky130_fd_sc_hd__nand2_1_247/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_367 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_251 sky130_fd_sc_hd__nand2_1_251/Y sky130_fd_sc_hd__nor2_1_78/Y
+ sky130_fd_sc_hd__nand2_1_256/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_378 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_850 sky130_fd_sc_hd__clkinv_1_850/Y sky130_fd_sc_hd__clkinv_8_8/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_262 sky130_fd_sc_hd__nor2_1_74/B sky130_fd_sc_hd__nor2_1_84/Y
+ sky130_fd_sc_hd__nor2_1_89/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_389 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_861 sky130_fd_sc_hd__clkinv_1_861/Y sky130_fd_sc_hd__inv_2_196/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_273 sky130_fd_sc_hd__xnor2_1_47/A sky130_fd_sc_hd__nand2_1_274/Y
+ sky130_fd_sc_hd__nand2_1_273/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_872 sky130_fd_sc_hd__buf_2_37/A sky130_fd_sc_hd__clkinv_4_84/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_284 sky130_fd_sc_hd__nand2_1_284/Y sky130_fd_sc_hd__nor2_1_96/Y
+ sky130_fd_sc_hd__nor2_1_44/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_883 sky130_fd_sc_hd__clkinv_1_883/Y sky130_fd_sc_hd__clkinv_4_87/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_295 sky130_fd_sc_hd__nand2_1_295/Y sky130_fd_sc_hd__or2_0_16/A
+ sky130_fd_sc_hd__or2_0_16/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_894 sky130_fd_sc_hd__clkinv_1_894/Y sky130_fd_sc_hd__clkinv_1_894/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1300 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_2_0 vccd1 vssd1 sky130_fd_sc_hd__xor2_2_0/X sky130_fd_sc_hd__xor2_2_0/B
+ sky130_fd_sc_hd__xor2_2_0/A vssd1 vccd1 sky130_fd_sc_hd__xor2_2
Xsky130_fd_sc_hd__decap_12_1311 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_50 sky130_fd_sc_hd__conb_1_50/LO sky130_fd_sc_hd__conb_1_50/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1322 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_61 sky130_fd_sc_hd__conb_1_61/LO sky130_fd_sc_hd__conb_1_61/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1333 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_72 sky130_fd_sc_hd__conb_1_72/LO sky130_fd_sc_hd__conb_1_72/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1344 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_83 sky130_fd_sc_hd__conb_1_83/LO sky130_fd_sc_hd__conb_1_83/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1355 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_94 sky130_fd_sc_hd__conb_1_94/LO sky130_fd_sc_hd__conb_1_94/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1366 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1377 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_808 vssd1 vccd1 sky130_fd_sc_hd__inv_2_52/Y sky130_fd_sc_hd__nand2_1_599/Y
+ sky130_fd_sc_hd__a21oi_1_124/Y sky130_fd_sc_hd__xor2_2_2/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1388 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_819 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_9/X sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__o21ai_1_819/B1 sky130_fd_sc_hd__xor2_1_592/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1399 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__mux2_2_1 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_1/A1 sky130_fd_sc_hd__mux2_2_1/A0
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__or2_0_77/A vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__decap_12_890 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2b_2_9 la_data_out[36] sky130_fd_sc_hd__nand2b_2_9/Y la_data_out[56]
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_2
Xsky130_fd_sc_hd__xor2_1_602 sky130_fd_sc_hd__xor2_1_602/B sky130_fd_sc_hd__xor2_1_602/X
+ sky130_fd_sc_hd__xor2_1_602/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_613 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__xor2_1_613/X
+ sky130_fd_sc_hd__xor2_1_613/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_624 sky130_fd_sc_hd__xor2_1_624/B sky130_fd_sc_hd__xor2_1_624/X
+ sky130_fd_sc_hd__xor2_1_624/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_635 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__xor2_1_635/X
+ sky130_fd_sc_hd__xor2_1_635/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_646 sky130_fd_sc_hd__xor2_1_646/B sky130_fd_sc_hd__xor2_1_646/X
+ sky130_fd_sc_hd__xor2_1_646/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_657 sky130_fd_sc_hd__xor2_1_657/B sky130_fd_sc_hd__xor2_1_657/X
+ sky130_fd_sc_hd__xor2_1_657/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_668 sky130_fd_sc_hd__mux2_4_4/X sky130_fd_sc_hd__xor2_1_668/X
+ sky130_fd_sc_hd__xnor2_2_4/B vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_679 sky130_fd_sc_hd__xor2_1_679/B sky130_fd_sc_hd__xor2_1_679/X
+ sky130_fd_sc_hd__xor2_1_679/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__fa_2_9 sky130_fd_sc_hd__fa_2_8/B sky130_fd_sc_hd__fa_2_9/SUM sky130_fd_sc_hd__fa_2_9/A
+ sky130_fd_sc_hd__fa_2_9/B sky130_fd_sc_hd__fa_2_9/CIN vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a211o_1_15 vssd1 vccd1 sky130_fd_sc_hd__fa_2_250/B sky130_fd_sc_hd__dfxtp_1_78/Q
+ sky130_fd_sc_hd__nor2_1_19/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_15/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__a211o_1_26 vssd1 vccd1 sky130_fd_sc_hd__fa_2_179/A sky130_fd_sc_hd__dfxtp_1_89/Q
+ sky130_fd_sc_hd__nor2_1_30/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_26/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__clkinv_1_102 io_oeb[37] sky130_fd_sc_hd__conb_1_40/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_113 io_oeb[26] sky130_fd_sc_hd__conb_1_29/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_124 io_oeb[15] sky130_fd_sc_hd__conb_1_18/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_135 io_oeb[4] sky130_fd_sc_hd__conb_1_7/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_146 sky130_fd_sc_hd__and2_0_251/A sky130_fd_sc_hd__a222oi_1_47/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_157 sky130_fd_sc_hd__o22ai_1_34/B1 sky130_fd_sc_hd__dfxtp_1_186/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_168 sky130_fd_sc_hd__o21ai_1_7/A2 sky130_fd_sc_hd__dfxtp_1_120/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_179 sky130_fd_sc_hd__nor2_1_26/A sky130_fd_sc_hd__dfxtp_1_149/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_15 sky130_fd_sc_hd__inv_2_66/Y sky130_fd_sc_hd__or2_0_90/B
+ sky130_fd_sc_hd__a22o_1_15/X sky130_fd_sc_hd__nor2_1_233/Y sky130_fd_sc_hd__xor2_1_655/X
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_26 sky130_fd_sc_hd__buf_2_63/A sky130_fd_sc_hd__buf_2_101/X
+ sky130_fd_sc_hd__a22o_1_26/X sky130_fd_sc_hd__a22o_1_26/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_37 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__buf_2_112/X
+ sky130_fd_sc_hd__a22o_1_37/X sky130_fd_sc_hd__a22o_1_37/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_48 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__a22o_1_48/A2
+ sky130_fd_sc_hd__a22o_1_48/X sky130_fd_sc_hd__a22o_1_48/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__o21ai_1_2 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_2/A2 sky130_fd_sc_hd__nor2_4_4/B
+ sky130_fd_sc_hd__o21ai_1_2/B1 sky130_fd_sc_hd__fa_2_12/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a22o_1_59 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__buf_2_49/A
+ sky130_fd_sc_hd__a22o_1_59/X sky130_fd_sc_hd__ha_2_30/SUM sky130_fd_sc_hd__a22o_1_71/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__nor2_1_240 sky130_fd_sc_hd__nor2_1_240/B sky130_fd_sc_hd__nor2_1_240/Y
+ sky130_fd_sc_hd__nor2_1_240/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_251 sky130_fd_sc_hd__nor2_1_251/B sky130_fd_sc_hd__nor2_1_251/Y
+ sky130_fd_sc_hd__nor2_1_251/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_2_5 sky130_fd_sc_hd__clkinv_2_5/Y sky130_fd_sc_hd__clkinv_2_5/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__nor2_1_262 sky130_fd_sc_hd__nor2_1_262/B sky130_fd_sc_hd__nor2_1_262/Y
+ sky130_fd_sc_hd__nor2_1_262/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_273 sky130_fd_sc_hd__nor2_1_273/B sky130_fd_sc_hd__nor2_1_273/Y
+ sky130_fd_sc_hd__nor2_1_273/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_284 sky130_fd_sc_hd__or3_1_0/X sky130_fd_sc_hd__a21o_2_2/B1
+ wbs_adr_i[5] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_480 sky130_fd_sc_hd__buf_12_480/A sky130_fd_sc_hd__buf_12_538/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_491 sky130_fd_sc_hd__buf_12_491/A sky130_fd_sc_hd__buf_12_517/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_120 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_131 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_142 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_153 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_164 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_175 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_210 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_210/B sky130_fd_sc_hd__a22o_1_11/B1
+ sky130_fd_sc_hd__xnor2_1_210/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_186 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_16 sky130_fd_sc_hd__nand2_1_16/Y sky130_fd_sc_hd__nand2_1_16/B
+ sky130_fd_sc_hd__nand2_1_16/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_221 vssd1 vccd1 sky130_fd_sc_hd__buf_2_207/X sky130_fd_sc_hd__xnor2_1_221/Y
+ sky130_fd_sc_hd__buf_4_41/X vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_197 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_27 sky130_fd_sc_hd__nand2_1_27/Y sky130_fd_sc_hd__nand2_1_8/B
+ sky130_fd_sc_hd__or2_0_79/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_232 vssd1 vccd1 sky130_fd_sc_hd__buf_2_207/X sky130_fd_sc_hd__xnor2_1_232/Y
+ la_data_out[68] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_680 sky130_fd_sc_hd__nand2_1_757/A sky130_fd_sc_hd__nor2_1_243/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_38 sky130_fd_sc_hd__nand2_1_38/Y sky130_fd_sc_hd__nand2_1_8/B
+ sky130_fd_sc_hd__or2_0_81/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_243 vssd1 vccd1 sky130_fd_sc_hd__buf_2_207/X sky130_fd_sc_hd__xnor2_1_243/Y
+ la_data_out[67] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_49 sky130_fd_sc_hd__nor2_1_0/A sky130_fd_sc_hd__nor2_4_0/B
+ sky130_fd_sc_hd__nor2_4_0/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_691 sky130_fd_sc_hd__nand2_1_765/A sky130_fd_sc_hd__nor2_1_249/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_254 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_5/B sky130_fd_sc_hd__xnor2_1_254/Y
+ sky130_fd_sc_hd__or2_1_10/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_265 vssd1 vccd1 sky130_fd_sc_hd__buf_2_207/X sky130_fd_sc_hd__xnor2_1_265/Y
+ la_data_out[72] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_276 vssd1 vccd1 sky130_fd_sc_hd__buf_2_207/X sky130_fd_sc_hd__xnor2_1_276/Y
+ sky130_fd_sc_hd__mux2_4_2/X vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_287 vssd1 vccd1 la_data_out[67] sky130_fd_sc_hd__xnor2_1_287/Y
+ sky130_fd_sc_hd__or2_0_77/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_298 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_298/B sky130_fd_sc_hd__xnor2_1_298/Y
+ sky130_fd_sc_hd__xnor2_1_298/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_1130 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1141 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1152 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1163 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1174 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_605 vssd1 vccd1 sky130_fd_sc_hd__buf_2_11/X sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_605/B1 sky130_fd_sc_hd__xor2_1_397/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1185 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_616 vssd1 vccd1 sky130_fd_sc_hd__inv_2_27/Y sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__nand2_1_330/Y sky130_fd_sc_hd__xor2_1_408/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1196 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_627 vssd1 vccd1 sky130_fd_sc_hd__buf_2_7/X sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_627/B1 sky130_fd_sc_hd__xor2_1_420/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_638 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_861/A2 sky130_fd_sc_hd__nand2b_2_6/Y
+ sky130_fd_sc_hd__nand2_1_498/Y sky130_fd_sc_hd__xor2_1_608/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_649 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_649/A2 sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_649/B1 sky130_fd_sc_hd__xor2_1_436/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fah_1_3 sky130_fd_sc_hd__nor2_2_14/A sky130_fd_sc_hd__fah_1_3/B
+ sky130_fd_sc_hd__fah_1_3/A sky130_fd_sc_hd__or2_0_37/B sky130_fd_sc_hd__fah_1_3/CI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__fah_1
Xsky130_fd_sc_hd__sdlclkp_2_10 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_8_61/Y
+ sky130_fd_sc_hd__dfxtp_4_3/CLK sky130_fd_sc_hd__o21ai_2_2/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__xor2_1_410 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__or2_0_43/A
+ sky130_fd_sc_hd__xor2_1_410/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_80 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_80/B sky130_fd_sc_hd__xnor2_1_80/Y
+ sky130_fd_sc_hd__xnor2_1_80/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_421 sky130_fd_sc_hd__o21a_1_3/A1 sky130_fd_sc_hd__xor2_1_421/X
+ sky130_fd_sc_hd__xor2_1_421/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_91 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_91/B sky130_fd_sc_hd__xnor2_1_91/Y
+ sky130_fd_sc_hd__xnor2_1_91/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_432 sky130_fd_sc_hd__fa_2_389/A sky130_fd_sc_hd__xor3_1_28/B
+ sky130_fd_sc_hd__xor2_1_432/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_443 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__fa_2_284/A
+ sky130_fd_sc_hd__xor2_1_443/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_454 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__fa_2_293/B
+ sky130_fd_sc_hd__xor2_1_454/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_465 sky130_fd_sc_hd__fah_1_14/A sky130_fd_sc_hd__fa_2_303/A
+ sky130_fd_sc_hd__xor2_1_465/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_476 sky130_fd_sc_hd__xor2_1_548/B sky130_fd_sc_hd__fa_2_311/A
+ sky130_fd_sc_hd__xor2_1_476/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_487 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__xor2_1_487/X
+ sky130_fd_sc_hd__xor2_1_487/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_498 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__fa_2_332/B
+ sky130_fd_sc_hd__xor2_1_498/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a222oi_1_507 vccd1 vssd1 sky130_fd_sc_hd__and3_4_20/X sky130_fd_sc_hd__buf_2_30/X
+ sky130_fd_sc_hd__buf_2_26/X sky130_fd_sc_hd__nor2_4_16/Y sky130_fd_sc_hd__buf_2_24/X
+ sky130_fd_sc_hd__o21ai_1_805/B1 sky130_fd_sc_hd__and2b_4_11/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_518 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__buf_2_20/X
+ sky130_fd_sc_hd__buf_2_21/X sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__o21ai_1_817/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_529 vccd1 vssd1 sky130_fd_sc_hd__and3_4_21/X sky130_fd_sc_hd__buf_2_25/A
+ sky130_fd_sc_hd__inv_6_0/Y sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__buf_8_0/A
+ sky130_fd_sc_hd__o21ai_1_836/B1 sky130_fd_sc_hd__and2b_4_12/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nor2b_1_107 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_107/Y
+ sky130_fd_sc_hd__nor2b_1_107/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_118 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_118/Y
+ sky130_fd_sc_hd__nor2b_1_118/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_129 sky130_fd_sc_hd__clkinv_4_48/Y sky130_fd_sc_hd__nor2b_1_129/Y
+ wb_rst_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__buf_6_8 vccd1 vssd1 sky130_fd_sc_hd__buf_6_8/X sky130_fd_sc_hd__buf_6_8/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__clkinv_2_10 sky130_fd_sc_hd__clkinv_4_6/A sky130_fd_sc_hd__clkinv_2_10/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_21 sky130_fd_sc_hd__inv_2_115/A sky130_fd_sc_hd__buf_8_99/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_32 sky130_fd_sc_hd__clkinv_2_32/Y sky130_fd_sc_hd__clkinv_2_32/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_43 sky130_fd_sc_hd__inv_2_171/A sky130_fd_sc_hd__inv_2_169/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__and2_0_401 vccd1 vssd1 sky130_fd_sc_hd__edfxbp_1_0/D sky130_fd_sc_hd__and2_0_401/B
+ sky130_fd_sc_hd__nor2_1_273/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_2_54 sky130_fd_sc_hd__inv_8_3/A sky130_fd_sc_hd__nand2_1_14/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__or2_1_3 sky130_fd_sc_hd__or2_1_3/A sky130_fd_sc_hd__or2_1_3/X sky130_fd_sc_hd__or2_1_3/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_1
Xsky130_fd_sc_hd__sdlclkp_4_6 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_4_0/Y
+ sky130_fd_sc_hd__dfxtp_1_94/CLK sky130_fd_sc_hd__o21ai_2_0/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_9 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_9/Y
+ sky130_fd_sc_hd__nor2_1_9/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_180 sky130_fd_sc_hd__xor2_1_411/X sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xor2_1_199/X sky130_fd_sc_hd__a22oi_1_180/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_191 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__nor2b_1_2/Y sky130_fd_sc_hd__nor2_1_48/Y sky130_fd_sc_hd__a22oi_1_191/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22o_4_0 sky130_fd_sc_hd__nand2_1_8/B sky130_fd_sc_hd__or2_0_73/A
+ sky130_fd_sc_hd__or2_0_61/A sky130_fd_sc_hd__or2_0_73/B sky130_fd_sc_hd__nand2_1_7/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_4
Xsky130_fd_sc_hd__o21ai_1_402 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_505/A2 sky130_fd_sc_hd__nand2b_2_3/Y
+ sky130_fd_sc_hd__o21ai_1_402/B1 sky130_fd_sc_hd__xor2_1_214/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_413 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_7/X sky130_fd_sc_hd__or2_0_32/X
+ sky130_fd_sc_hd__o21a_1_2/X sky130_fd_sc_hd__xnor2_1_69/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_424 vssd1 vccd1 sky130_fd_sc_hd__inv_2_41/Y sky130_fd_sc_hd__nand2b_2_3/Y
+ sky130_fd_sc_hd__o21ai_1_424/B1 sky130_fd_sc_hd__xor2_1_231/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_435 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_7/X sky130_fd_sc_hd__nand2_1_346/Y
+ sky130_fd_sc_hd__a21oi_1_75/Y sky130_fd_sc_hd__xnor2_1_72/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_446 vssd1 vccd1 sky130_fd_sc_hd__buf_2_8/X sky130_fd_sc_hd__nand2b_1_13/Y
+ sky130_fd_sc_hd__o21ai_1_446/B1 sky130_fd_sc_hd__xor2_1_249/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_457 vssd1 vccd1 sky130_fd_sc_hd__inv_2_40/Y sky130_fd_sc_hd__nand2b_2_3/Y
+ sky130_fd_sc_hd__o21ai_1_457/B1 sky130_fd_sc_hd__xor2_1_259/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_468 vssd1 vccd1 sky130_fd_sc_hd__buf_2_7/X sky130_fd_sc_hd__nand2b_1_12/Y
+ sky130_fd_sc_hd__o21ai_1_468/B1 sky130_fd_sc_hd__xor2_1_271/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_479 vssd1 vccd1 sky130_fd_sc_hd__buf_2_8/X sky130_fd_sc_hd__nand2b_1_14/Y
+ sky130_fd_sc_hd__o21ai_1_479/B1 sky130_fd_sc_hd__xor2_1_280/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2_4_11 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__or2b_2_1/A
+ sky130_fd_sc_hd__and3_4_9/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__nand2_1_806 sky130_fd_sc_hd__xnor2_1_294/A sky130_fd_sc_hd__nand2_1_807/Y
+ sky130_fd_sc_hd__or2_0_103/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_817 sky130_fd_sc_hd__nand2_1_817/Y sky130_fd_sc_hd__nor2_1_260/A
+ sky130_fd_sc_hd__nor2_1_260/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_828 sky130_fd_sc_hd__xor2_1_685/B sky130_fd_sc_hd__nand2_1_829/Y
+ sky130_fd_sc_hd__nand2_1_828/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_839 sky130_fd_sc_hd__nand2_1_839/Y sky130_fd_sc_hd__or2_0_111/A
+ sky130_fd_sc_hd__or2_0_111/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o21ai_1_17 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_16/B1 sky130_fd_sc_hd__inv_2_53/A
+ sky130_fd_sc_hd__o21ai_1_17/B1 sky130_fd_sc_hd__fa_2_104/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_240 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__xor2_1_240/X
+ sky130_fd_sc_hd__xor2_1_240/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__o21ai_1_28 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_5/B1 sky130_fd_sc_hd__nor2_4_4/B
+ sky130_fd_sc_hd__o21ai_1_28/B1 sky130_fd_sc_hd__fa_2_139/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_251 sky130_fd_sc_hd__fa_2_170/A sky130_fd_sc_hd__fa_2_161/B
+ sky130_fd_sc_hd__xor2_1_251/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__o21ai_1_39 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_41/A2 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_87/Y sky130_fd_sc_hd__and2_0_14/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_262 sky130_fd_sc_hd__fa_2_170/A sky130_fd_sc_hd__and3_1_1/B
+ sky130_fd_sc_hd__xor2_1_262/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_273 sky130_fd_sc_hd__dfxtp_2_5/Q sky130_fd_sc_hd__fa_2_182/A
+ sky130_fd_sc_hd__xor2_1_273/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_284 sky130_fd_sc_hd__fa_2_250/A sky130_fd_sc_hd__xor2_1_284/X
+ sky130_fd_sc_hd__xor2_1_284/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_295 sky130_fd_sc_hd__fa_2_250/A sky130_fd_sc_hd__fa_2_195/A
+ sky130_fd_sc_hd__xor2_1_295/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_200 vssd1 vccd1 sky130_fd_sc_hd__buf_12_27/A sky130_fd_sc_hd__inv_12_0/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_211 vssd1 vccd1 sky130_fd_sc_hd__buf_8_24/A sky130_fd_sc_hd__buf_2_61/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_222 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_54/A1 sky130_fd_sc_hd__clkbuf_1_222/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_233 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_39/A1 sky130_fd_sc_hd__clkbuf_1_233/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_304 vccd1 vssd1 sky130_fd_sc_hd__and3_4_10/X sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__buf_6_1/X sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__and2_0_38/A
+ sky130_fd_sc_hd__o21ai_1_519/B1 sky130_fd_sc_hd__and2b_4_7/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_244 vssd1 vccd1 sky130_fd_sc_hd__buf_8_115/A sky130_fd_sc_hd__clkbuf_1_302/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_315 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__buf_4_2/X sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__o21ai_1_530/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_255 vssd1 vccd1 sky130_fd_sc_hd__buf_12_52/A sky130_fd_sc_hd__clkbuf_1_255/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_2_2 sky130_fd_sc_hd__fah_1_14/A sky130_fd_sc_hd__dfxtp_2_2/CLK
+ sky130_fd_sc_hd__dfxtp_2_2/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_2
Xsky130_fd_sc_hd__a222oi_1_326 vccd1 vssd1 sky130_fd_sc_hd__and3_4_16/X sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__inv_6_0/Y sky130_fd_sc_hd__nor2_2_19/Y sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__o21ai_1_545/B1 sky130_fd_sc_hd__nor2b_2_3/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_266 vssd1 vccd1 sky130_fd_sc_hd__buf_8_129/A sky130_fd_sc_hd__clkbuf_1_34/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_337 vccd1 vssd1 sky130_fd_sc_hd__and3_4_11/X sky130_fd_sc_hd__buf_2_31/X
+ sky130_fd_sc_hd__buf_2_19/X sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__o21ai_1_559/B1 sky130_fd_sc_hd__and2b_4_8/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_277 vssd1 vccd1 sky130_fd_sc_hd__buf_8_144/A sky130_fd_sc_hd__clkbuf_1_277/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_348 vccd1 vssd1 sky130_fd_sc_hd__and3_4_10/X sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__buf_6_2/X sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__buf_4_7/X
+ sky130_fd_sc_hd__o21ai_1_575/B1 sky130_fd_sc_hd__and2b_4_7/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_288 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_288/X sky130_fd_sc_hd__clkbuf_1_288/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_359 vccd1 vssd1 sky130_fd_sc_hd__and3_4_11/X sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__buf_6_2/X sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__buf_4_7/X
+ sky130_fd_sc_hd__o21ai_1_593/B1 sky130_fd_sc_hd__and2b_4_8/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_299 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_299/X sky130_fd_sc_hd__clkbuf_1_299/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_4_5 vccd1 vssd1 sky130_fd_sc_hd__buf_4_5/X sky130_fd_sc_hd__buf_4_5/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__and2_0_220 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_86/D sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__o21ai_1_66/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_231 vccd1 vssd1 sky130_fd_sc_hd__and2_0_231/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_231/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_242 vccd1 vssd1 sky130_fd_sc_hd__and2_0_242/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__o21ai_1_49/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_253 vccd1 vssd1 sky130_fd_sc_hd__and2_0_253/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__and2_0_253/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_264 vccd1 vssd1 sky130_fd_sc_hd__and2_0_264/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__xor2_1_646/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_275 vccd1 vssd1 sky130_fd_sc_hd__and2_0_275/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__and2_0_275/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__a21oi_2_16 sky130_fd_sc_hd__a21oi_2_16/B1 sky130_fd_sc_hd__or2_1_6/X
+ sky130_fd_sc_hd__xnor2_1_145/B sky130_fd_sc_hd__xor2_1_489/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_2
Xsky130_fd_sc_hd__and2_0_286 vccd1 vssd1 sky130_fd_sc_hd__and2_0_286/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_7/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_297 vccd1 vssd1 sky130_fd_sc_hd__and2_0_297/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_18/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__sdlclkp_2_3 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_4_0/Y
+ sky130_fd_sc_hd__dfxtp_1_126/CLK sky130_fd_sc_hd__clkbuf_1_11/X vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__inv_4_5 sky130_fd_sc_hd__inv_4_5/Y sky130_fd_sc_hd__inv_4_5/A vccd1
+ vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__o21ai_1_210 vssd1 vccd1 sky130_fd_sc_hd__inv_2_23/Y sky130_fd_sc_hd__nand2b_2_0/Y
+ sky130_fd_sc_hd__a222oi_1_82/Y sky130_fd_sc_hd__xor2_1_35/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_221 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_59/Y sky130_fd_sc_hd__nor2_1_54/A
+ sky130_fd_sc_hd__nor2_1_53/Y sky130_fd_sc_hd__o21ai_1_221/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_232 vssd1 vccd1 sky130_fd_sc_hd__inv_2_9/Y sky130_fd_sc_hd__nand2b_1_7/Y
+ sky130_fd_sc_hd__o21ai_1_232/B1 sky130_fd_sc_hd__xor2_1_57/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_50 la_data_out[84] sky130_fd_sc_hd__mux2_2_48/X vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_243 vssd1 vccd1 sky130_fd_sc_hd__inv_2_23/Y sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__o21ai_1_243/B1 sky130_fd_sc_hd__xor2_1_66/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_254 vssd1 vccd1 sky130_fd_sc_hd__buf_2_3/X sky130_fd_sc_hd__nand2b_1_5/Y
+ sky130_fd_sc_hd__o21ai_1_254/B1 sky130_fd_sc_hd__xor2_1_76/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_265 vssd1 vccd1 sky130_fd_sc_hd__inv_2_18/Y sky130_fd_sc_hd__nand2b_1_7/Y
+ sky130_fd_sc_hd__o21ai_1_265/B1 sky130_fd_sc_hd__xor2_1_87/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_276 vssd1 vccd1 sky130_fd_sc_hd__inv_2_17/Y sky130_fd_sc_hd__nand2b_1_1/Y
+ sky130_fd_sc_hd__o21ai_1_276/B1 sky130_fd_sc_hd__xor2_1_97/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_287 vssd1 vccd1 sky130_fd_sc_hd__inv_2_19/Y sky130_fd_sc_hd__nand2b_1_1/Y
+ sky130_fd_sc_hd__o21ai_1_287/B1 sky130_fd_sc_hd__xor2_1_108/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_298 vssd1 vccd1 sky130_fd_sc_hd__inv_2_12/Y sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__o21ai_1_298/B1 sky130_fd_sc_hd__xor2_1_119/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_708 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_719 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_603 sky130_fd_sc_hd__nand2_1_603/Y sky130_fd_sc_hd__nand2_1_616/Y
+ sky130_fd_sc_hd__nand2_1_611/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_614 sky130_fd_sc_hd__nand2_1_614/Y sky130_fd_sc_hd__nand2_1_624/Y
+ sky130_fd_sc_hd__nand2_1_620/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_625 sky130_fd_sc_hd__nand2_1_625/Y sky130_fd_sc_hd__nand2_1_634/Y
+ sky130_fd_sc_hd__nand2_1_630/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_636 sky130_fd_sc_hd__xnor2_1_179/B sky130_fd_sc_hd__nand2_1_637/Y
+ sky130_fd_sc_hd__or2_0_62/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_647 sky130_fd_sc_hd__nand2_1_647/Y sky130_fd_sc_hd__or2_0_68/A
+ sky130_fd_sc_hd__or2_0_68/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_658 sky130_fd_sc_hd__xor2_1_634/A sky130_fd_sc_hd__o21a_1_5/B1
+ sky130_fd_sc_hd__nand2_1_658/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_669 sky130_fd_sc_hd__nand2_1_669/Y sky130_fd_sc_hd__mux2_2_20/X
+ sky130_fd_sc_hd__mux2_2_43/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_2_5 sky130_fd_sc_hd__nor2_2_32/A sky130_fd_sc_hd__nor2b_2_5/A
+ sky130_fd_sc_hd__nor2b_2_5/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_2
Xsky130_fd_sc_hd__decap_12_1707 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_410 sky130_fd_sc_hd__dfxtp_1_410/Q sky130_fd_sc_hd__dfxtp_1_410/CLK
+ sky130_fd_sc_hd__nor2b_1_105/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1718 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_17 sky130_fd_sc_hd__inv_2_17/A sky130_fd_sc_hd__inv_2_17/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_421 sky130_fd_sc_hd__dfxtp_1_421/Q sky130_fd_sc_hd__dfxtp_1_427/CLK
+ sky130_fd_sc_hd__nor2b_1_94/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1729 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_28 sky130_fd_sc_hd__inv_2_28/A sky130_fd_sc_hd__inv_2_28/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_432 sky130_fd_sc_hd__dfxtp_1_432/Q sky130_fd_sc_hd__clkinv_4_9/Y
+ sky130_fd_sc_hd__nor2b_1_115/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_39 sky130_fd_sc_hd__inv_2_39/A sky130_fd_sc_hd__inv_2_39/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_443 sky130_fd_sc_hd__dfxtp_1_443/Q sky130_fd_sc_hd__dfxtp_1_446/CLK
+ sky130_fd_sc_hd__nor2b_1_104/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_454 sky130_fd_sc_hd__dfxtp_1_454/Q sky130_fd_sc_hd__clkinv_4_9/Y
+ sky130_fd_sc_hd__nor2b_1_93/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_465 sky130_fd_sc_hd__ha_2_49/A sky130_fd_sc_hd__dfxtp_1_520/CLK
+ sky130_fd_sc_hd__and2_0_360/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_476 sky130_fd_sc_hd__dfxtp_1_476/Q sky130_fd_sc_hd__dfxtp_1_480/CLK
+ sky130_fd_sc_hd__and2_0_389/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_487 la_data_out[54] sky130_fd_sc_hd__dfxtp_1_489/CLK sky130_fd_sc_hd__and2_0_372/X
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_2_7 sky130_fd_sc_hd__nand2_2_7/Y sky130_fd_sc_hd__nand2_2_7/A
+ sky130_fd_sc_hd__nand2_2_7/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__dfxtp_1_498 la_data_out[47] sky130_fd_sc_hd__dfxtp_1_498/CLK sky130_fd_sc_hd__and2_0_380/X
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a222oi_1_101 vccd1 vssd1 sky130_fd_sc_hd__and3_4_4/X sky130_fd_sc_hd__clkbuf_1_3/X
+ sky130_fd_sc_hd__or2_0_53/A sky130_fd_sc_hd__nor2_1_61/Y sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__o21ai_1_233/B1 sky130_fd_sc_hd__nor2b_1_4/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2b_1_13 sky130_fd_sc_hd__nand2b_1_13/Y sky130_fd_sc_hd__and3_4_14/C
+ sky130_fd_sc_hd__and3_4_14/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a222oi_1_112 vccd1 vssd1 sky130_fd_sc_hd__and3_4_7/X sky130_fd_sc_hd__nor2_2_4/B
+ sky130_fd_sc_hd__buf_2_4/X sky130_fd_sc_hd__nor2_2_7/Y sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__o21ai_1_248/B1 sky130_fd_sc_hd__nor2b_2_1/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2b_1_24 sky130_fd_sc_hd__nand2b_1_24/Y sky130_fd_sc_hd__or2_0_84/A
+ la_data_out[77] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a222oi_1_123 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__or2_0_66/A sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__or2_0_60/B
+ sky130_fd_sc_hd__o21ai_1_261/B1 sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_134 vccd1 vssd1 sky130_fd_sc_hd__and3_4_8/X sky130_fd_sc_hd__nor2_2_4/B
+ sky130_fd_sc_hd__buf_2_4/X sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__o21ai_1_276/B1 sky130_fd_sc_hd__nor2b_2_2/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_145 vccd1 vssd1 sky130_fd_sc_hd__and3_4_8/X sky130_fd_sc_hd__nor2_2_5/A
+ sky130_fd_sc_hd__nor2_2_5/B sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__nor2_2_4/B
+ sky130_fd_sc_hd__o21ai_1_290/B1 sky130_fd_sc_hd__nor2b_2_2/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_156 vccd1 vssd1 sky130_fd_sc_hd__and3_4_1/X sky130_fd_sc_hd__nor2_2_4/B
+ sky130_fd_sc_hd__buf_2_4/X sky130_fd_sc_hd__nor2_2_9/Y sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__o21ai_1_304/B1 sky130_fd_sc_hd__and2b_4_3/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_304 sky130_fd_sc_hd__fa_2_293/A sky130_fd_sc_hd__fa_2_303/B
+ sky130_fd_sc_hd__fa_2_304/A sky130_fd_sc_hd__fa_2_304/B sky130_fd_sc_hd__xor2_1_462/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_167 vccd1 vssd1 sky130_fd_sc_hd__and3_4_7/X sky130_fd_sc_hd__clkbuf_1_3/X
+ sky130_fd_sc_hd__or2_0_53/A sky130_fd_sc_hd__nor2_2_7/Y sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__o21ai_1_318/B1 sky130_fd_sc_hd__nor2b_2_1/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_315 sky130_fd_sc_hd__fa_2_300/B sky130_fd_sc_hd__fa_2_317/CIN
+ sky130_fd_sc_hd__fa_2_315/A sky130_fd_sc_hd__fa_2_315/B sky130_fd_sc_hd__fa_2_316/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_178 vccd1 vssd1 sky130_fd_sc_hd__and3_4_2/X sky130_fd_sc_hd__nor2_2_5/B
+ sky130_fd_sc_hd__nor2_2_4/B sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__buf_2_4/A
+ sky130_fd_sc_hd__o21ai_1_334/B1 sky130_fd_sc_hd__and2b_4_4/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_326 sky130_fd_sc_hd__fa_2_323/CIN sky130_fd_sc_hd__fa_2_333/A
+ sky130_fd_sc_hd__fa_2_326/A sky130_fd_sc_hd__fa_2_326/B sky130_fd_sc_hd__fa_2_330/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_189 vccd1 vssd1 sky130_fd_sc_hd__and3_4_2/X sky130_fd_sc_hd__buf_4_6/X
+ sky130_fd_sc_hd__and2_0_25/A sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__nor2_2_5/A
+ sky130_fd_sc_hd__o21ai_1_351/B1 sky130_fd_sc_hd__and2b_4_4/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_337 sky130_fd_sc_hd__fa_2_333/B sky130_fd_sc_hd__fa_2_341/CIN
+ sky130_fd_sc_hd__fa_2_337/A sky130_fd_sc_hd__fa_2_337/B sky130_fd_sc_hd__fa_2_337/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_348 sky130_fd_sc_hd__or2_1_6/A sky130_fd_sc_hd__nor2_2_23/B
+ sky130_fd_sc_hd__fa_2_348/A sky130_fd_sc_hd__fa_2_348/B sky130_fd_sc_hd__fa_2_348/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_359 sky130_fd_sc_hd__fa_2_355/B sky130_fd_sc_hd__fa_2_362/CIN
+ sky130_fd_sc_hd__fa_2_359/A sky130_fd_sc_hd__fa_2_359/B sky130_fd_sc_hd__fa_2_359/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_8_20 sky130_fd_sc_hd__clkinv_8_22/A sky130_fd_sc_hd__clkinv_8_20/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_31 sky130_fd_sc_hd__clkinv_8_31/Y sky130_fd_sc_hd__clkinv_8_89/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_42 sky130_fd_sc_hd__clkinv_8_43/A sky130_fd_sc_hd__clkinv_8_42/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_53 sky130_fd_sc_hd__clkinv_8_58/A sky130_fd_sc_hd__clkinv_8_53/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_64 sky130_fd_sc_hd__clkinv_8_65/A sky130_fd_sc_hd__clkinv_8_4/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_75 sky130_fd_sc_hd__clkinv_8_75/Y sky130_fd_sc_hd__clkinv_8_75/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_86 sky130_fd_sc_hd__dfxtp_1_9/CLK sky130_fd_sc_hd__clkinv_8_86/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_40 sky130_fd_sc_hd__inv_2_178/Y sky130_fd_sc_hd__buf_12_40/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_51 sky130_fd_sc_hd__inv_2_182/Y sky130_fd_sc_hd__buf_12_51/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_62 sky130_fd_sc_hd__inv_2_188/Y sky130_fd_sc_hd__buf_12_62/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_73 sky130_fd_sc_hd__buf_8_154/X sky130_fd_sc_hd__buf_12_73/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_84 sky130_fd_sc_hd__buf_8_56/X sky130_fd_sc_hd__buf_12_84/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_95 sky130_fd_sc_hd__buf_8_31/X sky130_fd_sc_hd__buf_12_95/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_2_2 vccd1 vssd1 sky130_fd_sc_hd__buf_2_2/X sky130_fd_sc_hd__buf_2_2/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_12_309 sky130_fd_sc_hd__buf_12_309/A sky130_fd_sc_hd__buf_12_309/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__inv_2_2 sky130_fd_sc_hd__inv_2_2/A sky130_fd_sc_hd__inv_2_2/Y vccd1
+ vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__clkinv_1_509 sky130_fd_sc_hd__nand2_1_488/A sky130_fd_sc_hd__o21a_1_3/A2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_12 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_12/Y
+ sky130_fd_sc_hd__nor2_1_12/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_23 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_23/Y
+ sky130_fd_sc_hd__nor2_1_23/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_34 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_34/Y
+ sky130_fd_sc_hd__nor2_1_34/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_45 sky130_fd_sc_hd__nor2_1_45/B sky130_fd_sc_hd__nor2_1_45/Y
+ sky130_fd_sc_hd__nor2_1_45/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_56 sky130_fd_sc_hd__and3_1_0/B sky130_fd_sc_hd__nor2_1_56/Y
+ sky130_fd_sc_hd__and3_1_0/C vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_67 sky130_fd_sc_hd__nor2_1_67/B sky130_fd_sc_hd__nor2_1_67/Y
+ sky130_fd_sc_hd__nor2_1_67/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_78 sky130_fd_sc_hd__nor2_1_81/Y sky130_fd_sc_hd__nor2_1_78/Y
+ sky130_fd_sc_hd__nor2_1_85/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_89 sky130_fd_sc_hd__nor2_1_95/Y sky130_fd_sc_hd__nor2_1_89/Y
+ sky130_fd_sc_hd__nor2_1_92/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_12_505 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_516 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_400 sky130_fd_sc_hd__nand2_1_400/Y sky130_fd_sc_hd__nand2_1_410/Y
+ sky130_fd_sc_hd__nand2_1_406/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_527 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_411 sky130_fd_sc_hd__nand2_1_411/Y sky130_fd_sc_hd__nand2_1_424/Y
+ sky130_fd_sc_hd__nand2_1_418/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_538 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_422 sky130_fd_sc_hd__nand2_1_422/Y sky130_fd_sc_hd__nor2_1_136/Y
+ sky130_fd_sc_hd__nand2_1_427/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_549 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_433 sky130_fd_sc_hd__nor2_1_132/B sky130_fd_sc_hd__nor2_1_143/Y
+ sky130_fd_sc_hd__nor2_1_105/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_444 sky130_fd_sc_hd__xnor2_1_110/A sky130_fd_sc_hd__nand2_1_445/Y
+ sky130_fd_sc_hd__nand2_1_444/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_455 sky130_fd_sc_hd__nand2_1_455/Y sky130_fd_sc_hd__nor2_1_153/Y
+ sky130_fd_sc_hd__nor2_1_156/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_466 sky130_fd_sc_hd__nand2_1_466/Y sky130_fd_sc_hd__or2_0_43/A
+ sky130_fd_sc_hd__or2_0_43/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_477 sky130_fd_sc_hd__xnor2_1_121/A sky130_fd_sc_hd__nand2_1_478/Y
+ sky130_fd_sc_hd__nand2_1_477/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_488 sky130_fd_sc_hd__xor2_1_421/A sky130_fd_sc_hd__o21a_1_3/B1
+ sky130_fd_sc_hd__nand2_1_488/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_499 sky130_fd_sc_hd__nand2_1_499/Y sky130_fd_sc_hd__nor2_2_32/Y
+ sky130_fd_sc_hd__or2_0_72/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_13 sky130_fd_sc_hd__nor2_1_167/B sky130_fd_sc_hd__nor2b_1_13/Y
+ sky130_fd_sc_hd__nor2b_1_13/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_24 sky130_fd_sc_hd__or2_0_84/A sky130_fd_sc_hd__fa_2_448/A
+ sky130_fd_sc_hd__nor2b_1_24/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_35 sky130_fd_sc_hd__fa_2_419/A sky130_fd_sc_hd__nor2b_1_35/Y
+ sky130_fd_sc_hd__buf_2_214/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1002 sky130_fd_sc_hd__clkinv_1_1003/A sky130_fd_sc_hd__inv_4_2/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_46 sky130_fd_sc_hd__mux2_2_42/X sky130_fd_sc_hd__fa_2_474/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1013 sky130_fd_sc_hd__clkinv_1_1013/Y sky130_fd_sc_hd__clkinv_1_1013/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_57 sky130_fd_sc_hd__or2_0_77/B sky130_fd_sc_hd__nor2b_1_57/Y
+ sky130_fd_sc_hd__buf_2_214/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1024 sky130_fd_sc_hd__buf_8_52/A sky130_fd_sc_hd__clkinv_2_37/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_68 sky130_fd_sc_hd__or2_0_80/A sky130_fd_sc_hd__fa_2_485/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1035 sky130_fd_sc_hd__inv_2_162/A sky130_fd_sc_hd__clkbuf_1_160/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_79 sky130_fd_sc_hd__buf_4_41/X sky130_fd_sc_hd__nor2b_1_79/Y
+ sky130_fd_sc_hd__mux2_4_5/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1046 sky130_fd_sc_hd__inv_2_179/A sky130_fd_sc_hd__clkbuf_1_195/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1504 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1057 sky130_fd_sc_hd__clkbuf_1_297/A sky130_fd_sc_hd__buf_8_74/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1515 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1068 sky130_fd_sc_hd__and2_0_401/B sky130_fd_sc_hd__nor2_1_267/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_9 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_9/B sky130_fd_sc_hd__xnor2_1_9/Y
+ sky130_fd_sc_hd__xnor2_1_9/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_1526 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1079 sky130_fd_sc_hd__and2_0_402/A sky130_fd_sc_hd__ha_2_53/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1537 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_240 sky130_fd_sc_hd__xor2_1_291/A sky130_fd_sc_hd__dfxtp_2_4/CLK
+ sky130_fd_sc_hd__and2_0_68/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1548 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_251 sky130_fd_sc_hd__xnor2_1_55/A sky130_fd_sc_hd__dfxtp_1_264/CLK
+ sky130_fd_sc_hd__and2_0_23/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1559 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_262 sky130_fd_sc_hd__xnor2_1_34/A sky130_fd_sc_hd__dfxtp_1_266/CLK
+ sky130_fd_sc_hd__and2_0_85/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_273 sky130_fd_sc_hd__fa_2_28/A sky130_fd_sc_hd__dfxtp_1_275/CLK
+ sky130_fd_sc_hd__and2_0_90/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_284 sky130_fd_sc_hd__dfxtp_1_284/Q sky130_fd_sc_hd__dfxtp_1_2/CLK
+ sky130_fd_sc_hd__and2_0_260/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_295 sky130_fd_sc_hd__dfxtp_1_295/Q sky130_fd_sc_hd__clkinv_8_6/Y
+ sky130_fd_sc_hd__and2_0_271/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__mux2_4_5 sky130_fd_sc_hd__mux2_4_5/X sky130_fd_sc_hd__mux2_8_1/S
+ sky130_fd_sc_hd__buf_2_69/X sky130_fd_sc_hd__mux2_4_5/A1 vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__mux2_4
Xsky130_fd_sc_hd__o22ai_1_4 sky130_fd_sc_hd__o22ai_1_4/A2 sky130_fd_sc_hd__o22ai_1_4/B1
+ sky130_fd_sc_hd__o22ai_1_4/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__o22ai_1_9/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_101 sky130_fd_sc_hd__fa_2_98/B sky130_fd_sc_hd__fa_2_103/CIN
+ sky130_fd_sc_hd__fa_2_101/A sky130_fd_sc_hd__fa_2_101/B sky130_fd_sc_hd__fa_2_99/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_112 sky130_fd_sc_hd__fa_2_107/A sky130_fd_sc_hd__fa_2_111/B
+ sky130_fd_sc_hd__fa_2_112/A sky130_fd_sc_hd__fa_2_112/B sky130_fd_sc_hd__fa_2_112/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_123 sky130_fd_sc_hd__nor2_1_83/A sky130_fd_sc_hd__nor2_1_86/B
+ sky130_fd_sc_hd__fa_2_123/A sky130_fd_sc_hd__fa_2_123/B sky130_fd_sc_hd__fa_2_123/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_134 sky130_fd_sc_hd__nor2_1_94/A sky130_fd_sc_hd__nor2_1_97/B
+ sky130_fd_sc_hd__fa_2_134/A sky130_fd_sc_hd__fa_2_134/B sky130_fd_sc_hd__xor2_1_188/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_145 sky130_fd_sc_hd__xor3_1_12/A sky130_fd_sc_hd__fa_2_146/B
+ sky130_fd_sc_hd__fa_2_145/A sky130_fd_sc_hd__fa_2_145/B sky130_fd_sc_hd__xor2_1_231/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_156 sky130_fd_sc_hd__fa_2_147/A sky130_fd_sc_hd__fa_2_157/B
+ sky130_fd_sc_hd__fa_2_156/A sky130_fd_sc_hd__fa_2_156/B sky130_fd_sc_hd__fa_2_156/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_167 sky130_fd_sc_hd__fa_2_159/B sky130_fd_sc_hd__fa_2_167/SUM
+ sky130_fd_sc_hd__fa_2_167/A sky130_fd_sc_hd__fa_2_167/B sky130_fd_sc_hd__fa_2_168/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and3_4_6 sky130_fd_sc_hd__and3_4_6/A sky130_fd_sc_hd__and3_4_6/B
+ sky130_fd_sc_hd__and3_4_6/C sky130_fd_sc_hd__and3_4_6/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__fa_2_178 sky130_fd_sc_hd__fa_2_176/CIN sky130_fd_sc_hd__fa_2_184/B
+ sky130_fd_sc_hd__fa_2_178/A sky130_fd_sc_hd__fa_2_178/B sky130_fd_sc_hd__xor2_1_274/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_189 sky130_fd_sc_hd__fa_2_185/B sky130_fd_sc_hd__fa_2_193/CIN
+ sky130_fd_sc_hd__fa_2_189/A sky130_fd_sc_hd__fa_2_189/B sky130_fd_sc_hd__fa_2_189/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o22ai_1_11 sky130_fd_sc_hd__o22ai_1_52/B1 sky130_fd_sc_hd__o22ai_1_11/B1
+ sky130_fd_sc_hd__o22ai_1_11/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__inv_4_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_22 sky130_fd_sc_hd__o22ai_1_41/B1 sky130_fd_sc_hd__o22ai_1_22/B1
+ sky130_fd_sc_hd__o22ai_1_22/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__inv_4_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_140 vccd1 vssd1 sky130_fd_sc_hd__buf_2_140/X sky130_fd_sc_hd__buf_2_140/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_33 sky130_fd_sc_hd__nor2_1_32/A sky130_fd_sc_hd__o22ai_1_33/B1
+ sky130_fd_sc_hd__o22ai_1_33/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_151 vccd1 vssd1 sky130_fd_sc_hd__buf_2_151/X sky130_fd_sc_hd__buf_2_151/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_44 sky130_fd_sc_hd__nor2_1_23/A sky130_fd_sc_hd__o22ai_1_44/B1
+ sky130_fd_sc_hd__o22ai_1_44/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_162 vccd1 vssd1 sky130_fd_sc_hd__buf_2_162/X sky130_fd_sc_hd__buf_6_19/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_55 sky130_fd_sc_hd__nor2_1_12/A sky130_fd_sc_hd__o22ai_1_8/A2
+ sky130_fd_sc_hd__o22ai_1_55/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_173 vccd1 vssd1 sky130_fd_sc_hd__nor2_4_0/B la_data_out[34]
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_66 sky130_fd_sc_hd__xnor2_1_258/Y sky130_fd_sc_hd__xnor2_1_219/Y
+ sky130_fd_sc_hd__fa_2_426/A sky130_fd_sc_hd__nor2b_1_19/A sky130_fd_sc_hd__o22ai_1_66/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_184 vccd1 vssd1 sky130_fd_sc_hd__buf_2_184/X sky130_fd_sc_hd__buf_2_184/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_77 sky130_fd_sc_hd__xnor2_2_4/Y sky130_fd_sc_hd__xnor2_1_230/Y
+ sky130_fd_sc_hd__o22ai_1_77/Y sky130_fd_sc_hd__xnor2_1_228/Y sky130_fd_sc_hd__o22ai_1_96/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_195 vccd1 vssd1 la_data_out[82] sky130_fd_sc_hd__xnor2_2_5/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_88 sky130_fd_sc_hd__xnor2_1_236/Y sky130_fd_sc_hd__xnor2_1_235/Y
+ sky130_fd_sc_hd__or2_0_97/B sky130_fd_sc_hd__inv_2_65/Y sky130_fd_sc_hd__o22ai_1_99/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_99 sky130_fd_sc_hd__xnor2_1_248/Y sky130_fd_sc_hd__xnor2_1_247/Y
+ sky130_fd_sc_hd__ha_2_15/B sky130_fd_sc_hd__inv_2_65/Y sky130_fd_sc_hd__o22ai_1_99/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_4_13 vccd1 vssd1 sky130_fd_sc_hd__buf_4_13/X sky130_fd_sc_hd__buf_4_13/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_24 vccd1 vssd1 sky130_fd_sc_hd__buf_4_24/X sky130_fd_sc_hd__buf_4_24/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_35 vccd1 vssd1 sky130_fd_sc_hd__buf_4_35/X sky130_fd_sc_hd__buf_8_21/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_12_106 sky130_fd_sc_hd__buf_8_33/X sky130_fd_sc_hd__buf_12_339/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_117 sky130_fd_sc_hd__buf_8_36/X sky130_fd_sc_hd__buf_12_341/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_40 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_40/X sky130_fd_sc_hd__buf_2_184/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_128 sky130_fd_sc_hd__buf_8_46/X sky130_fd_sc_hd__buf_12_409/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_51 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_51/X sky130_fd_sc_hd__clkbuf_1_52/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_139 sky130_fd_sc_hd__buf_8_124/X sky130_fd_sc_hd__buf_12_139/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_62 vssd1 vccd1 sky130_fd_sc_hd__buf_8_42/A sky130_fd_sc_hd__buf_2_61/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_73 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_10/A1 sky130_fd_sc_hd__clkbuf_1_73/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_84 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_32/A1 sky130_fd_sc_hd__clkbuf_1_84/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_95 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_7/A1 sky130_fd_sc_hd__clkbuf_1_95/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_4_9 sky130_fd_sc_hd__clkbuf_4_9/X sky130_fd_sc_hd__clkbuf_4_9/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_1_306 sky130_fd_sc_hd__nand3_1_3/A sky130_fd_sc_hd__ha_2_5/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_317 sky130_fd_sc_hd__a21oi_1_39/A1 sky130_fd_sc_hd__nor2_1_49/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_328 sky130_fd_sc_hd__o21ai_1_219/A2 sky130_fd_sc_hd__xnor2_1_13/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_339 sky130_fd_sc_hd__nand2_1_199/A sky130_fd_sc_hd__nor2_1_60/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__or2_0_20 sky130_fd_sc_hd__or2_0_66/A sky130_fd_sc_hd__or2_0_20/X
+ sky130_fd_sc_hd__buf_4_5/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_31 sky130_fd_sc_hd__or2_0_9/A sky130_fd_sc_hd__or2_0_31/X
+ sky130_fd_sc_hd__or2_0_4/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_42 sky130_fd_sc_hd__or2_0_61/A sky130_fd_sc_hd__or2_0_42/X
+ sky130_fd_sc_hd__or2_0_42/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_53 sky130_fd_sc_hd__or2_0_53/A sky130_fd_sc_hd__or2_0_53/X
+ sky130_fd_sc_hd__inv_6_0/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_64 sky130_fd_sc_hd__buf_4_2/X sky130_fd_sc_hd__or2_0_64/X
+ sky130_fd_sc_hd__buf_4_4/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_75 sky130_fd_sc_hd__or2_0_75/A sky130_fd_sc_hd__or2_0_75/X
+ sky130_fd_sc_hd__or2_0_75/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__clkinv_4_9 sky130_fd_sc_hd__clkinv_4_9/A sky130_fd_sc_hd__clkinv_4_9/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__or2_0_86 sky130_fd_sc_hd__or2_0_86/A sky130_fd_sc_hd__or2_0_86/X
+ sky130_fd_sc_hd__or2_0_86/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_97 sky130_fd_sc_hd__or2_0_97/A sky130_fd_sc_hd__or2_0_97/X
+ sky130_fd_sc_hd__or2_0_97/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__clkinv_4_100 sky130_fd_sc_hd__clkinv_4_99/Y sky130_fd_sc_hd__clkinv_8_55/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_12_640 sky130_fd_sc_hd__buf_12_640/A sky130_fd_sc_hd__buf_12_640/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_4_111 sky130_fd_sc_hd__clkinv_4_114/A sky130_fd_sc_hd__clkinv_8_66/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_12_651 sky130_fd_sc_hd__buf_12_651/A sky130_fd_sc_hd__buf_12_651/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_4_122 sky130_fd_sc_hd__clkinv_8_86/A sky130_fd_sc_hd__dfxtp_1_1/CLK
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_12_662 sky130_fd_sc_hd__buf_12_662/A sky130_fd_sc_hd__buf_12_662/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_673 sky130_fd_sc_hd__buf_12_673/A sky130_fd_sc_hd__buf_12_673/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_302 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_313 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_324 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_335 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_346 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_230 sky130_fd_sc_hd__xnor2_1_30/A sky130_fd_sc_hd__nand2_1_231/Y
+ sky130_fd_sc_hd__or2_0_18/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_357 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_241 sky130_fd_sc_hd__nor2_1_74/A sky130_fd_sc_hd__nor2_1_75/Y
+ sky130_fd_sc_hd__nor2_1_78/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_368 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_840 sky130_fd_sc_hd__inv_2_74/A la_data_out[50] vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_252 sky130_fd_sc_hd__xnor2_1_39/A sky130_fd_sc_hd__nand2_1_253/Y
+ sky130_fd_sc_hd__nand2_1_252/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_379 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_851 sky130_fd_sc_hd__clkinv_1_851/Y sky130_fd_sc_hd__clkinv_8_8/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_263 sky130_fd_sc_hd__xnor2_1_42/A sky130_fd_sc_hd__nand2_1_264/Y
+ sky130_fd_sc_hd__nand2_1_263/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_862 sky130_fd_sc_hd__clkinv_1_862/Y sky130_fd_sc_hd__inv_2_196/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_274 sky130_fd_sc_hd__nand2_1_274/Y sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__buf_6_1/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_873 sky130_fd_sc_hd__clkinv_1_873/Y sky130_fd_sc_hd__clkinv_4_84/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_285 sky130_fd_sc_hd__xor2_1_187/A sky130_fd_sc_hd__nand2_1_286/Y
+ sky130_fd_sc_hd__nand2_1_285/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_884 sky130_fd_sc_hd__clkinv_1_884/Y sky130_fd_sc_hd__clkinv_4_87/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_296 sky130_fd_sc_hd__xnor2_1_2/B sky130_fd_sc_hd__nand2_1_297/Y
+ sky130_fd_sc_hd__nand2_1_296/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_895 sky130_fd_sc_hd__clkinv_1_895/Y sky130_fd_sc_hd__inv_2_199/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1301 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_2_1 vccd1 vssd1 sky130_fd_sc_hd__xor2_2_1/X sky130_fd_sc_hd__xor2_2_1/B
+ sky130_fd_sc_hd__xor2_2_1/A vssd1 vccd1 sky130_fd_sc_hd__xor2_2
Xsky130_fd_sc_hd__conb_1_40 sky130_fd_sc_hd__conb_1_40/LO sky130_fd_sc_hd__conb_1_40/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1312 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_51 sky130_fd_sc_hd__conb_1_51/LO sky130_fd_sc_hd__conb_1_51/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1323 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_62 sky130_fd_sc_hd__conb_1_62/LO sky130_fd_sc_hd__conb_1_62/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1334 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_73 sky130_fd_sc_hd__conb_1_73/LO sky130_fd_sc_hd__conb_1_73/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1345 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_84 sky130_fd_sc_hd__conb_1_84/LO sky130_fd_sc_hd__conb_1_84/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1356 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_95 sky130_fd_sc_hd__conb_1_95/LO sky130_fd_sc_hd__conb_1_95/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1367 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1378 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_809 vssd1 vccd1 sky130_fd_sc_hd__buf_2_13/X sky130_fd_sc_hd__nand2b_1_16/Y
+ sky130_fd_sc_hd__o21ai_1_809/B1 sky130_fd_sc_hd__xor2_1_584/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1389 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__mux2_2_2 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_2/A1 sky130_fd_sc_hd__buf_4_18/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__or2_1_10/A vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__decap_12_880 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_891 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_603 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__xor2_1_603/X
+ sky130_fd_sc_hd__xor2_1_603/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_614 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__xor2_1_614/X
+ sky130_fd_sc_hd__xor2_1_614/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_625 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__xor2_1_625/X
+ sky130_fd_sc_hd__xor2_1_625/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_636 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__xor2_1_636/X
+ sky130_fd_sc_hd__xor2_1_636/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_647 sky130_fd_sc_hd__xor2_1_647/B sky130_fd_sc_hd__xor2_1_647/X
+ sky130_fd_sc_hd__xor2_1_647/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_658 sky130_fd_sc_hd__xor2_1_658/B sky130_fd_sc_hd__a22o_1_8/B1
+ sky130_fd_sc_hd__xor2_1_658/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_669 sky130_fd_sc_hd__xnor2_2_5/A sky130_fd_sc_hd__xor2_1_669/X
+ sky130_fd_sc_hd__buf_2_207/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a211o_1_16 vssd1 vccd1 sky130_fd_sc_hd__fa_2_246/A sky130_fd_sc_hd__dfxtp_1_79/Q
+ sky130_fd_sc_hd__nor2_1_20/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_16/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__a211o_1_27 vssd1 vccd1 sky130_fd_sc_hd__fa_2_170/B sky130_fd_sc_hd__dfxtp_1_90/Q
+ sky130_fd_sc_hd__nor2_1_31/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_27/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__clkinv_1_103 io_oeb[36] sky130_fd_sc_hd__conb_1_39/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_114 io_oeb[25] sky130_fd_sc_hd__conb_1_28/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_125 io_oeb[14] sky130_fd_sc_hd__conb_1_17/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_136 io_oeb[3] sky130_fd_sc_hd__conb_1_6/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_147 sky130_fd_sc_hd__and2_0_249/A sky130_fd_sc_hd__a222oi_1_48/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_158 sky130_fd_sc_hd__nor2_1_31/A sky130_fd_sc_hd__dfxtp_1_154/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_169 sky130_fd_sc_hd__o22ai_1_38/B1 sky130_fd_sc_hd__dfxtp_1_183/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_16 sky130_fd_sc_hd__inv_2_66/Y sky130_fd_sc_hd__xor2_1_662/X
+ sky130_fd_sc_hd__a22o_1_16/X sky130_fd_sc_hd__nor2_1_233/Y sky130_fd_sc_hd__xor2_1_654/X
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_27 sky130_fd_sc_hd__buf_2_63/A sky130_fd_sc_hd__buf_2_102/X
+ sky130_fd_sc_hd__a22o_1_27/X sky130_fd_sc_hd__a22o_1_27/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_38 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__buf_2_113/X
+ sky130_fd_sc_hd__a22o_1_38/X sky130_fd_sc_hd__a22o_1_38/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_49 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__buf_2_123/X
+ sky130_fd_sc_hd__a22o_1_49/X sky130_fd_sc_hd__a22o_1_49/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__o21ai_1_3 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_3/A2 sky130_fd_sc_hd__nor2_4_4/B
+ sky130_fd_sc_hd__o21ai_1_3/B1 sky130_fd_sc_hd__fa_2_19/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2_1_230 sky130_fd_sc_hd__mux2_2_49/X sky130_fd_sc_hd__nor2_1_230/Y
+ la_data_out[72] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_241 sky130_fd_sc_hd__a22o_1_8/A2 sky130_fd_sc_hd__nor2_1_241/Y
+ sky130_fd_sc_hd__nor2_1_241/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_252 sky130_fd_sc_hd__nor2_1_252/B sky130_fd_sc_hd__nor2_1_252/Y
+ sky130_fd_sc_hd__nor2_1_252/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_2_6 sky130_fd_sc_hd__clkinv_2_7/A sky130_fd_sc_hd__clkinv_4_3/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__nor2_1_263 sky130_fd_sc_hd__nor2_1_263/B sky130_fd_sc_hd__nor2_1_263/Y
+ sky130_fd_sc_hd__nor2_1_263/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_274 sky130_fd_sc_hd__ha_2_46/B sky130_fd_sc_hd__nor2_1_274/Y
+ sky130_fd_sc_hd__ha_2_46/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_470 sky130_fd_sc_hd__buf_12_470/A sky130_fd_sc_hd__buf_12_539/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_481 sky130_fd_sc_hd__buf_12_481/A sky130_fd_sc_hd__buf_12_519/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_110 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_492 sky130_fd_sc_hd__buf_12_492/A sky130_fd_sc_hd__buf_12_632/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_121 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_132 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_143 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_154 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_165 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_200 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_200/B sky130_fd_sc_hd__and2_0_253/A
+ sky130_fd_sc_hd__xnor2_1_200/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_176 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_211 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_211/B sky130_fd_sc_hd__a22o_1_9/B1
+ sky130_fd_sc_hd__xnor2_1_211/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_187 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_17 sky130_fd_sc_hd__nand2_1_17/Y sky130_fd_sc_hd__nand2_1_17/B
+ sky130_fd_sc_hd__nand2_1_17/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_222 vssd1 vccd1 la_data_out[85] sky130_fd_sc_hd__xnor2_1_222/Y
+ la_data_out[68] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_198 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_670 sky130_fd_sc_hd__xnor2_1_208/B sky130_fd_sc_hd__a21oi_1_156/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_28 sky130_fd_sc_hd__nand2_1_28/Y sky130_fd_sc_hd__nand2_1_7/B
+ sky130_fd_sc_hd__or2_0_79/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_233 vssd1 vccd1 la_data_out[77] sky130_fd_sc_hd__xnor2_1_233/Y
+ sky130_fd_sc_hd__mux2_4_2/X vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_681 sky130_fd_sc_hd__clkinv_1_681/Y sky130_fd_sc_hd__nand2_1_773/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_39 sky130_fd_sc_hd__nand2_1_39/Y sky130_fd_sc_hd__nand2_1_7/B
+ la_data_out[71] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_244 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_5/B sky130_fd_sc_hd__xnor2_1_244/Y
+ la_data_out[68] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_692 sky130_fd_sc_hd__nand2_1_767/A sky130_fd_sc_hd__nor2_1_248/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_255 vssd1 vccd1 la_data_out[85] sky130_fd_sc_hd__xnor2_1_255/Y
+ sky130_fd_sc_hd__or2_0_82/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_266 vssd1 vccd1 sky130_fd_sc_hd__buf_2_207/X sky130_fd_sc_hd__xnor2_1_266/Y
+ sky130_fd_sc_hd__or2_1_10/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_277 vssd1 vccd1 sky130_fd_sc_hd__or2_0_84/A sky130_fd_sc_hd__xnor2_1_277/Y
+ sky130_fd_sc_hd__or2_0_77/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_288 vssd1 vccd1 la_data_out[77] sky130_fd_sc_hd__xnor2_1_288/Y
+ sky130_fd_sc_hd__mux2_2_27/X vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_299 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_299/B sky130_fd_sc_hd__xnor2_1_299/Y
+ sky130_fd_sc_hd__xnor2_1_299/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_1120 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1131 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1142 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1153 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1164 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1175 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_606 vssd1 vccd1 sky130_fd_sc_hd__buf_2_9/X sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_606/B1 sky130_fd_sc_hd__xor2_1_398/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1186 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_617 vssd1 vccd1 sky130_fd_sc_hd__buf_2_11/X sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_617/B1 sky130_fd_sc_hd__xor2_1_410/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1197 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_628 vssd1 vccd1 sky130_fd_sc_hd__nand2_2_12/Y sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__a22oi_1_211/Y sky130_fd_sc_hd__xor2_1_422/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_639 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_742/A2 sky130_fd_sc_hd__nand2b_2_6/Y
+ sky130_fd_sc_hd__o21ai_1_639/B1 sky130_fd_sc_hd__xor2_1_427/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fah_1_4 sky130_fd_sc_hd__fa_2_245/B sky130_fd_sc_hd__fah_1_4/B sky130_fd_sc_hd__fah_1_4/A
+ sky130_fd_sc_hd__fah_1_3/CI sky130_fd_sc_hd__fah_1_4/CI vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__fah_1
Xsky130_fd_sc_hd__sdlclkp_2_11 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_8_5/Y
+ sky130_fd_sc_hd__dfxtp_2_4/CLK sky130_fd_sc_hd__o21ai_2_3/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__a222oi_1_90 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__or2_0_61/A
+ sky130_fd_sc_hd__or2_0_42/B sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__or2_0_58/B
+ sky130_fd_sc_hd__a222oi_1_90/Y sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__xor2_1_400 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__xor2_1_400/X
+ sky130_fd_sc_hd__xor2_1_400/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_70 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_70/B sky130_fd_sc_hd__xnor2_1_70/Y
+ sky130_fd_sc_hd__xnor2_1_70/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_411 sky130_fd_sc_hd__xor2_1_411/B sky130_fd_sc_hd__xor2_1_411/X
+ sky130_fd_sc_hd__xor2_1_411/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_81 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_291/A sky130_fd_sc_hd__nor2b_1_9/A
+ sky130_fd_sc_hd__xnor2_1_84/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_422 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__xor2_1_422/X
+ sky130_fd_sc_hd__xor2_1_422/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_92 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_92/B sky130_fd_sc_hd__inv_2_37/A
+ sky130_fd_sc_hd__xnor2_1_92/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_433 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__xor3_1_27/A
+ sky130_fd_sc_hd__xor2_1_433/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_444 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__xor2_1_444/X
+ sky130_fd_sc_hd__xor2_1_444/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_455 sky130_fd_sc_hd__fah_1_14/A sky130_fd_sc_hd__xor2_1_455/X
+ sky130_fd_sc_hd__xor2_1_455/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_466 sky130_fd_sc_hd__xor2_1_548/B sky130_fd_sc_hd__xor2_1_466/X
+ sky130_fd_sc_hd__xor2_1_466/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_477 sky130_fd_sc_hd__fah_1_14/A sky130_fd_sc_hd__xor2_1_477/X
+ sky130_fd_sc_hd__xor2_1_477/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_488 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__fa_2_318/B
+ sky130_fd_sc_hd__xor2_1_488/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_499 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__fa_2_336/B
+ sky130_fd_sc_hd__xor2_1_499/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a222oi_1_508 vccd1 vssd1 sky130_fd_sc_hd__and3_4_21/X sky130_fd_sc_hd__buf_2_27/X
+ sky130_fd_sc_hd__buf_2_15/X sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__buf_2_4/A
+ sky130_fd_sc_hd__o21ai_1_637/B1 sky130_fd_sc_hd__and2b_4_12/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_519 vccd1 vssd1 sky130_fd_sc_hd__and3_4_21/X sky130_fd_sc_hd__buf_2_30/X
+ sky130_fd_sc_hd__buf_2_26/X sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__buf_4_0/X
+ sky130_fd_sc_hd__o21ai_1_819/B1 sky130_fd_sc_hd__and2b_4_12/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nor2b_1_108 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_108/Y
+ sky130_fd_sc_hd__nor2b_1_108/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_119 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_119/Y
+ sky130_fd_sc_hd__nor2b_1_119/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__decap_12_0 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_9 vccd1 vssd1 sky130_fd_sc_hd__buf_6_9/X sky130_fd_sc_hd__buf_6_9/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__clkinv_2_11 sky130_fd_sc_hd__clkinv_2_12/A sky130_fd_sc_hd__clkinv_2_11/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_22 sky130_fd_sc_hd__inv_2_120/A sky130_fd_sc_hd__o21ai_1_925/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_33 sky130_fd_sc_hd__clkinv_2_33/Y sky130_fd_sc_hd__clkinv_2_33/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_44 sky130_fd_sc_hd__inv_2_172/A sky130_fd_sc_hd__buf_8_72/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__and2_0_402 vccd1 vssd1 sky130_fd_sc_hd__nor3_1_3/B la_data_out[47]
+ sky130_fd_sc_hd__and2_0_402/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_2_55 la_data_out[91] sky130_fd_sc_hd__clkinv_4_93/Y vccd1
+ vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__or2_1_4 sky130_fd_sc_hd__or2_1_4/A sky130_fd_sc_hd__or2_1_4/X sky130_fd_sc_hd__or2_1_4/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_1
Xsky130_fd_sc_hd__sdlclkp_4_7 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_4_3/Y
+ sky130_fd_sc_hd__dfxtp_1_85/CLK sky130_fd_sc_hd__o21ai_2_0/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__a22oi_1_170 sky130_fd_sc_hd__nand2_1_127/A sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xor2_1_176/X sky130_fd_sc_hd__a22oi_1_170/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_181 sky130_fd_sc_hd__xor2_1_411/X sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xor2_1_199/X sky130_fd_sc_hd__a22oi_1_181/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_192 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__nor2b_1_3/Y sky130_fd_sc_hd__nor2_1_56/Y sky130_fd_sc_hd__a22oi_1_192/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22o_4_1 sky130_fd_sc_hd__nand2_1_8/B sky130_fd_sc_hd__mux2_2_35/X
+ sky130_fd_sc_hd__or2_0_60/A sky130_fd_sc_hd__mux2_2_15/X sky130_fd_sc_hd__nand2_1_7/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_4
Xsky130_fd_sc_hd__o21ai_1_403 vssd1 vccd1 sky130_fd_sc_hd__buf_2_8/X sky130_fd_sc_hd__nand2b_1_12/Y
+ sky130_fd_sc_hd__o21ai_1_403/B1 sky130_fd_sc_hd__xor2_1_215/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_414 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_111/Y sky130_fd_sc_hd__nor2_1_107/A
+ sky130_fd_sc_hd__nor2_1_106/Y sky130_fd_sc_hd__o21ai_1_414/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_425 vssd1 vccd1 sky130_fd_sc_hd__buf_2_10/X sky130_fd_sc_hd__nand2b_1_11/Y
+ sky130_fd_sc_hd__o21ai_1_425/B1 sky130_fd_sc_hd__xor2_1_232/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_436 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_444/A2 sky130_fd_sc_hd__nor2_1_112/A
+ sky130_fd_sc_hd__nor2_1_111/Y sky130_fd_sc_hd__o21ai_1_436/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_447 vssd1 vccd1 sky130_fd_sc_hd__inv_2_28/Y sky130_fd_sc_hd__nand2b_1_12/Y
+ sky130_fd_sc_hd__o21ai_1_447/B1 sky130_fd_sc_hd__xor2_1_250/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_458 vssd1 vccd1 sky130_fd_sc_hd__buf_2_10/X sky130_fd_sc_hd__nand2b_1_12/Y
+ sky130_fd_sc_hd__o21ai_1_458/B1 sky130_fd_sc_hd__xor2_1_260/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_469 vssd1 vccd1 sky130_fd_sc_hd__inv_2_29/Y sky130_fd_sc_hd__nand2b_1_13/Y
+ sky130_fd_sc_hd__o21ai_1_469/B1 sky130_fd_sc_hd__xor2_1_272/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2_4_12 sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__nor2_4_12/A
+ sky130_fd_sc_hd__nor2_4_12/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__nand2_1_807 sky130_fd_sc_hd__nand2_1_807/Y sky130_fd_sc_hd__or2_0_103/A
+ sky130_fd_sc_hd__or2_0_103/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_818 sky130_fd_sc_hd__xnor2_1_297/A sky130_fd_sc_hd__nand2_1_819/Y
+ sky130_fd_sc_hd__or2_0_106/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_829 sky130_fd_sc_hd__nand2_1_829/Y sky130_fd_sc_hd__nor2_1_263/A
+ sky130_fd_sc_hd__nor2_1_263/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_230 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__fa_2_144/A
+ sky130_fd_sc_hd__xor2_1_230/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__o21ai_1_18 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_15/B1 sky130_fd_sc_hd__inv_2_53/A
+ sky130_fd_sc_hd__o21ai_1_18/B1 sky130_fd_sc_hd__fa_2_110/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_241 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__fa_2_153/B
+ sky130_fd_sc_hd__xor2_1_241/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__o21ai_1_29 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_4/B1 sky130_fd_sc_hd__nor2_4_4/B
+ sky130_fd_sc_hd__o21ai_1_29/B1 sky130_fd_sc_hd__fa_2_140/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_252 sky130_fd_sc_hd__xor2_1_383/B sky130_fd_sc_hd__fa_2_163/A
+ sky130_fd_sc_hd__xor2_1_252/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_263 sky130_fd_sc_hd__xor2_1_362/B sky130_fd_sc_hd__fa_2_171/A
+ sky130_fd_sc_hd__xor2_1_263/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_274 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__xor2_1_274/X
+ sky130_fd_sc_hd__xor2_1_274/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_285 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__fa_2_192/B
+ sky130_fd_sc_hd__xor2_1_285/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_296 sky130_fd_sc_hd__xor2_1_296/B sky130_fd_sc_hd__xor2_1_296/X
+ sky130_fd_sc_hd__xor2_1_296/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_201 vssd1 vccd1 sky130_fd_sc_hd__buf_12_31/A la_data_out[42]
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_212 vssd1 vccd1 sky130_fd_sc_hd__buf_8_60/A sky130_fd_sc_hd__buf_8_118/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_223 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4_27/A sky130_fd_sc_hd__nand2_2_7/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_234 vssd1 vccd1 sky130_fd_sc_hd__buf_12_46/A sky130_fd_sc_hd__inv_2_160/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_305 vccd1 vssd1 sky130_fd_sc_hd__and3_4_11/X sky130_fd_sc_hd__and2_0_49/A
+ sky130_fd_sc_hd__and2_0_45/A sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__and2_0_87/A
+ sky130_fd_sc_hd__o21ai_1_520/B1 sky130_fd_sc_hd__and2b_4_8/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_245 vssd1 vccd1 sky130_fd_sc_hd__buf_8_127/A sky130_fd_sc_hd__clkbuf_1_286/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_316 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__and2_0_45/A
+ sky130_fd_sc_hd__and2_0_87/A sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__o21ai_1_532/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_256 vssd1 vccd1 sky130_fd_sc_hd__buf_8_145/A sky130_fd_sc_hd__buf_8_44/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_2_3 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__clkinv_4_6/Y
+ sky130_fd_sc_hd__dfxtp_2_3/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_2
Xsky130_fd_sc_hd__a222oi_1_327 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__and2_0_49/A
+ sky130_fd_sc_hd__and2_0_45/A sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__and2_0_87/A
+ sky130_fd_sc_hd__o21ai_1_547/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_267 vssd1 vccd1 sky130_fd_sc_hd__buf_8_156/A sky130_fd_sc_hd__clkbuf_4_29/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_338 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__and2_0_45/A
+ sky130_fd_sc_hd__and2_0_87/A sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__o21ai_1_560/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_278 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_278/X sky130_fd_sc_hd__clkinv_1_902/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_349 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__buf_2_31/X
+ sky130_fd_sc_hd__buf_2_19/X sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__o21ai_1_577/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_289 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_290/A sky130_fd_sc_hd__buf_8_72/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_2_90 vccd1 vssd1 sky130_fd_sc_hd__buf_2_90/X sky130_fd_sc_hd__buf_2_90/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_4_6 vccd1 vssd1 sky130_fd_sc_hd__buf_4_6/X sky130_fd_sc_hd__buf_6_2/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__and2_0_210 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_84/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_74/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_221 vccd1 vssd1 sky130_fd_sc_hd__and2_0_221/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_221/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_232 vccd1 vssd1 sky130_fd_sc_hd__and2_0_232/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__o21ai_1_57/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_243 vccd1 vssd1 sky130_fd_sc_hd__and2_0_243/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__o21ai_1_48/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_254 vccd1 vssd1 sky130_fd_sc_hd__and2_0_254/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__xor2_1_651/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_265 vccd1 vssd1 sky130_fd_sc_hd__and2_0_265/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__and2_0_265/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_276 vccd1 vssd1 sky130_fd_sc_hd__and2_0_276/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__xor2_1_640/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__a21oi_2_17 sky130_fd_sc_hd__a21oi_2_17/B1 sky130_fd_sc_hd__or2_1_4/X
+ sky130_fd_sc_hd__o21ai_2_14/Y sky130_fd_sc_hd__xor2_1_526/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_2
Xsky130_fd_sc_hd__and2_0_287 vccd1 vssd1 sky130_fd_sc_hd__and2_0_287/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_8/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_298 vccd1 vssd1 sky130_fd_sc_hd__and2_0_298/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_19/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__sdlclkp_2_4 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_8_3/Y
+ sky130_fd_sc_hd__dfxtp_1_118/CLK sky130_fd_sc_hd__clkbuf_1_11/X vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__inv_4_6 sky130_fd_sc_hd__inv_4_6/Y sky130_fd_sc_hd__inv_4_6/A vccd1
+ vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__o21ai_1_200 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_2/X sky130_fd_sc_hd__nand2_1_175/Y
+ sky130_fd_sc_hd__a21oi_1_40/Y sky130_fd_sc_hd__xnor2_1_9/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_211 vssd1 vccd1 sky130_fd_sc_hd__buf_2_5/X sky130_fd_sc_hd__nand2b_1_5/Y
+ sky130_fd_sc_hd__a222oi_1_83/Y sky130_fd_sc_hd__xor2_1_36/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_222 vssd1 vccd1 sky130_fd_sc_hd__inv_2_24/Y sky130_fd_sc_hd__nand2b_2_0/Y
+ sky130_fd_sc_hd__a222oi_1_91/Y sky130_fd_sc_hd__xor2_1_46/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_40 la_data_out[61] sky130_fd_sc_hd__dfxtp_1_476/Q vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_233 vssd1 vccd1 sky130_fd_sc_hd__buf_2_2/X sky130_fd_sc_hd__nand2b_1_4/Y
+ sky130_fd_sc_hd__o21ai_1_233/B1 sky130_fd_sc_hd__xor2_1_58/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_51 la_data_out[81] sky130_fd_sc_hd__xnor2_2_5/B vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_244 vssd1 vccd1 sky130_fd_sc_hd__buf_2_5/X sky130_fd_sc_hd__nand2b_1_6/Y
+ sky130_fd_sc_hd__o21ai_1_244/B1 sky130_fd_sc_hd__xor2_1_67/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_255 vssd1 vccd1 sky130_fd_sc_hd__inv_2_26/Y sky130_fd_sc_hd__nand2b_1_4/Y
+ sky130_fd_sc_hd__nand2_1_154/Y sky130_fd_sc_hd__xor2_1_77/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_266 vssd1 vccd1 sky130_fd_sc_hd__inv_2_13/Y sky130_fd_sc_hd__nand2b_2_0/Y
+ sky130_fd_sc_hd__o21ai_1_266/B1 sky130_fd_sc_hd__xor2_1_88/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_277 vssd1 vccd1 sky130_fd_sc_hd__inv_2_22/Y sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__o21ai_1_277/B1 sky130_fd_sc_hd__xor2_1_98/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_288 vssd1 vccd1 sky130_fd_sc_hd__inv_2_24/Y sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__o21ai_1_288/B1 sky130_fd_sc_hd__xor2_1_109/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_299 vssd1 vccd1 sky130_fd_sc_hd__inv_2_23/Y sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__o21ai_1_299/B1 sky130_fd_sc_hd__xor2_1_120/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_709 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_604 sky130_fd_sc_hd__nand2_1_604/Y sky130_fd_sc_hd__nor2_1_197/Y
+ sky130_fd_sc_hd__nor2_1_201/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_615 sky130_fd_sc_hd__xnor2_1_172/A sky130_fd_sc_hd__nand2_1_616/Y
+ sky130_fd_sc_hd__nand2_1_615/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_626 sky130_fd_sc_hd__o21ai_2_17/A1 sky130_fd_sc_hd__nor2_1_208/Y
+ sky130_fd_sc_hd__nor2_1_213/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_637 sky130_fd_sc_hd__nand2_1_637/Y sky130_fd_sc_hd__or2_0_62/A
+ sky130_fd_sc_hd__or2_0_62/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_648 sky130_fd_sc_hd__xnor2_1_183/A sky130_fd_sc_hd__nand2_1_649/Y
+ sky130_fd_sc_hd__nand2_1_648/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_659 sky130_fd_sc_hd__o21a_1_5/B1 sky130_fd_sc_hd__nor2_1_220/A
+ sky130_fd_sc_hd__xor2_1_635/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_400 sky130_fd_sc_hd__dfxtp_1_400/Q sky130_fd_sc_hd__clkinv_4_8/Y
+ sky130_fd_sc_hd__nor2b_1_115/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1708 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_411 sky130_fd_sc_hd__dfxtp_1_411/Q sky130_fd_sc_hd__dfxtp_1_423/CLK
+ sky130_fd_sc_hd__nor2b_1_104/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1719 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_2_18 sky130_fd_sc_hd__inv_2_18/A sky130_fd_sc_hd__inv_2_18/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_422 sky130_fd_sc_hd__dfxtp_1_422/Q sky130_fd_sc_hd__dfxtp_1_423/CLK
+ sky130_fd_sc_hd__nor2b_1_93/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_29 sky130_fd_sc_hd__inv_2_29/A sky130_fd_sc_hd__inv_2_29/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_433 sky130_fd_sc_hd__dfxtp_1_433/Q sky130_fd_sc_hd__dfxtp_1_439/CLK
+ sky130_fd_sc_hd__nor2b_1_114/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_444 sky130_fd_sc_hd__dfxtp_1_444/Q sky130_fd_sc_hd__dfxtp_1_446/CLK
+ sky130_fd_sc_hd__nor2b_1_103/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_455 sky130_fd_sc_hd__dfxtp_1_455/Q sky130_fd_sc_hd__clkinv_4_9/Y
+ sky130_fd_sc_hd__nor2b_1_92/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_466 sky130_fd_sc_hd__ha_2_47/A sky130_fd_sc_hd__dfxtp_1_515/CLK
+ sky130_fd_sc_hd__and2_0_355/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_477 sky130_fd_sc_hd__dfxtp_1_477/Q sky130_fd_sc_hd__dfxtp_1_480/CLK
+ sky130_fd_sc_hd__and2_0_385/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_488 sky130_fd_sc_hd__ha_2_33/A sky130_fd_sc_hd__dfxtp_1_489/CLK
+ sky130_fd_sc_hd__and2_0_371/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_2_8 sky130_fd_sc_hd__buf_6_5/A sky130_fd_sc_hd__nand2_2_8/A
+ sky130_fd_sc_hd__nand2_2_8/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__dfxtp_1_499 sky130_fd_sc_hd__buf_4_37/A sky130_fd_sc_hd__edfxbp_1_0/CLK
+ sky130_fd_sc_hd__and2_0_399/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a222oi_1_102 vccd1 vssd1 sky130_fd_sc_hd__and3_4_5/X sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__buf_4_6/X sky130_fd_sc_hd__nor2_1_68/Y sky130_fd_sc_hd__buf_4_1/X
+ sky130_fd_sc_hd__o21ai_1_234/B1 sky130_fd_sc_hd__nor2b_1_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2b_1_14 sky130_fd_sc_hd__nand2b_1_14/Y sky130_fd_sc_hd__and3_4_15/C
+ sky130_fd_sc_hd__and3_4_15/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a222oi_1_113 vccd1 vssd1 sky130_fd_sc_hd__and3_4_1/X sky130_fd_sc_hd__nor2_2_10/B
+ sky130_fd_sc_hd__buf_6_4/X sky130_fd_sc_hd__nor2_2_9/Y sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__o21ai_1_249/B1 sky130_fd_sc_hd__and2b_4_3/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2b_1_25 sky130_fd_sc_hd__o22ai_1_92/A1 sky130_fd_sc_hd__or2_0_84/A
+ sky130_fd_sc_hd__buf_2_207/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a222oi_1_124 vccd1 vssd1 sky130_fd_sc_hd__and3_4_2/X sky130_fd_sc_hd__buf_6_4/X
+ sky130_fd_sc_hd__buf_6_0/X sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__o21ai_1_264/B1 sky130_fd_sc_hd__and2b_4_4/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_135 vccd1 vssd1 sky130_fd_sc_hd__and3_4_2/X sky130_fd_sc_hd__nor2_2_10/B
+ sky130_fd_sc_hd__buf_6_4/X sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__o21ai_1_277/B1 sky130_fd_sc_hd__and2b_4_4/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_146 vccd1 vssd1 sky130_fd_sc_hd__and3_4_1/X sky130_fd_sc_hd__buf_2_4/X
+ sky130_fd_sc_hd__buf_6_5/X sky130_fd_sc_hd__nor2_2_9/Y sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__o21ai_1_291/B1 sky130_fd_sc_hd__and2b_4_3/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_157 vccd1 vssd1 sky130_fd_sc_hd__and3_4_2/X sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__buf_6_1/X sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__o21ai_1_305/B1 sky130_fd_sc_hd__and2b_4_4/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_305 sky130_fd_sc_hd__fa_2_296/B sky130_fd_sc_hd__fa_2_306/B
+ sky130_fd_sc_hd__fa_2_305/A sky130_fd_sc_hd__fa_2_305/B sky130_fd_sc_hd__xor2_1_466/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_168 vccd1 vssd1 sky130_fd_sc_hd__and3_4_8/X sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__buf_6_2/X sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__and2_0_25/A
+ sky130_fd_sc_hd__o21ai_1_319/B1 sky130_fd_sc_hd__nor2b_2_2/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_316 sky130_fd_sc_hd__fa_2_300/A sky130_fd_sc_hd__fa_2_316/SUM
+ sky130_fd_sc_hd__fa_2_316/A sky130_fd_sc_hd__fa_2_316/B sky130_fd_sc_hd__fa_2_316/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_179 vccd1 vssd1 sky130_fd_sc_hd__and3_4_2/X sky130_fd_sc_hd__nor2_2_5/A
+ sky130_fd_sc_hd__nor2_2_5/B sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__nor2_2_4/B
+ sky130_fd_sc_hd__o21ai_1_336/B1 sky130_fd_sc_hd__and2b_4_4/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_327 sky130_fd_sc_hd__fa_2_319/B sky130_fd_sc_hd__fa_2_331/A
+ sky130_fd_sc_hd__fa_2_327/A sky130_fd_sc_hd__fa_2_327/B sky130_fd_sc_hd__fa_2_327/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_338 sky130_fd_sc_hd__fa_2_327/CIN sky130_fd_sc_hd__fa_2_340/A
+ sky130_fd_sc_hd__fa_2_338/A sky130_fd_sc_hd__fa_2_338/B sky130_fd_sc_hd__xor2_1_503/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_349 sky130_fd_sc_hd__fa_2_345/CIN sky130_fd_sc_hd__fa_2_355/A
+ sky130_fd_sc_hd__fa_2_349/A sky130_fd_sc_hd__fa_2_349/B sky130_fd_sc_hd__fa_2_353/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_8_10 sky130_fd_sc_hd__clkinv_8_11/A sky130_fd_sc_hd__clkinv_8_10/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_21 sky130_fd_sc_hd__clkinv_8_21/Y sky130_fd_sc_hd__clkinv_8_22/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_32 sky130_fd_sc_hd__clkinv_8_32/Y sky130_fd_sc_hd__clkinv_8_80/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_43 sky130_fd_sc_hd__clkinv_8_43/Y sky130_fd_sc_hd__clkinv_8_43/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_54 sky130_fd_sc_hd__clkinv_8_54/Y sky130_fd_sc_hd__clkinv_8_58/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_65 sky130_fd_sc_hd__clkinv_8_65/Y sky130_fd_sc_hd__clkinv_8_65/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_76 sky130_fd_sc_hd__clkinv_8_76/Y sky130_fd_sc_hd__clkinv_8_76/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_30 sky130_fd_sc_hd__buf_12_30/A sky130_fd_sc_hd__buf_12_30/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_8_87 sky130_fd_sc_hd__clkinv_8_88/A sky130_fd_sc_hd__clkinv_8_87/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_41 sky130_fd_sc_hd__buf_12_41/A sky130_fd_sc_hd__buf_12_41/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_52 sky130_fd_sc_hd__buf_12_52/A sky130_fd_sc_hd__buf_12_52/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_63 sky130_fd_sc_hd__inv_2_190/Y sky130_fd_sc_hd__buf_12_63/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_74 sky130_fd_sc_hd__buf_8_131/X sky130_fd_sc_hd__buf_12_74/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_85 sky130_fd_sc_hd__buf_8_23/X sky130_fd_sc_hd__buf_12_85/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_96 sky130_fd_sc_hd__buf_8_93/X sky130_fd_sc_hd__buf_12_96/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_2_3 vccd1 vssd1 sky130_fd_sc_hd__buf_2_3/X sky130_fd_sc_hd__buf_2_3/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__inv_2_3 sky130_fd_sc_hd__inv_2_3/A sky130_fd_sc_hd__inv_2_3/Y vccd1
+ vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__nor2_1_13 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_13/Y
+ sky130_fd_sc_hd__nor2_1_13/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_24 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_24/Y
+ sky130_fd_sc_hd__nor2_1_24/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_35 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_35/Y
+ sky130_fd_sc_hd__nor2_1_35/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_46 sky130_fd_sc_hd__nor2_1_50/A sky130_fd_sc_hd__nor2_1_46/Y
+ sky130_fd_sc_hd__nor2_1_46/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_57 sky130_fd_sc_hd__nor2_1_57/B sky130_fd_sc_hd__nor2_1_57/Y
+ sky130_fd_sc_hd__nor2_1_60/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_68 sky130_fd_sc_hd__and3_4_5/A sky130_fd_sc_hd__nor2_1_68/Y
+ sky130_fd_sc_hd__and3_4_5/C vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_79 sky130_fd_sc_hd__nor2_1_80/Y sky130_fd_sc_hd__nor2_1_79/Y
+ sky130_fd_sc_hd__nor2_1_83/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_12_506 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_517 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_401 sky130_fd_sc_hd__xnor2_1_93/A sky130_fd_sc_hd__nand2_1_402/Y
+ sky130_fd_sc_hd__or2_0_44/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_528 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_412 sky130_fd_sc_hd__nor2_1_132/A sky130_fd_sc_hd__nor2_1_133/Y
+ sky130_fd_sc_hd__nor2_1_136/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_539 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__and2_0_90 vccd1 vssd1 sky130_fd_sc_hd__and2_0_90/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__or2_0_9/B vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_423 sky130_fd_sc_hd__xnor2_1_102/A sky130_fd_sc_hd__nand2_1_424/Y
+ sky130_fd_sc_hd__nand2_1_423/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_434 sky130_fd_sc_hd__xnor2_1_105/A sky130_fd_sc_hd__nand2_1_435/Y
+ sky130_fd_sc_hd__nand2_1_434/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_445 sky130_fd_sc_hd__nand2_1_445/Y sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__buf_6_1/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_456 sky130_fd_sc_hd__xor2_1_399/A sky130_fd_sc_hd__nand2_1_457/Y
+ sky130_fd_sc_hd__nand2_1_456/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_467 sky130_fd_sc_hd__xnor2_1_65/B sky130_fd_sc_hd__nand2_1_468/Y
+ sky130_fd_sc_hd__nand2_1_467/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_478 sky130_fd_sc_hd__nand2_1_478/Y sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__buf_8_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_489 sky130_fd_sc_hd__o21a_1_3/B1 sky130_fd_sc_hd__a211o_1_1/X
+ sky130_fd_sc_hd__xor2_1_422/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_14 sky130_fd_sc_hd__and3_1_2/C sky130_fd_sc_hd__nor2b_1_14/Y
+ sky130_fd_sc_hd__and3_1_2/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_25 sky130_fd_sc_hd__or2_0_84/A sky130_fd_sc_hd__fa_2_457/A
+ sky130_fd_sc_hd__nor2b_1_25/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_36 sky130_fd_sc_hd__or2_0_73/A sky130_fd_sc_hd__fa_2_469/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1003 sky130_fd_sc_hd__clkinv_1_1003/Y sky130_fd_sc_hd__clkinv_1_1003/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_47 sky130_fd_sc_hd__mux2_2_22/X sky130_fd_sc_hd__nor2b_1_47/Y
+ sky130_fd_sc_hd__buf_2_214/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1014 sky130_fd_sc_hd__clkinv_1_1015/A sky130_fd_sc_hd__clkinv_2_0/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_58 sky130_fd_sc_hd__mux2_2_47/X sky130_fd_sc_hd__fa_2_480/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1025 sky130_fd_sc_hd__buf_12_30/A sky130_fd_sc_hd__clkinv_2_38/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_69 sky130_fd_sc_hd__or2_0_80/B sky130_fd_sc_hd__nor2b_1_69/Y
+ sky130_fd_sc_hd__mux2_4_5/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1036 sky130_fd_sc_hd__inv_4_13/A sky130_fd_sc_hd__inv_2_74/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1047 sky130_fd_sc_hd__inv_2_180/A sky130_fd_sc_hd__buf_8_27/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1505 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1058 sky130_fd_sc_hd__clkbuf_4_31/A sky130_fd_sc_hd__buf_8_58/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1516 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1069 sky130_fd_sc_hd__a31o_1_0/A3 sky130_fd_sc_hd__nand2_1_856/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1527 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_230 sky130_fd_sc_hd__xnor2_1_99/A sky130_fd_sc_hd__dfxtp_1_230/CLK
+ sky130_fd_sc_hd__and2_0_87/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1538 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_241 sky130_fd_sc_hd__fa_2_198/A sky130_fd_sc_hd__clkinv_4_4/Y
+ sky130_fd_sc_hd__and2_0_97/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1549 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_252 sky130_fd_sc_hd__xor2_1_197/A sky130_fd_sc_hd__dfxtp_1_264/CLK
+ sky130_fd_sc_hd__and2_0_26/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_263 sky130_fd_sc_hd__xor2_1_131/A sky130_fd_sc_hd__dfxtp_1_266/CLK
+ sky130_fd_sc_hd__and2_0_84/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_274 sky130_fd_sc_hd__xnor2_1_8/A sky130_fd_sc_hd__dfxtp_1_275/CLK
+ sky130_fd_sc_hd__and2_0_99/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_285 sky130_fd_sc_hd__dfxtp_1_285/Q sky130_fd_sc_hd__dfxtp_1_2/CLK
+ sky130_fd_sc_hd__and2_0_261/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_296 sky130_fd_sc_hd__dfxtp_1_296/Q sky130_fd_sc_hd__clkinv_8_6/Y
+ sky130_fd_sc_hd__and2_0_272/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o22ai_1_5 sky130_fd_sc_hd__o22ai_1_5/A2 sky130_fd_sc_hd__o22ai_1_5/B1
+ sky130_fd_sc_hd__o22ai_1_5/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__o22ai_1_9/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_102 sky130_fd_sc_hd__fa_2_94/CIN sky130_fd_sc_hd__fa_2_100/B
+ sky130_fd_sc_hd__fa_2_102/A sky130_fd_sc_hd__fa_2_102/B sky130_fd_sc_hd__xor2_1_138/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_113 sky130_fd_sc_hd__fa_2_112/CIN sky130_fd_sc_hd__fah_1_1/B
+ sky130_fd_sc_hd__fa_2_113/A sky130_fd_sc_hd__fa_2_113/B sky130_fd_sc_hd__xor2_1_158/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_124 sky130_fd_sc_hd__fa_2_123/B sky130_fd_sc_hd__fa_2_126/CIN
+ sky130_fd_sc_hd__fa_2_124/A sky130_fd_sc_hd__fa_2_124/B sky130_fd_sc_hd__xor2_1_172/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_135 sky130_fd_sc_hd__fa_2_133/B sky130_fd_sc_hd__fa_2_136/A
+ sky130_fd_sc_hd__fa_2_135/A sky130_fd_sc_hd__fa_2_135/B sky130_fd_sc_hd__fa_2_135/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_146 sky130_fd_sc_hd__xor3_1_11/A sky130_fd_sc_hd__fa_2_147/B
+ sky130_fd_sc_hd__fa_2_146/A sky130_fd_sc_hd__fa_2_146/B sky130_fd_sc_hd__fa_2_146/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_157 sky130_fd_sc_hd__fa_2_142/B sky130_fd_sc_hd__fa_2_159/CIN
+ sky130_fd_sc_hd__fa_2_157/A sky130_fd_sc_hd__fa_2_157/B sky130_fd_sc_hd__fa_2_158/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_168 sky130_fd_sc_hd__fa_2_159/A sky130_fd_sc_hd__fa_2_168/SUM
+ sky130_fd_sc_hd__fa_2_168/A sky130_fd_sc_hd__fa_2_168/B sky130_fd_sc_hd__fa_2_168/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and3_4_7 sky130_fd_sc_hd__nor2_2_7/B sky130_fd_sc_hd__and3_4_7/B
+ sky130_fd_sc_hd__nor2_2_7/A sky130_fd_sc_hd__and3_4_7/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__fa_2_179 sky130_fd_sc_hd__fa_2_172/CIN sky130_fd_sc_hd__fa_2_181/B
+ sky130_fd_sc_hd__fa_2_179/A sky130_fd_sc_hd__fa_2_179/B sky130_fd_sc_hd__xor2_1_271/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o22ai_1_12 sky130_fd_sc_hd__o22ai_1_51/B1 sky130_fd_sc_hd__o22ai_1_12/B1
+ sky130_fd_sc_hd__o22ai_1_12/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__inv_4_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_130 vccd1 vssd1 sky130_fd_sc_hd__buf_2_130/X la_data_out[93]
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_23 sky130_fd_sc_hd__o22ai_1_40/B1 sky130_fd_sc_hd__o22ai_1_23/B1
+ sky130_fd_sc_hd__o22ai_1_23/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__inv_4_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_141 vccd1 vssd1 sky130_fd_sc_hd__buf_8_76/A sky130_fd_sc_hd__buf_2_52/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_34 sky130_fd_sc_hd__nor2_1_31/A sky130_fd_sc_hd__o22ai_1_34/B1
+ sky130_fd_sc_hd__o22ai_1_34/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_152 vccd1 vssd1 sky130_fd_sc_hd__mux2_2_1/A0 sky130_fd_sc_hd__buf_2_152/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_45 sky130_fd_sc_hd__nor2_1_22/A sky130_fd_sc_hd__o22ai_1_45/B1
+ sky130_fd_sc_hd__o22ai_1_45/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_163 vccd1 vssd1 sky130_fd_sc_hd__buf_8_118/A sky130_fd_sc_hd__inv_2_81/Y
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_56 sky130_fd_sc_hd__nor2_1_11/A sky130_fd_sc_hd__o22ai_1_7/A2
+ sky130_fd_sc_hd__o22ai_1_56/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_174 vccd1 vssd1 sky130_fd_sc_hd__nor2_4_0/A la_data_out[33]
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_67 sky130_fd_sc_hd__xnor2_2_5/Y sky130_fd_sc_hd__xnor2_1_221/Y
+ sky130_fd_sc_hd__fa_2_425/B sky130_fd_sc_hd__xnor2_1_257/Y sky130_fd_sc_hd__o22ai_1_95/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_185 vccd1 vssd1 sky130_fd_sc_hd__buf_2_40/A sky130_fd_sc_hd__buf_2_39/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_78 sky130_fd_sc_hd__nor2b_1_20/A sky130_fd_sc_hd__o22ai_1_78/B1
+ sky130_fd_sc_hd__fa_2_436/B sky130_fd_sc_hd__o22ai_1_78/A1 sky130_fd_sc_hd__o22ai_1_78/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_196 vccd1 vssd1 la_data_out[76] sky130_fd_sc_hd__buf_2_211/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_89 sky130_fd_sc_hd__xnor2_2_6/Y sky130_fd_sc_hd__xnor2_1_237/Y
+ sky130_fd_sc_hd__o22ai_1_89/Y sky130_fd_sc_hd__xnor2_1_249/Y sky130_fd_sc_hd__o22ai_1_98/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_4_14 vccd1 vssd1 sky130_fd_sc_hd__buf_4_14/X sky130_fd_sc_hd__buf_4_14/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_25 vccd1 vssd1 sky130_fd_sc_hd__buf_4_25/X sky130_fd_sc_hd__buf_4_25/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_36 vccd1 vssd1 sky130_fd_sc_hd__buf_4_36/X sky130_fd_sc_hd__buf_8_61/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_12_107 sky130_fd_sc_hd__buf_8_136/X sky130_fd_sc_hd__buf_12_364/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_30 vssd1 vccd1 sky130_fd_sc_hd__and2_0_87/A sky130_fd_sc_hd__buf_6_4/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_118 sky130_fd_sc_hd__buf_12_24/X sky130_fd_sc_hd__buf_12_321/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_41 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_41/X sky130_fd_sc_hd__buf_2_186/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_129 sky130_fd_sc_hd__buf_12_37/X sky130_fd_sc_hd__buf_12_325/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_52 vssd1 vccd1 sky130_fd_sc_hd__buf_8_53/A sky130_fd_sc_hd__clkbuf_1_52/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_63 vssd1 vccd1 sky130_fd_sc_hd__buf_12_33/A sky130_fd_sc_hd__buf_8_2/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_74 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_14/A1 sky130_fd_sc_hd__clkbuf_1_74/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_85 vssd1 vccd1 sky130_fd_sc_hd__mux2_8_1/A1 sky130_fd_sc_hd__clkbuf_1_85/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_96 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_35/A1 sky130_fd_sc_hd__clkbuf_1_96/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkinv_1_307 sky130_fd_sc_hd__nor2_4_1/B sky130_fd_sc_hd__nor2b_1_1/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_318 sky130_fd_sc_hd__nand2_1_170/A sky130_fd_sc_hd__nor2_1_50/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_329 sky130_fd_sc_hd__nor2_1_53/B sky130_fd_sc_hd__nand2_1_194/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__or2_0_10 sky130_fd_sc_hd__or2_0_58/A sky130_fd_sc_hd__or2_0_10/X
+ sky130_fd_sc_hd__or2_0_9/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_21 sky130_fd_sc_hd__or2_0_21/A sky130_fd_sc_hd__or2_0_21/X
+ sky130_fd_sc_hd__or2_0_21/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_32 sky130_fd_sc_hd__or2_0_32/A sky130_fd_sc_hd__or2_0_32/X
+ sky130_fd_sc_hd__or2_0_32/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_43 sky130_fd_sc_hd__or2_0_43/A sky130_fd_sc_hd__or2_0_43/X
+ sky130_fd_sc_hd__or2_0_43/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_54 sky130_fd_sc_hd__or2_0_9/A sky130_fd_sc_hd__or2_0_54/X
+ sky130_fd_sc_hd__or2_0_4/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_65 sky130_fd_sc_hd__buf_4_5/X sky130_fd_sc_hd__or2_0_65/X
+ sky130_fd_sc_hd__buf_4_4/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_76 sky130_fd_sc_hd__or2_0_76/A sky130_fd_sc_hd__or2_0_76/X
+ sky130_fd_sc_hd__or2_0_76/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_87 sky130_fd_sc_hd__or2_0_87/A sky130_fd_sc_hd__or2_0_87/X
+ sky130_fd_sc_hd__or2_0_87/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_98 sky130_fd_sc_hd__or2_0_98/A sky130_fd_sc_hd__or2_0_98/X
+ sky130_fd_sc_hd__or2_0_98/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__buf_12_630 sky130_fd_sc_hd__buf_12_630/A sky130_fd_sc_hd__buf_12_630/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_4_101 sky130_fd_sc_hd__clkinv_8_55/A sky130_fd_sc_hd__dfxtp_1_29/CLK
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_12_641 sky130_fd_sc_hd__buf_12_641/A sky130_fd_sc_hd__buf_12_641/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_4_112 sky130_fd_sc_hd__clkinv_8_66/Y sky130_fd_sc_hd__clkinv_8_67/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_12_652 sky130_fd_sc_hd__buf_12_652/A sky130_fd_sc_hd__buf_12_652/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_4_123 sky130_fd_sc_hd__clkinv_8_83/Y sky130_fd_sc_hd__clkinv_8_87/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_12_663 sky130_fd_sc_hd__buf_12_663/A sky130_fd_sc_hd__buf_12_663/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_674 sky130_fd_sc_hd__buf_12_674/A sky130_fd_sc_hd__buf_12_678/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_303 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_314 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_325 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_336 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_220 sky130_fd_sc_hd__xnor2_1_26/A sky130_fd_sc_hd__nand2_1_221/Y
+ sky130_fd_sc_hd__or2_0_17/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_347 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_231 sky130_fd_sc_hd__nand2_1_231/Y sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__buf_4_2/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_358 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_830 sky130_fd_sc_hd__clkinv_1_830/Y sky130_fd_sc_hd__nand2_1_839/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_242 sky130_fd_sc_hd__o21ai_2_7/A1 sky130_fd_sc_hd__nand2_1_248/A
+ sky130_fd_sc_hd__nor2_1_79/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_369 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_841 sky130_fd_sc_hd__buf_8_59/A sky130_fd_sc_hd__inv_2_79/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_253 sky130_fd_sc_hd__nand2_1_253/Y sky130_fd_sc_hd__buf_6_4/X
+ sky130_fd_sc_hd__nor2_2_10/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_852 sky130_fd_sc_hd__clkbuf_1_36/A sky130_fd_sc_hd__clkinv_8_8/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_264 sky130_fd_sc_hd__nand2_1_264/Y sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__nor2_1_85/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_863 sky130_fd_sc_hd__clkinv_1_863/Y sky130_fd_sc_hd__inv_2_94/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_275 sky130_fd_sc_hd__xor2_1_176/B sky130_fd_sc_hd__nand2_1_276/Y
+ sky130_fd_sc_hd__nand2_1_275/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_874 sky130_fd_sc_hd__clkinv_1_874/Y sky130_fd_sc_hd__clkinv_4_84/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_286 sky130_fd_sc_hd__nand2_1_286/Y sky130_fd_sc_hd__nor2_1_97/A
+ sky130_fd_sc_hd__nor2_1_97/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_885 sky130_fd_sc_hd__clkinv_1_885/Y sky130_fd_sc_hd__clkinv_4_87/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_297 sky130_fd_sc_hd__nand2_1_297/Y sky130_fd_sc_hd__nor2_2_5/A
+ sky130_fd_sc_hd__buf_4_1/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_896 sky130_fd_sc_hd__clkinv_1_897/A sky130_fd_sc_hd__buf_2_46/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__conb_1_30 sky130_fd_sc_hd__conb_1_30/LO sky130_fd_sc_hd__conb_1_30/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1302 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_2_2 vccd1 vssd1 sky130_fd_sc_hd__xor2_2_2/X sky130_fd_sc_hd__xor2_2_2/B
+ sky130_fd_sc_hd__xor2_2_2/A vssd1 vccd1 sky130_fd_sc_hd__xor2_2
Xsky130_fd_sc_hd__conb_1_41 sky130_fd_sc_hd__conb_1_41/LO sky130_fd_sc_hd__conb_1_41/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1313 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_52 sky130_fd_sc_hd__conb_1_52/LO sky130_fd_sc_hd__conb_1_52/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1324 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_63 sky130_fd_sc_hd__conb_1_63/LO sky130_fd_sc_hd__conb_1_63/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1335 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_74 sky130_fd_sc_hd__conb_1_74/LO sky130_fd_sc_hd__conb_1_74/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1346 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_85 sky130_fd_sc_hd__conb_1_85/LO sky130_fd_sc_hd__conb_1_85/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1357 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_96 sky130_fd_sc_hd__conb_1_96/LO sky130_fd_sc_hd__conb_1_96/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1368 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1379 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__mux2_2_3 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_3/A1 sky130_fd_sc_hd__buf_4_24/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__or2_0_83/A vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__decap_12_870 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_881 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_892 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_604 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__fa_2_402/B
+ sky130_fd_sc_hd__xor2_1_604/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_615 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__fa_2_407/A
+ sky130_fd_sc_hd__xor2_1_615/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_626 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__or2_0_69/A
+ sky130_fd_sc_hd__xor2_1_626/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_637 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__nor2_4_15/B
+ sky130_fd_sc_hd__xor2_1_637/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_648 sky130_fd_sc_hd__xor2_1_648/B sky130_fd_sc_hd__xor2_1_648/X
+ sky130_fd_sc_hd__xor2_1_648/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_659 sky130_fd_sc_hd__xor2_1_659/B sky130_fd_sc_hd__xor2_1_659/X
+ sky130_fd_sc_hd__xor2_1_659/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a211o_1_17 vssd1 vccd1 sky130_fd_sc_hd__fa_2_244/A sky130_fd_sc_hd__dfxtp_1_80/Q
+ sky130_fd_sc_hd__nor2_1_21/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_17/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__a211o_1_28 vssd1 vccd1 sky130_fd_sc_hd__fa_2_161/A sky130_fd_sc_hd__dfxtp_1_91/Q
+ sky130_fd_sc_hd__nor2_1_32/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_28/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__clkinv_1_104 io_oeb[35] sky130_fd_sc_hd__conb_1_38/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_115 io_oeb[24] sky130_fd_sc_hd__conb_1_27/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_126 io_oeb[13] sky130_fd_sc_hd__conb_1_16/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_137 io_oeb[2] sky130_fd_sc_hd__conb_1_5/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_148 sky130_fd_sc_hd__o21ai_2_2/A1 sky130_fd_sc_hd__nor2_1_2/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_159 sky130_fd_sc_hd__o21ai_1_4/A2 sky130_fd_sc_hd__dfxtp_1_122/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_17 sky130_fd_sc_hd__inv_2_66/Y sky130_fd_sc_hd__nor2_1_237/B
+ sky130_fd_sc_hd__a22o_1_17/X sky130_fd_sc_hd__nor2_1_233/Y sky130_fd_sc_hd__a22o_1_17/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_28 sky130_fd_sc_hd__buf_2_63/A sky130_fd_sc_hd__buf_2_103/X
+ sky130_fd_sc_hd__a22o_1_28/X sky130_fd_sc_hd__a22o_1_28/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_39 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__buf_2_114/X
+ sky130_fd_sc_hd__a22o_1_39/X sky130_fd_sc_hd__a22o_1_39/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__o21ai_1_4 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_4/A2 sky130_fd_sc_hd__nor2_4_4/B
+ sky130_fd_sc_hd__o21ai_1_4/B1 sky130_fd_sc_hd__fa_2_28/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2_1_220 sky130_fd_sc_hd__xor2_1_635/X sky130_fd_sc_hd__o21a_1_5/A2
+ sky130_fd_sc_hd__nor2_1_220/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_231 sky130_fd_sc_hd__xnor2_2_4/A sky130_fd_sc_hd__nor2_1_231/Y
+ sky130_fd_sc_hd__buf_4_41/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_242 sky130_fd_sc_hd__nor2_1_243/Y sky130_fd_sc_hd__nor2_1_242/Y
+ sky130_fd_sc_hd__nor2_1_244/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_253 sky130_fd_sc_hd__nor2_1_253/B sky130_fd_sc_hd__nor2_1_253/Y
+ sky130_fd_sc_hd__nor2_1_253/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_2_7 sky130_fd_sc_hd__clkinv_2_7/Y sky130_fd_sc_hd__clkinv_2_7/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__nor2_1_264 sky130_fd_sc_hd__nor2_1_264/B sky130_fd_sc_hd__nor2_1_264/Y
+ sky130_fd_sc_hd__nor2_1_264/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_275 sky130_fd_sc_hd__o31ai_1_0/A1 sky130_fd_sc_hd__nor2_1_275/Y
+ sky130_fd_sc_hd__nor2_1_275/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_460 sky130_fd_sc_hd__buf_12_460/A sky130_fd_sc_hd__buf_12_512/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_471 sky130_fd_sc_hd__buf_12_471/A sky130_fd_sc_hd__buf_12_471/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_100 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_482 sky130_fd_sc_hd__buf_12_482/A sky130_fd_sc_hd__buf_12_620/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_111 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_493 sky130_fd_sc_hd__buf_12_493/A sky130_fd_sc_hd__buf_12_520/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_122 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_133 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_144 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_155 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_166 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_201 vssd1 vccd1 sky130_fd_sc_hd__buf_2_207/X sky130_fd_sc_hd__nor2b_1_20/A
+ la_data_out[84] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_177 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_212 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_212/B sky130_fd_sc_hd__a22o_1_7/B1
+ sky130_fd_sc_hd__xnor2_1_212/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_188 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_660 sky130_fd_sc_hd__nand2_1_725/A sky130_fd_sc_hd__nor2_1_235/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_18 sky130_fd_sc_hd__nand2_8_0/B sky130_fd_sc_hd__nand2_1_8/B
+ sky130_fd_sc_hd__or2_1_11/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_223 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_4/B sky130_fd_sc_hd__xnor2_1_223/Y
+ sky130_fd_sc_hd__mux2_4_2/X vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_199 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_671 sky130_fd_sc_hd__clkinv_1_671/Y sky130_fd_sc_hd__nand2_1_742/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_29 sky130_fd_sc_hd__nand2_2_8/B sky130_fd_sc_hd__nand2_1_8/B
+ sky130_fd_sc_hd__mux2_2_46/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_234 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_4/B sky130_fd_sc_hd__xnor2_1_234/Y
+ sky130_fd_sc_hd__or2_0_84/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_682 sky130_fd_sc_hd__xnor2_1_213/B sky130_fd_sc_hd__a21oi_1_164/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_245 vssd1 vccd1 la_data_out[77] sky130_fd_sc_hd__xnor2_1_245/Y
+ la_data_out[72] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_693 sky130_fd_sc_hd__clkinv_1_693/Y sky130_fd_sc_hd__nand2_1_771/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_256 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_4/B sky130_fd_sc_hd__xnor2_1_256/Y
+ sky130_fd_sc_hd__or2_0_80/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_267 vssd1 vccd1 la_data_out[85] sky130_fd_sc_hd__xnor2_1_267/Y
+ sky130_fd_sc_hd__buf_4_41/X vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_278 vssd1 vccd1 la_data_out[85] sky130_fd_sc_hd__xnor2_1_278/Y
+ la_data_out[72] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_289 vssd1 vccd1 la_data_out[77] sky130_fd_sc_hd__xnor2_1_289/Y
+ sky130_fd_sc_hd__or2_0_77/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_1110 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1121 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1132 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1143 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1154 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand3_1_0 sky130_fd_sc_hd__inv_2_6/A sky130_fd_sc_hd__nand3_1_3/A
+ sky130_fd_sc_hd__nand3_1_3/C sky130_fd_sc_hd__nor2_1_38/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__decap_12_1165 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1176 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_607 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_403/B sky130_fd_sc_hd__nor2_1_155/Y
+ sky130_fd_sc_hd__nand2_1_461/Y sky130_fd_sc_hd__o21ai_1_607/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1187 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_618 vssd1 vccd1 sky130_fd_sc_hd__nand2_1_469/Y sky130_fd_sc_hd__a21oi_1_102/Y
+ sky130_fd_sc_hd__a21oi_1_99/Y sky130_fd_sc_hd__xnor2_1_117/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1198 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_629 vssd1 vccd1 sky130_fd_sc_hd__inv_2_27/Y sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__nand2_1_331/Y sky130_fd_sc_hd__xor2_1_423/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fah_1_5 sky130_fd_sc_hd__fah_1_5/COUT sky130_fd_sc_hd__fah_1_5/B
+ sky130_fd_sc_hd__fah_1_5/A sky130_fd_sc_hd__fa_2_255/A sky130_fd_sc_hd__fah_1_5/CI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__fah_1
Xsky130_fd_sc_hd__sdlclkp_2_12 sky130_fd_sc_hd__conb_1_145/LO sky130_fd_sc_hd__clkinv_4_99/Y
+ sky130_fd_sc_hd__dfxtp_1_417/CLK sky130_fd_sc_hd__o21ai_1_891/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__a222oi_1_80 vccd1 vssd1 sky130_fd_sc_hd__and3_4_2/X sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__buf_4_5/X sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__a222oi_1_80/Y sky130_fd_sc_hd__and2b_4_4/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_91 vccd1 vssd1 sky130_fd_sc_hd__and3_4_1/X sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__nor2_1_73/B sky130_fd_sc_hd__nor2_2_9/Y sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__a222oi_1_91/Y sky130_fd_sc_hd__and2b_4_3/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__xnor2_1_60 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_60/B sky130_fd_sc_hd__xnor2_1_60/Y
+ sky130_fd_sc_hd__xnor2_1_60/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_401 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__xor2_1_401/X
+ sky130_fd_sc_hd__xor2_1_401/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_71 vssd1 vccd1 sky130_fd_sc_hd__fa_2_170/A sky130_fd_sc_hd__xnor2_1_71/Y
+ sky130_fd_sc_hd__xnor2_1_71/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_412 sky130_fd_sc_hd__fa_2_281/A sky130_fd_sc_hd__xor2_1_412/X
+ sky130_fd_sc_hd__xor2_1_412/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_82 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_82/B sky130_fd_sc_hd__xnor2_1_82/Y
+ sky130_fd_sc_hd__xnor2_1_82/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_423 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__xor2_1_423/X
+ sky130_fd_sc_hd__xor2_1_423/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_93 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_93/B sky130_fd_sc_hd__inv_2_39/A
+ sky130_fd_sc_hd__xnor2_1_93/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_434 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__xor3_1_29/C
+ sky130_fd_sc_hd__xor2_1_434/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_445 sky130_fd_sc_hd__fa_2_310/A sky130_fd_sc_hd__fa_2_288/B
+ sky130_fd_sc_hd__xor2_1_445/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_456 sky130_fd_sc_hd__fa_2_357/A sky130_fd_sc_hd__fa_2_295/B
+ sky130_fd_sc_hd__xor2_1_456/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_467 sky130_fd_sc_hd__fa_2_379/A sky130_fd_sc_hd__fa_2_305/B
+ sky130_fd_sc_hd__xor2_1_467/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_478 sky130_fd_sc_hd__fa_2_357/A sky130_fd_sc_hd__fa_2_313/B
+ sky130_fd_sc_hd__xor2_1_478/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_489 sky130_fd_sc_hd__xor2_1_489/B sky130_fd_sc_hd__inv_2_60/A
+ sky130_fd_sc_hd__xor2_1_489/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a222oi_1_509 vccd1 vssd1 sky130_fd_sc_hd__and3_4_21/X sky130_fd_sc_hd__buf_2_24/X
+ sky130_fd_sc_hd__buf_2_27/X sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__buf_2_15/X
+ sky130_fd_sc_hd__o21ai_1_806/B1 sky130_fd_sc_hd__and2b_4_12/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nor2b_1_109 sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nor2b_1_109/Y
+ sky130_fd_sc_hd__nor2b_1_109/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__decap_12_1 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_2_12 sky130_fd_sc_hd__clkinv_2_12/Y sky130_fd_sc_hd__clkinv_2_12/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_23 sky130_fd_sc_hd__buf_8_66/A sky130_fd_sc_hd__inv_2_126/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_34 sky130_fd_sc_hd__clkinv_2_34/Y sky130_fd_sc_hd__clkinv_4_28/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_45 sky130_fd_sc_hd__clkinv_2_45/Y sky130_fd_sc_hd__clkinv_8_68/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_56 la_data_out[90] sky130_fd_sc_hd__clkinv_4_94/Y vccd1
+ vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__or2_1_5 sky130_fd_sc_hd__or2_1_5/A sky130_fd_sc_hd__or2_1_5/X sky130_fd_sc_hd__or2_1_5/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_1
Xsky130_fd_sc_hd__sdlclkp_4_8 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_8_1/Y
+ sky130_fd_sc_hd__dfxtp_1_72/CLK sky130_fd_sc_hd__o21ai_2_0/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__buf_12_290 sky130_fd_sc_hd__buf_12_290/A sky130_fd_sc_hd__buf_12_467/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_160 sky130_fd_sc_hd__xor2_1_359/X sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xor2_1_146/X sky130_fd_sc_hd__a22oi_1_160/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_171 sky130_fd_sc_hd__nand2_1_127/A sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xor2_1_176/X sky130_fd_sc_hd__a22oi_1_171/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_182 sky130_fd_sc_hd__xnor2_1_120/Y sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xnor2_1_57/Y sky130_fd_sc_hd__a22oi_1_182/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_193 sky130_fd_sc_hd__clkbuf_1_3/X sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__nor2b_1_4/Y sky130_fd_sc_hd__nor2_1_61/Y sky130_fd_sc_hd__a22oi_1_193/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22o_4_2 sky130_fd_sc_hd__nand2_1_8/B sky130_fd_sc_hd__or2_0_74/A
+ sky130_fd_sc_hd__or2_0_60/B sky130_fd_sc_hd__or2_0_74/B sky130_fd_sc_hd__nand2_1_7/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_4
Xsky130_fd_sc_hd__clkinv_1_490 sky130_fd_sc_hd__nand2_1_450/A sky130_fd_sc_hd__nor2_1_152/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_404 vssd1 vccd1 sky130_fd_sc_hd__inv_2_28/Y sky130_fd_sc_hd__nand2b_1_11/Y
+ sky130_fd_sc_hd__o21ai_1_404/B1 sky130_fd_sc_hd__xor2_1_216/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_415 vssd1 vccd1 sky130_fd_sc_hd__inv_2_35/Y sky130_fd_sc_hd__nand2b_1_8/Y
+ sky130_fd_sc_hd__o21ai_1_415/B1 sky130_fd_sc_hd__xor2_1_224/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_426 vssd1 vccd1 sky130_fd_sc_hd__inv_2_27/Y sky130_fd_sc_hd__nand2b_1_10/Y
+ sky130_fd_sc_hd__nand2_1_322/Y sky130_fd_sc_hd__ha_2_1/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_437 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_0/Y sky130_fd_sc_hd__nand2b_1_9/Y
+ sky130_fd_sc_hd__o21ai_1_437/B1 sky130_fd_sc_hd__xor2_1_242/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_448 vssd1 vccd1 sky130_fd_sc_hd__nand2_2_12/Y sky130_fd_sc_hd__nand2b_1_11/Y
+ sky130_fd_sc_hd__a22oi_1_203/Y sky130_fd_sc_hd__xor2_1_251/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_459 vssd1 vccd1 sky130_fd_sc_hd__inv_2_27/Y sky130_fd_sc_hd__nand2b_1_11/Y
+ sky130_fd_sc_hd__nand2_1_323/Y sky130_fd_sc_hd__xor2_1_261/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2_4_13 sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__nor2_4_13/A
+ sky130_fd_sc_hd__nor2_4_13/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__nand2_1_808 sky130_fd_sc_hd__xor2_1_680/B sky130_fd_sc_hd__nand2_1_809/Y
+ sky130_fd_sc_hd__nand2_1_808/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_819 sky130_fd_sc_hd__nand2_1_819/Y sky130_fd_sc_hd__or2_0_106/A
+ sky130_fd_sc_hd__or2_0_106/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_220 sky130_fd_sc_hd__dfxtp_2_5/Q sky130_fd_sc_hd__xor3_1_17/A
+ sky130_fd_sc_hd__xor2_1_220/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_231 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__xor2_1_231/X
+ sky130_fd_sc_hd__xor2_1_231/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__o21ai_1_19 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_14/B1 sky130_fd_sc_hd__inv_2_53/A
+ sky130_fd_sc_hd__o21ai_1_19/B1 sky130_fd_sc_hd__fa_2_113/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_242 sky130_fd_sc_hd__xor2_1_383/B sky130_fd_sc_hd__xor2_1_242/X
+ sky130_fd_sc_hd__xor2_1_242/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_253 sky130_fd_sc_hd__xor2_1_362/B sky130_fd_sc_hd__xor2_1_253/X
+ sky130_fd_sc_hd__xor2_1_253/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_264 sky130_fd_sc_hd__xor2_1_383/B sky130_fd_sc_hd__xor2_1_264/X
+ sky130_fd_sc_hd__xor2_1_264/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_275 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__fa_2_178/B
+ sky130_fd_sc_hd__xor2_1_275/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_286 sky130_fd_sc_hd__dfxtp_2_5/Q sky130_fd_sc_hd__fa_2_196/B
+ sky130_fd_sc_hd__xor2_1_286/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_297 sky130_fd_sc_hd__dfxtp_2_5/Q sky130_fd_sc_hd__xor2_1_297/X
+ sky130_fd_sc_hd__xor2_1_297/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_202 vssd1 vccd1 sky130_fd_sc_hd__buf_12_56/A sky130_fd_sc_hd__ha_2_36/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_213 vssd1 vccd1 sky130_fd_sc_hd__buf_8_57/A sky130_fd_sc_hd__inv_12_0/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_224 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_225/A sky130_fd_sc_hd__nand2b_1_31/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_235 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_235/X sky130_fd_sc_hd__clkbuf_1_290/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_306 vccd1 vssd1 sky130_fd_sc_hd__and3_4_16/X sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__buf_4_7/X sky130_fd_sc_hd__nor2_2_19/Y sky130_fd_sc_hd__buf_4_0/X
+ sky130_fd_sc_hd__o21ai_1_521/B1 sky130_fd_sc_hd__nor2b_2_3/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_246 vssd1 vccd1 sky130_fd_sc_hd__buf_8_128/A sky130_fd_sc_hd__clkbuf_1_306/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_317 vccd1 vssd1 sky130_fd_sc_hd__and3_4_11/X sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__and2_0_38/A sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__and2_0_49/A
+ sky130_fd_sc_hd__o21ai_1_533/B1 sky130_fd_sc_hd__and2b_4_8/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_257 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_258/A sky130_fd_sc_hd__buf_8_73/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_2_4 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__dfxtp_2_4/CLK
+ sky130_fd_sc_hd__dfxtp_2_4/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_2
Xsky130_fd_sc_hd__a222oi_1_328 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__and2_0_87/A
+ sky130_fd_sc_hd__buf_6_0/X sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__o21ai_1_548/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_268 vssd1 vccd1 sky130_fd_sc_hd__buf_8_109/A sky130_fd_sc_hd__clkbuf_1_273/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_339 vccd1 vssd1 sky130_fd_sc_hd__and3_4_17/X sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__inv_6_0/Y sky130_fd_sc_hd__nor2_2_20/Y sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__o21ai_1_563/B1 sky130_fd_sc_hd__nor2b_2_4/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_279 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_280/A sky130_fd_sc_hd__buf_6_24/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_2_80 vccd1 vssd1 sky130_fd_sc_hd__buf_2_80/X sky130_fd_sc_hd__buf_2_80/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_91 vccd1 vssd1 sky130_fd_sc_hd__buf_2_91/X sky130_fd_sc_hd__buf_2_91/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_4_7 vccd1 vssd1 sky130_fd_sc_hd__buf_4_7/X sky130_fd_sc_hd__buf_4_7/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__and2_0_200 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_82/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_82/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_211 vccd1 vssd1 sky130_fd_sc_hd__and2_0_211/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_211/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_222 vccd1 vssd1 sky130_fd_sc_hd__and2_0_222/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__o21ai_1_65/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_233 vccd1 vssd1 sky130_fd_sc_hd__and2_0_233/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__o21ai_1_56/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_244 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_91/D sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__o21ai_1_47/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_255 vccd1 vssd1 sky130_fd_sc_hd__and2_0_255/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__and2_0_255/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_266 vccd1 vssd1 sky130_fd_sc_hd__and2_0_266/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__xor2_1_645/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_277 vccd1 vssd1 sky130_fd_sc_hd__and2_0_277/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__and2_0_277/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_288 vccd1 vssd1 sky130_fd_sc_hd__and2_0_288/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_9/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__a21oi_2_18 sky130_fd_sc_hd__a21oi_2_18/B1 sky130_fd_sc_hd__or2_1_2/X
+ sky130_fd_sc_hd__o21ai_2_15/Y sky130_fd_sc_hd__xor2_1_543/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_2
Xsky130_fd_sc_hd__and2_0_299 vccd1 vssd1 sky130_fd_sc_hd__and2_0_299/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_20/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__xor3_1_20 sky130_fd_sc_hd__xor3_1_20/X sky130_fd_sc_hd__xor3_1_21/X
+ sky130_fd_sc_hd__xor3_1_20/B sky130_fd_sc_hd__xor3_1_26/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__sdlclkp_2_5 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_4_0/Y
+ sky130_fd_sc_hd__dfxtp_1_158/CLK sky130_fd_sc_hd__o21ai_1_1/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__inv_4_7 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__inv_4_7/A vccd1
+ vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__o21ai_1_201 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_209/A2 sky130_fd_sc_hd__nor2_1_50/A
+ sky130_fd_sc_hd__nor2_1_49/Y sky130_fd_sc_hd__o21ai_1_201/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_212 vssd1 vccd1 sky130_fd_sc_hd__inv_2_15/Y sky130_fd_sc_hd__nand2b_1_4/Y
+ sky130_fd_sc_hd__a222oi_1_84/Y sky130_fd_sc_hd__xor2_1_37/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_30 sky130_fd_sc_hd__clkbuf_4_30/X sky130_fd_sc_hd__buf_12_74/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_223 vssd1 vccd1 sky130_fd_sc_hd__buf_2_3/X sky130_fd_sc_hd__nand2b_1_4/Y
+ sky130_fd_sc_hd__a222oi_1_92/Y sky130_fd_sc_hd__xor2_1_47/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_41 la_data_out[58] sky130_fd_sc_hd__dfxtp_1_473/Q vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_234 vssd1 vccd1 sky130_fd_sc_hd__inv_2_16/Y sky130_fd_sc_hd__nand2b_1_5/Y
+ sky130_fd_sc_hd__o21ai_1_234/B1 sky130_fd_sc_hd__xor2_1_59/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_52 la_data_out[79] sky130_fd_sc_hd__xnor2_2_4/B vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_245 vssd1 vccd1 sky130_fd_sc_hd__inv_2_15/Y sky130_fd_sc_hd__nand2b_1_5/Y
+ sky130_fd_sc_hd__o21ai_1_245/B1 sky130_fd_sc_hd__xor2_1_68/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_256 vssd1 vccd1 sky130_fd_sc_hd__inv_2_20/Y sky130_fd_sc_hd__nand2b_1_1/Y
+ sky130_fd_sc_hd__o21ai_1_256/B1 sky130_fd_sc_hd__xor2_1_79/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_267 vssd1 vccd1 sky130_fd_sc_hd__inv_2_9/Y sky130_fd_sc_hd__nand2b_1_1/Y
+ sky130_fd_sc_hd__o21ai_1_267/B1 sky130_fd_sc_hd__xor2_1_89/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_278 vssd1 vccd1 sky130_fd_sc_hd__inv_2_23/Y sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__o21ai_1_278/B1 sky130_fd_sc_hd__xor2_1_99/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_289 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_0/Y sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__o21ai_1_289/B1 sky130_fd_sc_hd__xor2_1_110/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nand2_1_605 sky130_fd_sc_hd__xnor2_1_167/A sky130_fd_sc_hd__nand2_1_606/Y
+ sky130_fd_sc_hd__nand2_1_605/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_616 sky130_fd_sc_hd__nand2_1_616/Y sky130_fd_sc_hd__buf_2_20/X
+ sky130_fd_sc_hd__buf_2_21/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_627 sky130_fd_sc_hd__xor2_1_612/A sky130_fd_sc_hd__nand2_1_628/Y
+ sky130_fd_sc_hd__nand2_1_627/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_638 sky130_fd_sc_hd__xnor2_1_128/B sky130_fd_sc_hd__nand2_1_639/Y
+ sky130_fd_sc_hd__nand2_1_638/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_649 sky130_fd_sc_hd__nand2_1_649/Y sky130_fd_sc_hd__buf_2_30/X
+ sky130_fd_sc_hd__buf_2_29/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_401 sky130_fd_sc_hd__dfxtp_1_401/Q sky130_fd_sc_hd__clkinv_4_8/Y
+ sky130_fd_sc_hd__nor2b_1_114/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1709 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_412 sky130_fd_sc_hd__dfxtp_1_412/Q sky130_fd_sc_hd__dfxtp_1_423/CLK
+ sky130_fd_sc_hd__nor2b_1_103/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_19 sky130_fd_sc_hd__inv_2_19/A sky130_fd_sc_hd__inv_2_19/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_423 sky130_fd_sc_hd__dfxtp_1_423/Q sky130_fd_sc_hd__dfxtp_1_423/CLK
+ sky130_fd_sc_hd__nor2b_1_92/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_434 sky130_fd_sc_hd__dfxtp_1_434/Q sky130_fd_sc_hd__dfxtp_1_439/CLK
+ sky130_fd_sc_hd__nor2b_1_113/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_445 sky130_fd_sc_hd__dfxtp_1_445/Q sky130_fd_sc_hd__dfxtp_1_446/CLK
+ sky130_fd_sc_hd__nor2b_1_102/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_456 sky130_fd_sc_hd__dfxtp_1_456/Q sky130_fd_sc_hd__clkinv_4_9/Y
+ sky130_fd_sc_hd__nor2b_1_91/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_467 sky130_fd_sc_hd__ha_2_50/A sky130_fd_sc_hd__dfxtp_1_515/CLK
+ sky130_fd_sc_hd__and2_0_356/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_478 sky130_fd_sc_hd__dfxtp_1_478/Q sky130_fd_sc_hd__dfxtp_1_480/CLK
+ sky130_fd_sc_hd__and2_0_387/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_489 sky130_fd_sc_hd__dfxtp_1_489/Q sky130_fd_sc_hd__dfxtp_1_489/CLK
+ sky130_fd_sc_hd__and2_0_370/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_2_9 sky130_fd_sc_hd__nand2_2_9/Y sky130_fd_sc_hd__inv_2_6/A
+ sky130_fd_sc_hd__inv_2_7/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__a222oi_1_103 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__or2_0_66/A sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__or2_0_60/B
+ sky130_fd_sc_hd__o21ai_1_235/B1 sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2b_1_15 sky130_fd_sc_hd__nand2b_1_15/Y sky130_fd_sc_hd__nor2_2_31/A
+ sky130_fd_sc_hd__nor2_2_31/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a222oi_1_114 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__buf_4_4/X sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__o21ai_1_250/B1 sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2b_1_26 sky130_fd_sc_hd__nand2b_1_26/Y sky130_fd_sc_hd__or2_0_84/A
+ la_data_out[81] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a222oi_1_125 vccd1 vssd1 sky130_fd_sc_hd__and3_4_7/X sky130_fd_sc_hd__nor2_2_5/A
+ sky130_fd_sc_hd__nor2_2_5/B sky130_fd_sc_hd__nor2_2_7/Y sky130_fd_sc_hd__nor2_2_4/B
+ sky130_fd_sc_hd__o21ai_1_265/B1 sky130_fd_sc_hd__nor2b_2_1/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_136 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__buf_4_3/X sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__o21ai_1_278/B1 sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_147 vccd1 vssd1 sky130_fd_sc_hd__and3_4_2/X sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__nor2_1_85/B sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__nor2_2_10/B
+ sky130_fd_sc_hd__o21ai_1_292/B1 sky130_fd_sc_hd__and2b_4_4/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_158 vccd1 vssd1 sky130_fd_sc_hd__and3_4_8/X sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__and2_0_25/A sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__nor2_2_5/A
+ sky130_fd_sc_hd__o21ai_1_306/B1 sky130_fd_sc_hd__nor2b_2_2/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_306 sky130_fd_sc_hd__fa_2_297/A sky130_fd_sc_hd__fa_2_307/B
+ sky130_fd_sc_hd__fa_2_306/A sky130_fd_sc_hd__fa_2_306/B sky130_fd_sc_hd__fa_2_306/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o21ai_1_790 vssd1 vccd1 sky130_fd_sc_hd__buf_2_13/X sky130_fd_sc_hd__nand2b_1_15/Y
+ sky130_fd_sc_hd__o21ai_1_790/B1 sky130_fd_sc_hd__xor2_1_564/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_169 vccd1 vssd1 sky130_fd_sc_hd__and3_4_1/X sky130_fd_sc_hd__and2_0_25/A
+ sky130_fd_sc_hd__nor2_2_5/A sky130_fd_sc_hd__nor2_2_9/Y sky130_fd_sc_hd__nor2_2_5/B
+ sky130_fd_sc_hd__o21ai_1_320/B1 sky130_fd_sc_hd__and2b_4_3/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_317 sky130_fd_sc_hd__or2_1_8/A sky130_fd_sc_hd__nor2_2_21/B
+ sky130_fd_sc_hd__fa_2_317/A sky130_fd_sc_hd__fa_2_317/B sky130_fd_sc_hd__fa_2_317/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_328 sky130_fd_sc_hd__fa_2_323/A sky130_fd_sc_hd__fa_2_329/B
+ sky130_fd_sc_hd__fa_2_328/A sky130_fd_sc_hd__fa_2_328/B sky130_fd_sc_hd__fa_2_328/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_339 sky130_fd_sc_hd__fa_2_326/B sky130_fd_sc_hd__fa_2_339/SUM
+ sky130_fd_sc_hd__fa_2_339/A sky130_fd_sc_hd__fa_2_339/B sky130_fd_sc_hd__xor2_1_501/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_8_11 sky130_fd_sc_hd__clkinv_8_12/A sky130_fd_sc_hd__clkinv_8_11/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_22 sky130_fd_sc_hd__clkinv_8_22/Y sky130_fd_sc_hd__clkinv_8_22/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_33 sky130_fd_sc_hd__clkinv_8_34/A sky130_fd_sc_hd__clkinv_8_33/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_44 sky130_fd_sc_hd__inv_2_105/A wbs_dat_i[4] vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_55 sky130_fd_sc_hd__dfxtp_2_7/CLK sky130_fd_sc_hd__clkinv_8_55/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_66 sky130_fd_sc_hd__clkinv_8_66/Y sky130_fd_sc_hd__clkinv_8_66/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_20 sky130_fd_sc_hd__inv_2_145/Y sky130_fd_sc_hd__buf_12_20/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_8_77 sky130_fd_sc_hd__clkinv_8_78/A sky130_fd_sc_hd__clkinv_8_77/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_31 sky130_fd_sc_hd__buf_12_31/A sky130_fd_sc_hd__buf_12_31/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_8_88 sky130_fd_sc_hd__clkinv_8_89/A sky130_fd_sc_hd__clkinv_8_88/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_42 sky130_fd_sc_hd__buf_12_42/A sky130_fd_sc_hd__buf_12_42/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_53 sky130_fd_sc_hd__buf_12_53/A sky130_fd_sc_hd__buf_12_53/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_64 sky130_fd_sc_hd__buf_12_64/A sky130_fd_sc_hd__buf_12_64/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_75 sky130_fd_sc_hd__buf_8_74/X sky130_fd_sc_hd__buf_12_75/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_86 sky130_fd_sc_hd__buf_8_70/X sky130_fd_sc_hd__buf_12_86/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_97 sky130_fd_sc_hd__buf_8_22/X sky130_fd_sc_hd__buf_12_97/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_2_4 vccd1 vssd1 sky130_fd_sc_hd__buf_2_4/X sky130_fd_sc_hd__buf_2_4/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__inv_2_4 sky130_fd_sc_hd__inv_2_4/A sky130_fd_sc_hd__inv_2_4/Y vccd1
+ vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__nor2_1_14 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_14/Y
+ sky130_fd_sc_hd__nor2_1_14/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_25 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_25/Y
+ sky130_fd_sc_hd__nor2_1_25/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_36 sky130_fd_sc_hd__nor2_4_7/B sky130_fd_sc_hd__nor2_1_36/Y
+ sky130_fd_sc_hd__nor2_1_36/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_47 sky130_fd_sc_hd__nor2_1_51/B sky130_fd_sc_hd__nor2_1_47/Y
+ sky130_fd_sc_hd__nor2_1_47/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_58 sky130_fd_sc_hd__nor2_1_58/B sky130_fd_sc_hd__nor2_1_58/Y
+ sky130_fd_sc_hd__nor2_1_58/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_69 sky130_fd_sc_hd__nor2_1_69/B sky130_fd_sc_hd__nor2_1_69/Y
+ sky130_fd_sc_hd__nor2_1_69/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_12_507 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_518 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_402 sky130_fd_sc_hd__nand2_1_402/Y sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__buf_4_2/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_529 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__and2_0_80 vccd1 vssd1 sky130_fd_sc_hd__and2_0_80/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__buf_4_5/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_413 sky130_fd_sc_hd__o21ai_2_10/A1 sky130_fd_sc_hd__or2_1_0/X
+ sky130_fd_sc_hd__nor2_1_138/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_91 vccd1 vssd1 sky130_fd_sc_hd__and2_0_91/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__or2_0_9/B vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_424 sky130_fd_sc_hd__nand2_1_424/Y sky130_fd_sc_hd__buf_6_4/X
+ sky130_fd_sc_hd__nor2_2_10/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_435 sky130_fd_sc_hd__nand2_1_435/Y sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__nor2_1_85/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_446 sky130_fd_sc_hd__xor2_1_389/B sky130_fd_sc_hd__nand2_1_447/Y
+ sky130_fd_sc_hd__nand2_1_446/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_457 sky130_fd_sc_hd__nand2_1_457/Y sky130_fd_sc_hd__nor2_1_154/A
+ sky130_fd_sc_hd__nor2_1_154/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_468 sky130_fd_sc_hd__nand2_1_468/Y sky130_fd_sc_hd__buf_4_0/X
+ sky130_fd_sc_hd__buf_4_7/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_479 sky130_fd_sc_hd__xnor2_1_123/B sky130_fd_sc_hd__nand2_1_480/Y
+ sky130_fd_sc_hd__or2_0_48/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_15 sky130_fd_sc_hd__and3_4_23/C sky130_fd_sc_hd__nor2b_1_15/Y
+ sky130_fd_sc_hd__and3_4_23/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_26 sky130_fd_sc_hd__fa_2_415/B sky130_fd_sc_hd__fa_2_461/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_37 sky130_fd_sc_hd__or2_0_73/B sky130_fd_sc_hd__nor2b_1_37/Y
+ sky130_fd_sc_hd__buf_2_214/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1004 sky130_fd_sc_hd__clkinv_1_1005/A sky130_fd_sc_hd__clkinv_2_2/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_48 sky130_fd_sc_hd__or2_0_76/A sky130_fd_sc_hd__fa_2_475/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1015 sky130_fd_sc_hd__clkinv_1_1015/Y sky130_fd_sc_hd__clkinv_1_1015/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_59 sky130_fd_sc_hd__mux2_2_27/X sky130_fd_sc_hd__nor2b_1_59/Y
+ sky130_fd_sc_hd__buf_2_214/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1026 sky130_fd_sc_hd__buf_12_6/A sky130_fd_sc_hd__clkinv_2_39/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1037 sky130_fd_sc_hd__clkinv_1_1038/A sky130_fd_sc_hd__inv_8_0/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1048 sky130_fd_sc_hd__inv_2_181/A sky130_fd_sc_hd__clkbuf_4_20/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_90 sky130_fd_sc_hd__buf_8_90/A sky130_fd_sc_hd__buf_8_90/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__decap_12_1506 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1059 sky130_fd_sc_hd__inv_16_2/A sky130_fd_sc_hd__buf_8_142/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1517 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_220 sky130_fd_sc_hd__xnor2_1_124/A sky130_fd_sc_hd__dfxtp_2_5/CLK
+ sky130_fd_sc_hd__and2_0_29/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1528 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_231 sky130_fd_sc_hd__xor2_1_362/A sky130_fd_sc_hd__dfxtp_1_234/CLK
+ sky130_fd_sc_hd__and2_0_81/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1539 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_242 sky130_fd_sc_hd__xnor2_1_77/B sky130_fd_sc_hd__clkinv_4_4/Y
+ sky130_fd_sc_hd__and2_0_96/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_253 sky130_fd_sc_hd__xnor2_1_51/A sky130_fd_sc_hd__clkinv_4_6/Y
+ sky130_fd_sc_hd__and2_0_56/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_264 sky130_fd_sc_hd__fa_2_97/A sky130_fd_sc_hd__dfxtp_1_264/CLK
+ sky130_fd_sc_hd__and2_0_83/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_275 sky130_fd_sc_hd__xnor2_1_5/A sky130_fd_sc_hd__dfxtp_1_275/CLK
+ sky130_fd_sc_hd__and2_0_57/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_286 sky130_fd_sc_hd__dfxtp_1_286/Q sky130_fd_sc_hd__clkinv_8_6/Y
+ sky130_fd_sc_hd__and2_0_262/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_297 sky130_fd_sc_hd__dfxtp_1_297/Q sky130_fd_sc_hd__clkinv_8_6/Y
+ sky130_fd_sc_hd__and2_0_273/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o22ai_1_6 sky130_fd_sc_hd__o22ai_1_6/A2 sky130_fd_sc_hd__o22ai_1_6/B1
+ sky130_fd_sc_hd__o22ai_1_6/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__o22ai_1_9/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_103 sky130_fd_sc_hd__or2_0_8/A sky130_fd_sc_hd__nor2_2_3/B
+ sky130_fd_sc_hd__fa_2_103/A sky130_fd_sc_hd__fa_2_103/B sky130_fd_sc_hd__fa_2_103/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_114 sky130_fd_sc_hd__fah_1_0/B sky130_fd_sc_hd__fa_2_115/CIN
+ sky130_fd_sc_hd__fa_2_114/A sky130_fd_sc_hd__fa_2_114/B sky130_fd_sc_hd__fa_2_114/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_125 sky130_fd_sc_hd__fa_2_120/CIN sky130_fd_sc_hd__fa_2_124/B
+ sky130_fd_sc_hd__fa_2_125/A sky130_fd_sc_hd__fa_2_125/B sky130_fd_sc_hd__xor2_1_173/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_136 sky130_fd_sc_hd__nor2_1_97/A sky130_fd_sc_hd__nor2_1_98/B
+ sky130_fd_sc_hd__fa_2_136/A sky130_fd_sc_hd__fa_2_136/B sky130_fd_sc_hd__xor2_1_192/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_147 sky130_fd_sc_hd__xor3_1_10/B sky130_fd_sc_hd__fa_2_147/SUM
+ sky130_fd_sc_hd__fa_2_147/A sky130_fd_sc_hd__fa_2_147/B sky130_fd_sc_hd__fa_2_147/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_158 sky130_fd_sc_hd__fa_2_142/A sky130_fd_sc_hd__fa_2_158/SUM
+ sky130_fd_sc_hd__fa_2_158/A sky130_fd_sc_hd__fa_2_158/B sky130_fd_sc_hd__fa_2_158/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_169 sky130_fd_sc_hd__fa_2_168/CIN sky130_fd_sc_hd__fa_2_176/B
+ sky130_fd_sc_hd__fa_2_169/A sky130_fd_sc_hd__fa_2_169/B sky130_fd_sc_hd__xor2_1_256/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and3_4_8 sky130_fd_sc_hd__nor2_2_8/B sky130_fd_sc_hd__and3_4_8/B
+ sky130_fd_sc_hd__nor2_2_8/A sky130_fd_sc_hd__and3_4_8/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__buf_2_120 vccd1 vssd1 sky130_fd_sc_hd__buf_2_120/X sky130_fd_sc_hd__buf_2_120/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_13 sky130_fd_sc_hd__o22ai_1_50/B1 sky130_fd_sc_hd__o22ai_1_13/B1
+ sky130_fd_sc_hd__o22ai_1_13/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__inv_4_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_131 vccd1 vssd1 sky130_fd_sc_hd__buf_2_131/X sky130_fd_sc_hd__buf_2_131/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_24 sky130_fd_sc_hd__o22ai_1_38/B1 sky130_fd_sc_hd__o21ai_1_8/A2
+ sky130_fd_sc_hd__o22ai_1_24/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__inv_4_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_142 vccd1 vssd1 sky130_fd_sc_hd__buf_2_142/X sky130_fd_sc_hd__buf_2_142/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_35 sky130_fd_sc_hd__nor2_1_34/A sky130_fd_sc_hd__o22ai_1_35/B1
+ sky130_fd_sc_hd__o22ai_1_35/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_153 vccd1 vssd1 sky130_fd_sc_hd__buf_2_153/X sky130_fd_sc_hd__buf_2_153/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_46 sky130_fd_sc_hd__nor2_1_21/A sky130_fd_sc_hd__o22ai_1_46/B1
+ sky130_fd_sc_hd__o22ai_1_46/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_164 vccd1 vssd1 sky130_fd_sc_hd__buf_8_108/A sky130_fd_sc_hd__inv_4_13/Y
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_57 sky130_fd_sc_hd__nor2_1_10/A sky130_fd_sc_hd__o22ai_1_6/A2
+ sky130_fd_sc_hd__o22ai_1_57/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_175 vccd1 vssd1 la_data_out[65] sky130_fd_sc_hd__buf_2_175/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_68 sky130_fd_sc_hd__xnor2_2_4/Y sky130_fd_sc_hd__xnor2_1_220/Y
+ sky130_fd_sc_hd__fa_2_425/A sky130_fd_sc_hd__xnor2_1_254/Y sky130_fd_sc_hd__o22ai_1_96/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_186 vccd1 vssd1 sky130_fd_sc_hd__buf_2_41/A sky130_fd_sc_hd__buf_2_186/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_79 sky130_fd_sc_hd__xnor2_2_5/Y sky130_fd_sc_hd__xnor2_1_232/Y
+ sky130_fd_sc_hd__fa_2_436/A sky130_fd_sc_hd__xnor2_1_229/Y sky130_fd_sc_hd__o22ai_1_95/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_197 vccd1 vssd1 la_data_out[75] sky130_fd_sc_hd__or2_0_80/B
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_4_15 vccd1 vssd1 sky130_fd_sc_hd__buf_4_15/X sky130_fd_sc_hd__buf_4_15/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_26 vccd1 vssd1 sky130_fd_sc_hd__buf_8_73/A sky130_fd_sc_hd__buf_4_26/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_37 vccd1 vssd1 la_data_out[36] sky130_fd_sc_hd__buf_4_37/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__clkbuf_1_20 vssd1 vccd1 sky130_fd_sc_hd__inv_2_53/A sky130_fd_sc_hd__nor2_4_4/B
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_108 sky130_fd_sc_hd__buf_8_62/X sky130_fd_sc_hd__buf_12_449/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_31 vssd1 vccd1 sky130_fd_sc_hd__a22o_1_9/B2 sky130_fd_sc_hd__nor2_1_233/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_119 sky130_fd_sc_hd__buf_8_44/X sky130_fd_sc_hd__buf_12_119/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_42 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_42/X wbs_dat_i[10]
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_53 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_53/X sky130_fd_sc_hd__conb_1_147/HI
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_64 vssd1 vccd1 sky130_fd_sc_hd__buf_8_49/A sky130_fd_sc_hd__buf_8_34/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_75 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_17/A1 sky130_fd_sc_hd__clkbuf_1_75/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_86 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_33/A1 sky130_fd_sc_hd__clkbuf_1_86/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_97 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_4/A1 sky130_fd_sc_hd__clkbuf_1_97/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkinv_1_308 sky130_fd_sc_hd__nand2_1_291/A sky130_fd_sc_hd__nor2_2_5/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_319 sky130_fd_sc_hd__nand2_1_173/A sky130_fd_sc_hd__nor2_2_2/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__or2_0_11 sky130_fd_sc_hd__or2_0_11/A sky130_fd_sc_hd__or2_0_11/X
+ sky130_fd_sc_hd__or2_0_11/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_22 sky130_fd_sc_hd__or2_0_22/A sky130_fd_sc_hd__or2_0_22/X
+ sky130_fd_sc_hd__or2_0_22/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_33 sky130_fd_sc_hd__or2_0_33/A sky130_fd_sc_hd__or2_0_33/X
+ sky130_fd_sc_hd__or2_0_33/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_44 sky130_fd_sc_hd__buf_4_3/X sky130_fd_sc_hd__or2_0_44/X
+ sky130_fd_sc_hd__buf_4_2/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_55 sky130_fd_sc_hd__or2_0_55/A sky130_fd_sc_hd__or2_0_55/X
+ sky130_fd_sc_hd__or2_0_55/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_66 sky130_fd_sc_hd__or2_0_66/A sky130_fd_sc_hd__or2_0_66/X
+ sky130_fd_sc_hd__buf_4_5/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_77 sky130_fd_sc_hd__or2_0_77/A sky130_fd_sc_hd__or2_0_77/X
+ sky130_fd_sc_hd__or2_0_77/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_88 sky130_fd_sc_hd__or2_0_88/A sky130_fd_sc_hd__or2_0_88/X
+ sky130_fd_sc_hd__or2_0_88/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_99 sky130_fd_sc_hd__or2_0_99/A sky130_fd_sc_hd__or2_0_99/X
+ sky130_fd_sc_hd__or2_0_99/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__buf_12_620 sky130_fd_sc_hd__buf_12_620/A sky130_fd_sc_hd__buf_12_620/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_631 sky130_fd_sc_hd__buf_12_631/A sky130_fd_sc_hd__buf_12_631/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_4_102 sky130_fd_sc_hd__clkinv_8_7/A sky130_fd_sc_hd__clkinv_2_11/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_12_642 sky130_fd_sc_hd__buf_12_642/A sky130_fd_sc_hd__buf_12_642/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_4_113 sky130_fd_sc_hd__clkinv_8_68/A sky130_fd_sc_hd__edfxbp_1_0/CLK
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_12_653 sky130_fd_sc_hd__buf_12_653/A sky130_fd_sc_hd__buf_12_653/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_4_124 sky130_fd_sc_hd__clkinv_4_97/Y sky130_fd_sc_hd__clkinv_8_90/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_12_664 sky130_fd_sc_hd__buf_12_664/A sky130_fd_sc_hd__buf_12_664/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_675 sky130_fd_sc_hd__buf_12_675/A sky130_fd_sc_hd__buf_12_675/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_304 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_315 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_326 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_210 sky130_fd_sc_hd__xnor2_1_22/A sky130_fd_sc_hd__nand2_1_211/Y
+ sky130_fd_sc_hd__or2_0_13/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_337 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_221 sky130_fd_sc_hd__nand2_1_221/Y sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__buf_4_4/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_348 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_820 sky130_fd_sc_hd__clkinv_1_820/Y sky130_fd_sc_hd__nand2_1_819/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_232 sky130_fd_sc_hd__xnor2_1_32/A sky130_fd_sc_hd__nand2_1_233/Y
+ sky130_fd_sc_hd__or2_0_8/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_359 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_831 sky130_fd_sc_hd__clkinv_1_831/Y sky130_fd_sc_hd__nand2_1_843/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_243 sky130_fd_sc_hd__xnor2_1_35/A sky130_fd_sc_hd__nand2_1_244/Y
+ sky130_fd_sc_hd__or2_0_11/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_842 sky130_fd_sc_hd__inv_2_83/A la_data_out[44] vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_254 sky130_fd_sc_hd__xor2_1_154/B sky130_fd_sc_hd__nand2_1_255/Y
+ sky130_fd_sc_hd__nand2_1_254/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_853 sky130_fd_sc_hd__clkinv_1_853/Y sky130_fd_sc_hd__clkinv_8_9/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_265 sky130_fd_sc_hd__xnor2_1_44/A sky130_fd_sc_hd__nand2_1_266/Y
+ sky130_fd_sc_hd__nand2_1_265/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_864 sky130_fd_sc_hd__clkinv_1_864/Y sky130_fd_sc_hd__inv_2_94/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_276 sky130_fd_sc_hd__nand2_1_276/Y sky130_fd_sc_hd__nor2_1_91/A
+ sky130_fd_sc_hd__nor2_1_91/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_875 sky130_fd_sc_hd__clkinv_1_875/Y sky130_fd_sc_hd__clkinv_4_85/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_287 sky130_fd_sc_hd__xnor2_1_52/A sky130_fd_sc_hd__nand2_1_288/Y
+ sky130_fd_sc_hd__nand2_1_287/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_886 sky130_fd_sc_hd__clkinv_1_886/Y sky130_fd_sc_hd__inv_4_17/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_298 sky130_fd_sc_hd__nand2_1_298/Y sky130_fd_sc_hd__or2_0_22/X
+ sky130_fd_sc_hd__or2_0_23/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_897 sky130_fd_sc_hd__clkinv_1_897/Y sky130_fd_sc_hd__clkinv_1_897/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__conb_1_20 sky130_fd_sc_hd__conb_1_20/LO sky130_fd_sc_hd__conb_1_20/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_31 sky130_fd_sc_hd__conb_1_31/LO sky130_fd_sc_hd__conb_1_31/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1303 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_42 sky130_fd_sc_hd__conb_1_42/LO sky130_fd_sc_hd__conb_1_42/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1314 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_53 sky130_fd_sc_hd__conb_1_53/LO sky130_fd_sc_hd__conb_1_53/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1325 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_64 sky130_fd_sc_hd__conb_1_64/LO sky130_fd_sc_hd__conb_1_64/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1336 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_75 sky130_fd_sc_hd__conb_1_75/LO sky130_fd_sc_hd__conb_1_75/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1347 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_86 sky130_fd_sc_hd__conb_1_86/LO sky130_fd_sc_hd__conb_1_86/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1358 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_97 sky130_fd_sc_hd__conb_1_97/LO sky130_fd_sc_hd__conb_1_97/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1369 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__mux2_2_4 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_4/A1 sky130_fd_sc_hd__buf_2_90/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__or2_0_74/A vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__decap_12_860 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_871 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_882 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_893 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_605 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__fah_1_12/B
+ sky130_fd_sc_hd__xor2_1_605/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_616 sky130_fd_sc_hd__xor2_1_616/B sky130_fd_sc_hd__xor2_1_616/X
+ sky130_fd_sc_hd__xor2_1_616/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_627 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__or2_0_68/B
+ sky130_fd_sc_hd__xor2_1_627/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_638 sky130_fd_sc_hd__xor2_1_638/B sky130_fd_sc_hd__xor2_1_638/X
+ sky130_fd_sc_hd__xor2_1_639/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_649 sky130_fd_sc_hd__xor2_1_649/B sky130_fd_sc_hd__xor2_1_649/X
+ sky130_fd_sc_hd__xor2_1_649/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1870 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a211o_1_18 vssd1 vccd1 sky130_fd_sc_hd__fa_2_239/B sky130_fd_sc_hd__dfxtp_1_81/Q
+ sky130_fd_sc_hd__nor2_1_22/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_18/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__a211o_1_29 vssd1 vccd1 sky130_fd_sc_hd__fa_2_154/A sky130_fd_sc_hd__dfxtp_1_92/Q
+ sky130_fd_sc_hd__nor2_1_33/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_29/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__o2bb2ai_1_0 sky130_fd_sc_hd__o2bb2ai_1_0/Y sky130_fd_sc_hd__nand2_1_167/Y
+ sky130_fd_sc_hd__o21ai_1_161/Y sky130_fd_sc_hd__o21ai_1_161/Y sky130_fd_sc_hd__nand2_1_167/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__clkinv_1_105 io_oeb[34] sky130_fd_sc_hd__conb_1_37/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_116 io_oeb[23] sky130_fd_sc_hd__conb_1_26/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_127 io_oeb[12] sky130_fd_sc_hd__conb_1_15/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_138 io_oeb[1] sky130_fd_sc_hd__conb_1_4/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_149 sky130_fd_sc_hd__nor2_1_40/A sky130_fd_sc_hd__ha_2_9/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_18 sky130_fd_sc_hd__inv_2_66/Y sky130_fd_sc_hd__or2_0_86/B
+ sky130_fd_sc_hd__a22o_1_18/X sky130_fd_sc_hd__nor2_1_233/Y sky130_fd_sc_hd__a22o_1_18/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_29 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__buf_2_104/X
+ sky130_fd_sc_hd__a22o_1_29/X sky130_fd_sc_hd__a22o_1_29/B2 sky130_fd_sc_hd__inv_2_69/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__o21ai_1_5 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_5/A2 sky130_fd_sc_hd__nor2_4_4/B
+ sky130_fd_sc_hd__o21ai_1_5/B1 sky130_fd_sc_hd__ha_2_0/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2_1_210 sky130_fd_sc_hd__buf_2_15/X sky130_fd_sc_hd__nor2_1_210/Y
+ sky130_fd_sc_hd__buf_2_27/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_221 sky130_fd_sc_hd__mux2_2_35/X sky130_fd_sc_hd__nor2_1_221/Y
+ sky130_fd_sc_hd__mux2_2_15/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_232 sky130_fd_sc_hd__mux2_4_4/X sky130_fd_sc_hd__nor2_1_232/Y
+ la_data_out[68] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_243 sky130_fd_sc_hd__nor2_1_243/B sky130_fd_sc_hd__nor2_1_243/Y
+ sky130_fd_sc_hd__nor2_1_243/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_254 sky130_fd_sc_hd__nor2_1_254/B sky130_fd_sc_hd__nor2_1_254/Y
+ sky130_fd_sc_hd__nor2_1_254/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_2_8 sky130_fd_sc_hd__clkinv_4_2/A sky130_fd_sc_hd__clkinv_2_8/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__nor2_1_265 sky130_fd_sc_hd__nor2_1_265/B sky130_fd_sc_hd__nor2_1_265/Y
+ sky130_fd_sc_hd__nor2_1_265/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_276 sky130_fd_sc_hd__nor2_1_277/Y sky130_fd_sc_hd__nand3_1_5/C
+ sky130_fd_sc_hd__a21o_2_0/B1 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_450 sky130_fd_sc_hd__buf_12_450/A sky130_fd_sc_hd__buf_12_469/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_461 sky130_fd_sc_hd__buf_12_461/A sky130_fd_sc_hd__buf_12_548/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_472 sky130_fd_sc_hd__buf_12_472/A sky130_fd_sc_hd__buf_12_558/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_101 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_483 sky130_fd_sc_hd__buf_12_483/A sky130_fd_sc_hd__buf_12_508/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_112 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_494 sky130_fd_sc_hd__buf_12_494/A sky130_fd_sc_hd__buf_12_522/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_123 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_134 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_145 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_156 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_167 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_202 vssd1 vccd1 sky130_fd_sc_hd__or2_0_80/A sky130_fd_sc_hd__nor2b_1_19/A
+ sky130_fd_sc_hd__mux2_2_46/X vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_178 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_650 sky130_fd_sc_hd__xnor2_1_200/A sky130_fd_sc_hd__and2_0_284/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_213 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_213/B sky130_fd_sc_hd__or2_0_86/B
+ sky130_fd_sc_hd__xnor2_1_213/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_189 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_661 sky130_fd_sc_hd__xor2_1_652/A sky130_fd_sc_hd__o21ai_1_875/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_19 sky130_fd_sc_hd__nand2_8_0/A sky130_fd_sc_hd__nand2_1_7/B
+ sky130_fd_sc_hd__or2_1_11/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_224 vssd1 vccd1 la_data_out[77] sky130_fd_sc_hd__xnor2_1_224/Y
+ sky130_fd_sc_hd__or2_0_80/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_672 sky130_fd_sc_hd__nand2_1_743/A sky130_fd_sc_hd__nor2_1_239/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_235 vssd1 vccd1 la_data_out[77] sky130_fd_sc_hd__xnor2_1_235/Y
+ la_data_out[67] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_683 sky130_fd_sc_hd__nand2_1_758/A sky130_fd_sc_hd__nor2_1_244/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_246 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_4/B sky130_fd_sc_hd__xnor2_1_246/Y
+ sky130_fd_sc_hd__buf_4_41/X vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_694 sky130_fd_sc_hd__clkinv_1_694/Y sky130_fd_sc_hd__nand2_1_777/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_257 vssd1 vccd1 sky130_fd_sc_hd__buf_2_207/X sky130_fd_sc_hd__xnor2_1_257/Y
+ la_data_out[71] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_268 vssd1 vccd1 sky130_fd_sc_hd__or2_0_84/A sky130_fd_sc_hd__xnor2_1_268/Y
+ sky130_fd_sc_hd__or2_0_78/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_279 vssd1 vccd1 la_data_out[79] sky130_fd_sc_hd__xnor2_1_279/Y
+ sky130_fd_sc_hd__mux2_2_24/X vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_1100 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1111 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1122 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1133 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1144 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1155 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand3_1_1 sky130_fd_sc_hd__nor2_1_38/A sky130_fd_sc_hd__nand3_1_4/A
+ sky130_fd_sc_hd__nand3_1_4/C sky130_fd_sc_hd__nor2_1_39/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__decap_12_1166 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1177 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_608 vssd1 vccd1 sky130_fd_sc_hd__inv_2_34/Y sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_608/B1 sky130_fd_sc_hd__xor2_1_400/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1188 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_619 vssd1 vccd1 sky130_fd_sc_hd__buf_2_7/X sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_619/B1 sky130_fd_sc_hd__xor2_1_412/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1199 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__fah_1_6 sky130_fd_sc_hd__or2_1_2/A sky130_fd_sc_hd__fah_1_6/B sky130_fd_sc_hd__fah_1_6/A
+ sky130_fd_sc_hd__nor2_2_27/B sky130_fd_sc_hd__fah_1_6/CI vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__fah_1
Xsky130_fd_sc_hd__sdlclkp_2_13 sky130_fd_sc_hd__conb_1_145/LO sky130_fd_sc_hd__clkinv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_451/CLK sky130_fd_sc_hd__o31ai_2_0/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__a222oi_1_70 vccd1 vssd1 sky130_fd_sc_hd__and3_1_0/X sky130_fd_sc_hd__or2_0_52/B
+ sky130_fd_sc_hd__or2_0_53/A sky130_fd_sc_hd__nor2_1_56/Y sky130_fd_sc_hd__buf_2_32/X
+ sky130_fd_sc_hd__a222oi_1_70/Y sky130_fd_sc_hd__nor2b_1_3/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_81 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__or2_0_42/B
+ sky130_fd_sc_hd__or2_0_39/B sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__or2_0_58/A
+ sky130_fd_sc_hd__a222oi_1_81/Y sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_92 vccd1 vssd1 sky130_fd_sc_hd__and3_4_4/X sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__inv_6_0/Y sky130_fd_sc_hd__nor2_1_61/Y sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__a222oi_1_92/Y sky130_fd_sc_hd__nor2b_1_4/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_690 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_50 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_50/B sky130_fd_sc_hd__xnor2_1_50/Y
+ sky130_fd_sc_hd__xnor2_1_50/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_61 vssd1 vccd1 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__and3_4_3/B
+ sky130_fd_sc_hd__xnor2_1_61/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_402 sky130_fd_sc_hd__fa_2_281/A sky130_fd_sc_hd__fa_2_274/A
+ sky130_fd_sc_hd__xor2_1_402/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_72 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_72/B sky130_fd_sc_hd__xnor2_1_72/Y
+ sky130_fd_sc_hd__xnor2_1_72/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_413 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__or2_0_49/A
+ sky130_fd_sc_hd__xor2_1_413/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_83 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_83/B sky130_fd_sc_hd__xnor2_1_83/Y
+ sky130_fd_sc_hd__xnor2_1_83/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_424 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__and3_4_9/B
+ sky130_fd_sc_hd__xor2_1_424/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_94 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_344/A sky130_fd_sc_hd__and3_4_15/B
+ sky130_fd_sc_hd__xnor2_1_97/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_435 sky130_fd_sc_hd__fah_1_14/A sky130_fd_sc_hd__xor3_1_29/B
+ sky130_fd_sc_hd__xor2_1_435/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_446 sky130_fd_sc_hd__fa_2_379/A sky130_fd_sc_hd__fa_2_285/A
+ sky130_fd_sc_hd__xor2_1_446/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_457 sky130_fd_sc_hd__xor2_1_548/B sky130_fd_sc_hd__fa_2_295/A
+ sky130_fd_sc_hd__xor2_1_457/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_468 sky130_fd_sc_hd__xor2_1_468/B sky130_fd_sc_hd__inv_2_59/A
+ sky130_fd_sc_hd__xor2_1_468/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_479 sky130_fd_sc_hd__fa_2_379/A sky130_fd_sc_hd__fa_2_313/A
+ sky130_fd_sc_hd__xor2_1_479/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__o32ai_1_0 sky130_fd_sc_hd__nor2_4_3/Y sky130_fd_sc_hd__inv_2_8/A
+ sky130_fd_sc_hd__nor2_4_4/B sky130_fd_sc_hd__nor2b_1_1/Y sky130_fd_sc_hd__nor2_4_3/Y
+ sky130_fd_sc_hd__nor2_4_3/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o32ai_1
Xsky130_fd_sc_hd__decap_12_2 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_2_13 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkinv_2_13/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_24 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_12_1/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_35 sky130_fd_sc_hd__clkinv_2_35/Y sky130_fd_sc_hd__nand2_1_11/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_46 sky130_fd_sc_hd__clkinv_2_46/Y sky130_fd_sc_hd__clkinv_8_40/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_57 la_data_out[89] sky130_fd_sc_hd__clkinv_4_95/Y vccd1
+ vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__or2_1_6 sky130_fd_sc_hd__or2_1_6/A sky130_fd_sc_hd__or2_1_6/X sky130_fd_sc_hd__or2_1_6/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_1
Xsky130_fd_sc_hd__sdlclkp_4_9 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_4_0/Y
+ sky130_fd_sc_hd__dfxtp_1_105/CLK sky130_fd_sc_hd__clkbuf_1_11/X vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__buf_12_280 sky130_fd_sc_hd__buf_12_79/X sky130_fd_sc_hd__buf_12_514/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_291 sky130_fd_sc_hd__buf_12_291/A sky130_fd_sc_hd__buf_12_618/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_150 sky130_fd_sc_hd__xnor2_1_91/Y sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xnor2_1_28/Y sky130_fd_sc_hd__o21ai_1_80/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_161 sky130_fd_sc_hd__xor2_1_367/X sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xor2_1_154/X sky130_fd_sc_hd__a22oi_1_161/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_172 sky130_fd_sc_hd__nand2_1_129/A sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xnor2_1_50/Y sky130_fd_sc_hd__a22oi_1_172/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_183 sky130_fd_sc_hd__xnor2_1_120/Y sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xnor2_1_57/Y sky130_fd_sc_hd__a22oi_1_183/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_194 sky130_fd_sc_hd__clkbuf_1_3/X sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__nor2b_1_5/Y sky130_fd_sc_hd__nor2_1_68/Y sky130_fd_sc_hd__a22oi_1_194/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22o_4_3 sky130_fd_sc_hd__nand2_1_8/B sky130_fd_sc_hd__mux2_2_43/X
+ sky130_fd_sc_hd__or2_0_66/A sky130_fd_sc_hd__mux2_2_20/X sky130_fd_sc_hd__nand2_1_7/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_4
Xsky130_fd_sc_hd__clkinv_1_480 sky130_fd_sc_hd__nand2_1_436/A sky130_fd_sc_hd__nor2_1_145/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_491 sky130_fd_sc_hd__nand2_1_452/A sky130_fd_sc_hd__nor2_2_18/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_405 vssd1 vccd1 sky130_fd_sc_hd__nand2_2_12/Y sky130_fd_sc_hd__nand2b_1_10/Y
+ sky130_fd_sc_hd__a22oi_1_202/Y sky130_fd_sc_hd__xor3_1_15/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_416 vssd1 vccd1 sky130_fd_sc_hd__buf_2_11/X sky130_fd_sc_hd__nand2b_1_12/Y
+ sky130_fd_sc_hd__o21ai_1_416/B1 sky130_fd_sc_hd__xor2_1_225/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_427 vssd1 vccd1 sky130_fd_sc_hd__inv_2_32/Y sky130_fd_sc_hd__nand2b_1_14/Y
+ sky130_fd_sc_hd__o21ai_1_427/B1 sky130_fd_sc_hd__xor2_1_233/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_438 vssd1 vccd1 sky130_fd_sc_hd__inv_2_34/Y sky130_fd_sc_hd__nand2b_1_13/Y
+ sky130_fd_sc_hd__o21ai_1_438/B1 sky130_fd_sc_hd__xor2_1_243/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_449 vssd1 vccd1 sky130_fd_sc_hd__inv_2_36/Y sky130_fd_sc_hd__nand2b_1_9/Y
+ sky130_fd_sc_hd__o21ai_1_449/B1 sky130_fd_sc_hd__xor2_1_252/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2_4_14 sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__nor2_4_14/A
+ sky130_fd_sc_hd__nor2_4_14/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__nand2_1_809 sky130_fd_sc_hd__nand2_1_809/Y sky130_fd_sc_hd__nor2_1_258/A
+ sky130_fd_sc_hd__nor2_1_258/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_210 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__xor2_1_210/X
+ sky130_fd_sc_hd__xor2_1_210/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_221 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__xor3_1_19/C
+ sky130_fd_sc_hd__xor2_1_221/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_232 sky130_fd_sc_hd__fa_2_170/A sky130_fd_sc_hd__fa_2_148/B
+ sky130_fd_sc_hd__xor2_1_232/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_243 sky130_fd_sc_hd__fa_2_217/A sky130_fd_sc_hd__fa_2_155/B
+ sky130_fd_sc_hd__xor2_1_243/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_254 sky130_fd_sc_hd__fa_2_239/A sky130_fd_sc_hd__fa_2_165/B
+ sky130_fd_sc_hd__xor2_1_254/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_265 sky130_fd_sc_hd__fa_2_217/A sky130_fd_sc_hd__fa_2_173/B
+ sky130_fd_sc_hd__xor2_1_265/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_276 sky130_fd_sc_hd__xor2_1_276/B sky130_fd_sc_hd__xor2_1_276/X
+ sky130_fd_sc_hd__a21oi_2_9/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_287 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__fa_2_196/A
+ sky130_fd_sc_hd__xor2_1_287/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_298 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__fa_2_204/B
+ sky130_fd_sc_hd__xor2_1_298/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_203 vssd1 vccd1 sky130_fd_sc_hd__buf_12_14/A sky130_fd_sc_hd__clkbuf_1_51/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_214 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_214/X sky130_fd_sc_hd__buf_8_44/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_225 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_225/X sky130_fd_sc_hd__clkbuf_1_225/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_236 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_236/X sky130_fd_sc_hd__clkinv_1_875/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_307 vccd1 vssd1 sky130_fd_sc_hd__and3_4_17/X sky130_fd_sc_hd__buf_2_23/X
+ sky130_fd_sc_hd__buf_2_31/X sky130_fd_sc_hd__nor2_2_20/Y sky130_fd_sc_hd__buf_2_19/X
+ sky130_fd_sc_hd__o21ai_1_522/B1 sky130_fd_sc_hd__nor2b_2_4/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_247 vssd1 vccd1 sky130_fd_sc_hd__buf_8_80/A sky130_fd_sc_hd__clkbuf_1_303/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_318 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__buf_4_3/X sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__o21ai_1_534/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_258 vssd1 vccd1 sky130_fd_sc_hd__buf_8_71/A sky130_fd_sc_hd__clkbuf_1_258/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_2_5 sky130_fd_sc_hd__dfxtp_2_5/Q sky130_fd_sc_hd__dfxtp_2_5/CLK
+ sky130_fd_sc_hd__dfxtp_2_5/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_2
Xsky130_fd_sc_hd__a222oi_1_329 vccd1 vssd1 sky130_fd_sc_hd__and3_4_10/X sky130_fd_sc_hd__buf_4_0/X
+ sky130_fd_sc_hd__buf_2_23/X sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__buf_2_31/X
+ sky130_fd_sc_hd__o21ai_1_550/B1 sky130_fd_sc_hd__and2b_4_7/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_269 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_269/X sky130_fd_sc_hd__clkbuf_1_288/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_2_70 vccd1 vssd1 sky130_fd_sc_hd__buf_2_70/X sky130_fd_sc_hd__buf_2_70/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_81 vccd1 vssd1 sky130_fd_sc_hd__buf_2_81/X sky130_fd_sc_hd__buf_2_81/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_92 vccd1 vssd1 sky130_fd_sc_hd__buf_2_92/X sky130_fd_sc_hd__buf_2_92/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_4_8 vccd1 vssd1 sky130_fd_sc_hd__buf_4_8/X sky130_fd_sc_hd__buf_4_8/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__and2_0_201 vccd1 vssd1 sky130_fd_sc_hd__and2_0_201/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_201/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_212 vccd1 vssd1 sky130_fd_sc_hd__and2_0_212/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_73/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_223 vccd1 vssd1 sky130_fd_sc_hd__and2_0_223/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_64/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_234 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_89/D sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__o21ai_1_55/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_245 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_59/D sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__o21ai_1_46/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_256 vccd1 vssd1 sky130_fd_sc_hd__and2_0_256/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__xor2_1_650/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_267 vccd1 vssd1 sky130_fd_sc_hd__and2_0_267/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__and2_0_267/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_278 vccd1 vssd1 sky130_fd_sc_hd__and2_0_278/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__fa_2_419/SUM vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_289 vccd1 vssd1 sky130_fd_sc_hd__and2_0_289/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_10/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__a21oi_2_19 sky130_fd_sc_hd__a21oi_2_19/B1 sky130_fd_sc_hd__or2_1_3/X
+ sky130_fd_sc_hd__o21ai_2_16/Y sky130_fd_sc_hd__xor2_1_559/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_2
Xsky130_fd_sc_hd__xor3_1_10 sky130_fd_sc_hd__xor3_1_10/X sky130_fd_sc_hd__xor3_1_11/X
+ sky130_fd_sc_hd__xor3_1_10/B sky130_fd_sc_hd__xor3_1_16/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__xor3_1_21 sky130_fd_sc_hd__xor3_1_21/X sky130_fd_sc_hd__xor3_1_21/C
+ sky130_fd_sc_hd__xor3_1_22/X sky130_fd_sc_hd__xor3_1_21/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__sdlclkp_2_6 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_4_1/Y
+ sky130_fd_sc_hd__dfxtp_1_141/CLK sky130_fd_sc_hd__o21ai_1_1/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__inv_4_8 sky130_fd_sc_hd__inv_4_8/Y sky130_fd_sc_hd__inv_4_8/A vccd1
+ vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__a22o_2_0 sky130_fd_sc_hd__nand2_1_7/B sky130_fd_sc_hd__fa_2_416/B
+ sky130_fd_sc_hd__or2_0_9/B sky130_fd_sc_hd__fa_2_416/A sky130_fd_sc_hd__nand2_1_8/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_2
Xsky130_fd_sc_hd__o21ai_1_202 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_0/Y sky130_fd_sc_hd__nand2b_1_1/Y
+ sky130_fd_sc_hd__a222oi_1_76/Y sky130_fd_sc_hd__xor2_1_29/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_20 sky130_fd_sc_hd__clkbuf_4_20/X sky130_fd_sc_hd__buf_8_76/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_213 vssd1 vccd1 sky130_fd_sc_hd__nand2_4_4/Y sky130_fd_sc_hd__nand2b_1_3/Y
+ sky130_fd_sc_hd__a22oi_1_192/Y sky130_fd_sc_hd__xor2_1_38/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_31 sky130_fd_sc_hd__clkinv_4_43/A sky130_fd_sc_hd__clkbuf_4_31/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_224 vssd1 vccd1 sky130_fd_sc_hd__inv_2_26/Y sky130_fd_sc_hd__nand2b_1_3/Y
+ sky130_fd_sc_hd__nand2_1_153/Y sky130_fd_sc_hd__xor2_1_48/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_42 la_data_out[57] sky130_fd_sc_hd__dfxtp_1_472/Q vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_235 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_261/A2 sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__o21ai_1_235/B1 sky130_fd_sc_hd__xor2_1_60/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_246 vssd1 vccd1 sky130_fd_sc_hd__nand2_4_4/Y sky130_fd_sc_hd__nand2b_1_4/Y
+ sky130_fd_sc_hd__a22oi_1_193/Y sky130_fd_sc_hd__xor2_1_69/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_257 vssd1 vccd1 sky130_fd_sc_hd__inv_2_21/Y sky130_fd_sc_hd__nand2b_2_0/Y
+ sky130_fd_sc_hd__o21ai_1_257/B1 sky130_fd_sc_hd__xor2_1_80/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_268 vssd1 vccd1 sky130_fd_sc_hd__buf_2_2/X sky130_fd_sc_hd__nand2b_1_5/Y
+ sky130_fd_sc_hd__o21ai_1_268/B1 sky130_fd_sc_hd__xor2_1_90/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_279 vssd1 vccd1 sky130_fd_sc_hd__inv_2_10/Y sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__o21ai_1_279/B1 sky130_fd_sc_hd__xor2_1_101/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nand2_1_606 sky130_fd_sc_hd__nand2_1_606/Y sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__nor2_1_85/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_617 sky130_fd_sc_hd__xor2_1_602/B sky130_fd_sc_hd__nand2_1_618/Y
+ sky130_fd_sc_hd__nand2_1_617/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_628 sky130_fd_sc_hd__nand2_1_628/Y sky130_fd_sc_hd__nor2_1_209/A
+ sky130_fd_sc_hd__nor2_1_209/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_639 sky130_fd_sc_hd__nand2_1_639/Y sky130_fd_sc_hd__buf_2_24/X
+ sky130_fd_sc_hd__buf_2_26/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_402 sky130_fd_sc_hd__dfxtp_1_402/Q sky130_fd_sc_hd__clkinv_4_8/Y
+ sky130_fd_sc_hd__nor2b_1_113/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_413 sky130_fd_sc_hd__dfxtp_1_413/Q sky130_fd_sc_hd__dfxtp_1_417/CLK
+ sky130_fd_sc_hd__nor2b_1_102/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_424 sky130_fd_sc_hd__dfxtp_1_424/Q sky130_fd_sc_hd__dfxtp_1_427/CLK
+ sky130_fd_sc_hd__nor2b_1_91/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_435 sky130_fd_sc_hd__dfxtp_1_435/Q sky130_fd_sc_hd__dfxtp_1_439/CLK
+ sky130_fd_sc_hd__nor2b_1_112/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_446 sky130_fd_sc_hd__dfxtp_1_446/Q sky130_fd_sc_hd__dfxtp_1_446/CLK
+ sky130_fd_sc_hd__nor2b_1_101/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_457 sky130_fd_sc_hd__dfxtp_1_457/Q sky130_fd_sc_hd__dfxtp_1_459/CLK
+ sky130_fd_sc_hd__nor2b_1_90/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_468 sky130_fd_sc_hd__ha_2_52/A sky130_fd_sc_hd__dfxtp_1_515/CLK
+ sky130_fd_sc_hd__and2_0_358/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_479 sky130_fd_sc_hd__ha_2_19/A sky130_fd_sc_hd__dfxtp_1_479/CLK
+ sky130_fd_sc_hd__and2_0_384/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a222oi_1_104 vccd1 vssd1 sky130_fd_sc_hd__and3_4_2/X sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__buf_4_2/X sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__o21ai_1_236/B1 sky130_fd_sc_hd__and2b_4_4/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2b_1_16 sky130_fd_sc_hd__nand2b_1_16/Y sky130_fd_sc_hd__nor2_2_32/A
+ sky130_fd_sc_hd__nor2_2_32/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a222oi_1_115 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__or2_0_60/B sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__or2_0_60/A
+ sky130_fd_sc_hd__o21ai_1_251/B1 sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2b_1_27 sky130_fd_sc_hd__nand2b_1_27/Y sky130_fd_sc_hd__or2_0_84/A
+ sky130_fd_sc_hd__or2_0_79/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a222oi_1_126 vccd1 vssd1 sky130_fd_sc_hd__and3_4_1/X sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__nor2_1_85/B sky130_fd_sc_hd__nor2_2_9/Y sky130_fd_sc_hd__nor2_2_10/B
+ sky130_fd_sc_hd__o21ai_1_266/B1 sky130_fd_sc_hd__and2b_4_3/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_137 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__buf_4_4/X sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__o21ai_1_279/B1 sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_148 vccd1 vssd1 sky130_fd_sc_hd__and3_4_6/X sky130_fd_sc_hd__clkbuf_1_3/X
+ sky130_fd_sc_hd__or2_0_53/A sky130_fd_sc_hd__nor2_1_72/Y sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__o21ai_1_293/B1 sky130_fd_sc_hd__nor2b_1_6/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__o21ai_1_780 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_780/A2 sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_780/B1 sky130_fd_sc_hd__xor2_1_554/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_159 vccd1 vssd1 sky130_fd_sc_hd__and3_4_1/X sky130_fd_sc_hd__nor2_2_5/B
+ sky130_fd_sc_hd__nor2_2_4/B sky130_fd_sc_hd__nor2_2_9/Y sky130_fd_sc_hd__buf_2_4/X
+ sky130_fd_sc_hd__o21ai_1_307/B1 sky130_fd_sc_hd__and2b_4_3/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_307 sky130_fd_sc_hd__fa_2_299/B sky130_fd_sc_hd__fa_2_307/SUM
+ sky130_fd_sc_hd__fa_2_307/A sky130_fd_sc_hd__fa_2_307/B sky130_fd_sc_hd__fa_2_308/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o21ai_1_791 vssd1 vccd1 sky130_fd_sc_hd__inv_2_48/Y sky130_fd_sc_hd__nand2b_1_16/Y
+ sky130_fd_sc_hd__o21ai_1_791/B1 sky130_fd_sc_hd__xor2_1_565/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_318 sky130_fd_sc_hd__fa_2_316/CIN sky130_fd_sc_hd__fa_2_324/B
+ sky130_fd_sc_hd__fa_2_318/A sky130_fd_sc_hd__fa_2_318/B sky130_fd_sc_hd__xor2_1_487/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_329 sky130_fd_sc_hd__fa_2_325/B sky130_fd_sc_hd__fa_2_333/CIN
+ sky130_fd_sc_hd__fa_2_329/A sky130_fd_sc_hd__fa_2_329/B sky130_fd_sc_hd__fa_2_329/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_8_12 sky130_fd_sc_hd__clkinv_8_12/Y sky130_fd_sc_hd__clkinv_8_12/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_23 sky130_fd_sc_hd__clkinv_8_25/A sky130_fd_sc_hd__clkinv_8_23/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_34 sky130_fd_sc_hd__clkinv_8_35/A sky130_fd_sc_hd__clkinv_8_34/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_45 sky130_fd_sc_hd__clkinv_8_46/A sky130_fd_sc_hd__clkinv_8_45/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_56 sky130_fd_sc_hd__clkinv_8_7/A sky130_fd_sc_hd__clkinv_8_56/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_10 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__buf_12_78/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_8_67 sky130_fd_sc_hd__clkinv_8_68/A sky130_fd_sc_hd__clkinv_8_67/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_21 sky130_fd_sc_hd__buf_12_21/A sky130_fd_sc_hd__buf_12_21/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_8_78 sky130_fd_sc_hd__clkinv_8_79/A sky130_fd_sc_hd__clkinv_8_78/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_32 sky130_fd_sc_hd__inv_2_90/Y sky130_fd_sc_hd__buf_12_32/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_8_89 sky130_fd_sc_hd__dfxtp_1_3/CLK sky130_fd_sc_hd__clkinv_8_89/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_43 sky130_fd_sc_hd__buf_12_43/A sky130_fd_sc_hd__buf_12_43/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_54 sky130_fd_sc_hd__buf_12_54/A sky130_fd_sc_hd__buf_12_54/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_65 sky130_fd_sc_hd__buf_12_65/A sky130_fd_sc_hd__buf_12_65/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_76 sky130_fd_sc_hd__buf_8_58/X sky130_fd_sc_hd__buf_12_76/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_87 sky130_fd_sc_hd__buf_8_122/X sky130_fd_sc_hd__buf_12_87/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_98 sky130_fd_sc_hd__buf_8_43/X sky130_fd_sc_hd__buf_12_98/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_2_5 vccd1 vssd1 sky130_fd_sc_hd__buf_2_5/X sky130_fd_sc_hd__buf_2_5/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__inv_2_5 sky130_fd_sc_hd__inv_2_5/A sky130_fd_sc_hd__inv_2_5/Y vccd1
+ vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__nor2_1_15 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_15/Y
+ sky130_fd_sc_hd__nor2_1_15/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_26 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_26/Y
+ sky130_fd_sc_hd__nor2_1_26/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_37 sky130_fd_sc_hd__nor2_4_7/B sky130_fd_sc_hd__nor2_1_37/Y
+ sky130_fd_sc_hd__nor2_1_37/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_48 sky130_fd_sc_hd__xnor2_1_8/Y sky130_fd_sc_hd__nor2_1_48/Y
+ sky130_fd_sc_hd__xnor2_1_5/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_59 sky130_fd_sc_hd__nor2_1_59/B sky130_fd_sc_hd__nor2_1_59/Y
+ sky130_fd_sc_hd__nor2_1_59/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_12_508 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_519 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__and2_0_70 vccd1 vssd1 sky130_fd_sc_hd__and2_0_70/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__or2_0_60/B vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_403 sky130_fd_sc_hd__xnor2_1_95/A sky130_fd_sc_hd__nand2_1_404/Y
+ sky130_fd_sc_hd__or2_0_35/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_81 vccd1 vssd1 sky130_fd_sc_hd__and2_0_81/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__buf_6_0/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_414 sky130_fd_sc_hd__xnor2_1_98/A sky130_fd_sc_hd__nand2_1_415/Y
+ sky130_fd_sc_hd__or2_0_37/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_92 vccd1 vssd1 sky130_fd_sc_hd__and2_0_92/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__or2_0_58/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_425 sky130_fd_sc_hd__xor2_1_367/B sky130_fd_sc_hd__nand2_1_426/Y
+ sky130_fd_sc_hd__nand2_1_425/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_436 sky130_fd_sc_hd__xnor2_1_107/A sky130_fd_sc_hd__nand2_1_437/Y
+ sky130_fd_sc_hd__nand2_1_436/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_447 sky130_fd_sc_hd__nand2_1_447/Y sky130_fd_sc_hd__nor2_1_149/A
+ sky130_fd_sc_hd__nor2_1_149/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_458 sky130_fd_sc_hd__xnor2_1_115/A sky130_fd_sc_hd__nand2_1_459/Y
+ sky130_fd_sc_hd__nand2_1_458/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_469 sky130_fd_sc_hd__nand2_1_469/Y sky130_fd_sc_hd__or2_0_50/X
+ sky130_fd_sc_hd__or2_0_49/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_16 sky130_fd_sc_hd__and3_4_24/C sky130_fd_sc_hd__nor2b_1_16/Y
+ sky130_fd_sc_hd__and3_4_24/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_27 sky130_fd_sc_hd__fa_2_415/A sky130_fd_sc_hd__nor2b_1_27/Y
+ sky130_fd_sc_hd__buf_2_214/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_38 sky130_fd_sc_hd__mux2_2_35/X sky130_fd_sc_hd__fa_2_470/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1005 sky130_fd_sc_hd__clkinv_1_1005/Y sky130_fd_sc_hd__clkinv_1_1005/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_49 sky130_fd_sc_hd__or2_0_76/B sky130_fd_sc_hd__nor2b_1_49/Y
+ sky130_fd_sc_hd__buf_2_214/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1016 sky130_fd_sc_hd__clkinv_1_1017/A sky130_fd_sc_hd__buf_6_6/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1027 sky130_fd_sc_hd__clkinv_1_1028/A sky130_fd_sc_hd__inv_4_9/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1038 sky130_fd_sc_hd__clkbuf_8_1/A sky130_fd_sc_hd__clkinv_1_1038/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_80 sky130_fd_sc_hd__buf_8_80/A sky130_fd_sc_hd__buf_8_80/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__clkinv_1_1049 sky130_fd_sc_hd__inv_2_182/A sky130_fd_sc_hd__clkbuf_1_235/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_91 sky130_fd_sc_hd__buf_8_91/A sky130_fd_sc_hd__buf_8_91/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__decap_12_1507 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_210 sky130_fd_sc_hd__xnor2_1_147/A sky130_fd_sc_hd__dfxtp_2_0/CLK
+ sky130_fd_sc_hd__and2_0_61/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1518 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_221 sky130_fd_sc_hd__xor2_1_418/A sky130_fd_sc_hd__dfxtp_1_234/CLK
+ sky130_fd_sc_hd__and2_0_17/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1529 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_232 sky130_fd_sc_hd__xor2_1_362/B sky130_fd_sc_hd__dfxtp_1_234/CLK
+ sky130_fd_sc_hd__and2_0_44/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_243 sky130_fd_sc_hd__xor2_1_262/A sky130_fd_sc_hd__clkinv_4_4/Y
+ sky130_fd_sc_hd__and2_0_92/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_254 sky130_fd_sc_hd__xor2_1_183/A sky130_fd_sc_hd__clkinv_4_6/Y
+ sky130_fd_sc_hd__and2_0_52/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_265 sky130_fd_sc_hd__xnor2_1_27/A sky130_fd_sc_hd__dfxtp_1_266/CLK
+ sky130_fd_sc_hd__and2_0_82/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_276 sky130_fd_sc_hd__dfxtp_1_276/Q sky130_fd_sc_hd__dfxtp_1_2/CLK
+ sky130_fd_sc_hd__and2_0_252/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_287 sky130_fd_sc_hd__a22oi_1_8/B2 sky130_fd_sc_hd__dfxtp_1_2/CLK
+ sky130_fd_sc_hd__and2_0_263/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_298 sky130_fd_sc_hd__dfxtp_1_298/Q sky130_fd_sc_hd__clkinv_8_6/Y
+ sky130_fd_sc_hd__and2_0_274/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o22ai_1_7 sky130_fd_sc_hd__o22ai_1_7/A2 sky130_fd_sc_hd__o22ai_1_7/B1
+ sky130_fd_sc_hd__o22ai_1_7/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__o22ai_1_9/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_104 sky130_fd_sc_hd__fa_2_102/B sky130_fd_sc_hd__fa_2_105/A
+ sky130_fd_sc_hd__fa_2_104/A sky130_fd_sc_hd__fa_2_104/B sky130_fd_sc_hd__fa_2_104/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_115 sky130_fd_sc_hd__nor2_1_43/A sky130_fd_sc_hd__nor2_1_80/B
+ sky130_fd_sc_hd__fa_2_115/A sky130_fd_sc_hd__fa_2_115/B sky130_fd_sc_hd__fa_2_115/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_126 sky130_fd_sc_hd__nor2_1_86/A sky130_fd_sc_hd__nor2_1_88/B
+ sky130_fd_sc_hd__fa_2_126/A sky130_fd_sc_hd__fa_2_126/B sky130_fd_sc_hd__fa_2_126/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_137 sky130_fd_sc_hd__fa_2_135/CIN sky130_fd_sc_hd__fa_2_138/A
+ sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__fa_2_137/B sky130_fd_sc_hd__xor2_1_196/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_148 sky130_fd_sc_hd__xor3_1_18/A sky130_fd_sc_hd__fa_2_145/B
+ sky130_fd_sc_hd__ha_2_1/SUM sky130_fd_sc_hd__fa_2_148/B sky130_fd_sc_hd__fa_2_148/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_159 sky130_fd_sc_hd__or2_0_27/A sky130_fd_sc_hd__nor2_1_110/A
+ sky130_fd_sc_hd__fa_2_159/A sky130_fd_sc_hd__fa_2_159/B sky130_fd_sc_hd__fa_2_159/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and3_4_9 sky130_fd_sc_hd__and3_4_9/A sky130_fd_sc_hd__and3_4_9/B
+ sky130_fd_sc_hd__or2b_2_1/A sky130_fd_sc_hd__and3_4_9/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__buf_2_110 vccd1 vssd1 sky130_fd_sc_hd__buf_2_110/X sky130_fd_sc_hd__buf_2_110/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_121 vccd1 vssd1 sky130_fd_sc_hd__buf_2_121/X sky130_fd_sc_hd__buf_2_121/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_14 sky130_fd_sc_hd__o22ai_1_49/B1 sky130_fd_sc_hd__o22ai_1_14/B1
+ sky130_fd_sc_hd__o22ai_1_14/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__o22ai_1_9/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_132 vccd1 vssd1 sky130_fd_sc_hd__buf_2_132/X sky130_fd_sc_hd__inv_2_4/Y
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_25 sky130_fd_sc_hd__o22ai_1_37/B1 sky130_fd_sc_hd__o21ai_1_7/A2
+ sky130_fd_sc_hd__o22ai_1_25/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__inv_4_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_143 vccd1 vssd1 sky130_fd_sc_hd__buf_2_143/X sky130_fd_sc_hd__buf_2_143/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_36 sky130_fd_sc_hd__nor2_1_30/A sky130_fd_sc_hd__o22ai_1_36/B1
+ sky130_fd_sc_hd__o22ai_1_36/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_154 vccd1 vssd1 sky130_fd_sc_hd__buf_2_154/X sky130_fd_sc_hd__buf_2_154/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_47 sky130_fd_sc_hd__nor2_1_20/A sky130_fd_sc_hd__o22ai_1_47/B1
+ sky130_fd_sc_hd__o22ai_1_47/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_165 vccd1 vssd1 sky130_fd_sc_hd__buf_2_165/X sky130_fd_sc_hd__buf_2_165/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_58 sky130_fd_sc_hd__nor2_1_9/A sky130_fd_sc_hd__o22ai_1_5/A2
+ sky130_fd_sc_hd__o22ai_1_58/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_176 vccd1 vssd1 la_data_out[64] sky130_fd_sc_hd__ha_2_19/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_69 sky130_fd_sc_hd__xnor2_2_4/Y sky130_fd_sc_hd__xnor2_1_228/Y
+ sky130_fd_sc_hd__o22ai_1_69/Y sky130_fd_sc_hd__xnor2_1_220/Y sky130_fd_sc_hd__o22ai_1_96/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_187 vccd1 vssd1 sky130_fd_sc_hd__buf_2_43/A sky130_fd_sc_hd__buf_2_42/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_198 vccd1 vssd1 la_data_out[95] sky130_fd_sc_hd__nand2_2_3/Y
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_4_16 vccd1 vssd1 sky130_fd_sc_hd__buf_4_16/X sky130_fd_sc_hd__buf_4_16/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_27 vccd1 vssd1 sky130_fd_sc_hd__buf_4_27/X sky130_fd_sc_hd__buf_8_57/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_38 vccd1 vssd1 sky130_fd_sc_hd__buf_4_38/X sky130_fd_sc_hd__buf_4_38/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__clkbuf_1_10 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_10/X sky130_fd_sc_hd__xnor2_1_126/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_21 vssd1 vccd1 sky130_fd_sc_hd__or2_0_39/B sky130_fd_sc_hd__or2_0_58/B
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_109 sky130_fd_sc_hd__buf_8_138/X sky130_fd_sc_hd__buf_12_456/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a222oi_1_490 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__nor2_1_73/B sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__o21ai_1_780/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_32 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_32/X sky130_fd_sc_hd__nor2_4_19/B
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_43 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_43/X sky130_fd_sc_hd__clkbuf_1_43/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_54 vssd1 vccd1 sky130_fd_sc_hd__buf_12_29/A sky130_fd_sc_hd__conb_1_147/HI
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_65 vssd1 vccd1 sky130_fd_sc_hd__buf_8_48/A sky130_fd_sc_hd__inv_2_150/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_76 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_20/A1 sky130_fd_sc_hd__clkbuf_1_76/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_87 vssd1 vccd1 sky130_fd_sc_hd__mux2_4_0/A1 sky130_fd_sc_hd__clkbuf_1_87/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_98 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_43/A1 sky130_fd_sc_hd__clkbuf_1_98/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkinv_1_309 sky130_fd_sc_hd__nand2_1_287/A sky130_fd_sc_hd__nor2_2_4/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__or2_0_12 sky130_fd_sc_hd__or2_0_58/A sky130_fd_sc_hd__or2_0_12/X
+ sky130_fd_sc_hd__or2_0_58/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_23 sky130_fd_sc_hd__or2_0_23/A sky130_fd_sc_hd__or2_0_23/X
+ sky130_fd_sc_hd__or2_0_23/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_34 sky130_fd_sc_hd__or2_0_34/A sky130_fd_sc_hd__or2_0_34/X
+ sky130_fd_sc_hd__or2_0_34/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_45 sky130_fd_sc_hd__buf_4_2/X sky130_fd_sc_hd__or2_0_45/X
+ sky130_fd_sc_hd__buf_4_4/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_56 sky130_fd_sc_hd__or2_0_9/A sky130_fd_sc_hd__or2_0_56/X
+ sky130_fd_sc_hd__or2_0_9/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_67 sky130_fd_sc_hd__or2_0_67/A sky130_fd_sc_hd__or2_0_67/X
+ sky130_fd_sc_hd__or2_0_67/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_78 sky130_fd_sc_hd__or2_0_78/A sky130_fd_sc_hd__or2_0_78/X
+ sky130_fd_sc_hd__or2_0_78/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_89 sky130_fd_sc_hd__or2_0_89/A sky130_fd_sc_hd__or2_0_89/X
+ sky130_fd_sc_hd__or2_0_89/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__buf_12_610 sky130_fd_sc_hd__buf_12_610/A sky130_fd_sc_hd__buf_12_610/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_621 sky130_fd_sc_hd__buf_12_621/A sky130_fd_sc_hd__buf_12_621/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_632 sky130_fd_sc_hd__buf_12_632/A sky130_fd_sc_hd__buf_12_632/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_4_103 sky130_fd_sc_hd__clkinv_2_11/A sky130_fd_sc_hd__clkinv_8_6/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_12_643 sky130_fd_sc_hd__buf_12_643/A sky130_fd_sc_hd__buf_12_643/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_4_114 sky130_fd_sc_hd__clkinv_4_114/A sky130_fd_sc_hd__clkinv_4_115/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_12_654 sky130_fd_sc_hd__buf_12_654/A sky130_fd_sc_hd__buf_12_654/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_665 sky130_fd_sc_hd__buf_12_665/A sky130_fd_sc_hd__buf_12_665/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_676 sky130_fd_sc_hd__buf_12_676/A sky130_fd_sc_hd__buf_12_676/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_305 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_316 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_200 sky130_fd_sc_hd__nand2_1_200/Y sky130_fd_sc_hd__or2_0_60/A
+ sky130_fd_sc_hd__or2_0_61/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_327 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_211 sky130_fd_sc_hd__nand2_1_211/Y sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__or2_0_60/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_338 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_810 sky130_fd_sc_hd__clkinv_1_810/Y sky130_fd_sc_hd__nand2_1_799/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_222 sky130_fd_sc_hd__xnor2_1_28/A sky130_fd_sc_hd__nand2_1_223/Y
+ sky130_fd_sc_hd__or2_0_7/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_349 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_821 sky130_fd_sc_hd__nand2_1_820/A sky130_fd_sc_hd__nor2_1_261/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_233 sky130_fd_sc_hd__nand2_1_233/Y sky130_fd_sc_hd__or2_0_8/A
+ sky130_fd_sc_hd__or2_0_8/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_832 sky130_fd_sc_hd__nand2_1_840/A sky130_fd_sc_hd__nor2_1_266/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_244 sky130_fd_sc_hd__nand2_1_244/Y sky130_fd_sc_hd__or2_0_11/A
+ sky130_fd_sc_hd__or2_0_11/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_843 sky130_fd_sc_hd__inv_2_84/A sky130_fd_sc_hd__clkbuf_1_35/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_255 sky130_fd_sc_hd__nand2_1_255/Y sky130_fd_sc_hd__nor2_1_80/A
+ sky130_fd_sc_hd__nor2_1_80/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_854 sky130_fd_sc_hd__clkinv_1_854/Y sky130_fd_sc_hd__clkinv_8_9/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_266 sky130_fd_sc_hd__nand2_1_266/Y sky130_fd_sc_hd__nor2_1_86/A
+ sky130_fd_sc_hd__nor2_1_86/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_865 sky130_fd_sc_hd__clkinv_1_865/Y sky130_fd_sc_hd__clkinv_4_81/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_277 sky130_fd_sc_hd__xnor2_1_49/A sky130_fd_sc_hd__nand2_1_278/Y
+ sky130_fd_sc_hd__nand2_1_277/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_876 sky130_fd_sc_hd__clkinv_1_876/Y sky130_fd_sc_hd__buf_4_42/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_288 sky130_fd_sc_hd__nand2_1_288/Y sky130_fd_sc_hd__nor2_2_5/B
+ sky130_fd_sc_hd__nor2_2_4/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_887 sky130_fd_sc_hd__clkinv_1_887/Y sky130_fd_sc_hd__inv_4_18/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_299 sky130_fd_sc_hd__xor2_1_199/B sky130_fd_sc_hd__nand2_1_300/Y
+ sky130_fd_sc_hd__or2_0_23/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_898 sky130_fd_sc_hd__clkinv_1_898/Y sky130_fd_sc_hd__clkinv_4_89/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__conb_1_10 sky130_fd_sc_hd__conb_1_10/LO sky130_fd_sc_hd__conb_1_10/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_21 sky130_fd_sc_hd__conb_1_21/LO sky130_fd_sc_hd__conb_1_21/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_32 sky130_fd_sc_hd__conb_1_32/LO sky130_fd_sc_hd__conb_1_32/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1304 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_43 sky130_fd_sc_hd__conb_1_43/LO sky130_fd_sc_hd__conb_1_43/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1315 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_54 sky130_fd_sc_hd__conb_1_54/LO sky130_fd_sc_hd__conb_1_54/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1326 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_65 sky130_fd_sc_hd__conb_1_65/LO sky130_fd_sc_hd__conb_1_65/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1337 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_76 sky130_fd_sc_hd__conb_1_76/LO sky130_fd_sc_hd__conb_1_76/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1348 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_87 sky130_fd_sc_hd__conb_1_87/LO sky130_fd_sc_hd__conb_1_87/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1359 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_98 sky130_fd_sc_hd__conb_1_98/LO sky130_fd_sc_hd__conb_1_98/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__mux2_2_5 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_5/A1 sky130_fd_sc_hd__buf_2_92/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__or2_0_75/A vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__decap_12_850 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_861 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_872 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_883 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_894 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_606 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__fa_2_403/B
+ sky130_fd_sc_hd__xor2_1_606/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_617 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__xor2_1_617/X
+ sky130_fd_sc_hd__xor2_1_617/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_628 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__fa_2_413/B
+ sky130_fd_sc_hd__xor2_1_628/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_639 sky130_fd_sc_hd__mux2_2_0/X sky130_fd_sc_hd__xor2_1_639/X
+ sky130_fd_sc_hd__buf_2_214/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1860 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1871 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a211o_1_19 vssd1 vccd1 sky130_fd_sc_hd__fa_2_232/A sky130_fd_sc_hd__dfxtp_1_82/Q
+ sky130_fd_sc_hd__nor2_1_23/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_19/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__o2bb2ai_1_1 sky130_fd_sc_hd__maj3_1_1/C sky130_fd_sc_hd__a21oi_1_192/Y
+ sky130_fd_sc_hd__xnor2_1_306/B sky130_fd_sc_hd__ha_2_32/A sky130_fd_sc_hd__ha_2_48/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__fa_2_490 sky130_fd_sc_hd__nor2_1_264/B sky130_fd_sc_hd__or2_0_110/A
+ sky130_fd_sc_hd__fa_2_490/A sky130_fd_sc_hd__fa_2_490/B sky130_fd_sc_hd__nor2b_1_79/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_1_106 io_oeb[33] sky130_fd_sc_hd__conb_1_36/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_117 io_oeb[22] sky130_fd_sc_hd__conb_1_25/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_128 io_oeb[11] sky130_fd_sc_hd__conb_1_14/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_139 io_oeb[0] sky130_fd_sc_hd__conb_1_3/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor3b_1_0 sky130_fd_sc_hd__buf_2_16/A sky130_fd_sc_hd__nor3b_1_0/Y
+ sky130_fd_sc_hd__ha_2_5/A sky130_fd_sc_hd__nor3b_1_0/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor3b_1
Xsky130_fd_sc_hd__a22o_1_19 sky130_fd_sc_hd__inv_2_66/Y sky130_fd_sc_hd__or2_0_87/B
+ sky130_fd_sc_hd__a22o_1_19/X sky130_fd_sc_hd__nor2_1_233/Y sky130_fd_sc_hd__xor2_1_653/X
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__o21ai_1_6 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_6/A2 sky130_fd_sc_hd__nor2_4_4/B
+ sky130_fd_sc_hd__o21ai_1_6/B1 sky130_fd_sc_hd__fa_2_37/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2_1_200 sky130_fd_sc_hd__nor2_1_200/B sky130_fd_sc_hd__nor2_1_200/Y
+ sky130_fd_sc_hd__nor2_1_200/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_211 sky130_fd_sc_hd__nor2_1_211/B sky130_fd_sc_hd__nor2_1_211/Y
+ sky130_fd_sc_hd__nor2_1_211/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_222 sky130_fd_sc_hd__mux2_2_43/X sky130_fd_sc_hd__nor2_1_222/Y
+ sky130_fd_sc_hd__mux2_2_20/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_233 sky130_fd_sc_hd__nor2_1_233/B sky130_fd_sc_hd__nor2_1_233/Y
+ sky130_fd_sc_hd__nor3_1_1/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_244 sky130_fd_sc_hd__nor2_1_244/B sky130_fd_sc_hd__nor2_1_244/Y
+ sky130_fd_sc_hd__nor2_1_244/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_255 sky130_fd_sc_hd__nor2_1_255/B sky130_fd_sc_hd__nor2_1_255/Y
+ sky130_fd_sc_hd__nor2_1_255/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_2_9 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkinv_2_9/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__nor2_1_266 sky130_fd_sc_hd__ha_2_18/SUM sky130_fd_sc_hd__nor2_1_266/Y
+ sky130_fd_sc_hd__nor2b_1_86/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_277 sky130_fd_sc_hd__nor2_1_277/B sky130_fd_sc_hd__nor2_1_277/Y
+ la_data_out[35] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_440 sky130_fd_sc_hd__buf_12_97/X sky130_fd_sc_hd__buf_12_465/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_451 sky130_fd_sc_hd__buf_12_91/X sky130_fd_sc_hd__buf_12_549/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_462 sky130_fd_sc_hd__buf_12_462/A sky130_fd_sc_hd__buf_12_565/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_473 sky130_fd_sc_hd__buf_12_473/A sky130_fd_sc_hd__buf_12_556/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_102 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_484 sky130_fd_sc_hd__buf_12_484/A sky130_fd_sc_hd__buf_12_511/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_113 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_495 sky130_fd_sc_hd__buf_12_495/A sky130_fd_sc_hd__buf_12_495/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_124 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_135 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_146 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_157 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_168 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_640 sky130_fd_sc_hd__nand2_1_692/A sky130_fd_sc_hd__nor2_1_228/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_203 vssd1 vccd1 sky130_fd_sc_hd__or2_0_79/A sky130_fd_sc_hd__nor2b_1_24/A
+ sky130_fd_sc_hd__mux2_2_38/X vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_179 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_651 sky130_fd_sc_hd__nor2_1_233/B sky130_fd_sc_hd__and2_0_1/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_214 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_214/B sky130_fd_sc_hd__nor2_1_237/B
+ sky130_fd_sc_hd__xnor2_1_214/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_662 sky130_fd_sc_hd__clkinv_1_662/Y sky130_fd_sc_hd__nand2_1_729/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_225 vssd1 vccd1 la_data_out[85] sky130_fd_sc_hd__xnor2_1_225/Y
+ sky130_fd_sc_hd__or2_0_84/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_673 sky130_fd_sc_hd__clkinv_1_673/Y sky130_fd_sc_hd__nand2_1_746/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_236 vssd1 vccd1 la_data_out[77] sky130_fd_sc_hd__xnor2_1_236/Y
+ la_data_out[68] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_684 sky130_fd_sc_hd__nand2_1_759/A sky130_fd_sc_hd__nor2_1_246/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_247 vssd1 vccd1 la_data_out[77] sky130_fd_sc_hd__xnor2_1_247/Y
+ sky130_fd_sc_hd__buf_4_41/X vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_695 sky130_fd_sc_hd__clkinv_1_695/Y sky130_fd_sc_hd__nand2_1_778/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_258 vssd1 vccd1 la_data_out[67] sky130_fd_sc_hd__xnor2_1_258/Y
+ sky130_fd_sc_hd__or2_0_79/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_269 vssd1 vccd1 la_data_out[79] sky130_fd_sc_hd__xnor2_1_269/Y
+ sky130_fd_sc_hd__or2_0_79/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_1101 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1112 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1123 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1134 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1145 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1156 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand3_1_2 sky130_fd_sc_hd__nor2_1_39/A sky130_fd_sc_hd__nand3_1_2/A
+ sky130_fd_sc_hd__nor2_1_40/Y sky130_fd_sc_hd__nor3_1_0/B vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__decap_12_1167 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1178 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_609 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_63/A sky130_fd_sc_hd__nor2_2_17/Y
+ sky130_fd_sc_hd__nand2_1_463/Y sky130_fd_sc_hd__xnor2_1_115/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1189 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__fah_1_7 sky130_fd_sc_hd__nor2_2_25/A sky130_fd_sc_hd__fah_1_7/B
+ sky130_fd_sc_hd__fah_1_7/A sky130_fd_sc_hd__or2_1_2/B sky130_fd_sc_hd__fah_1_7/CI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__fah_1
Xsky130_fd_sc_hd__sdlclkp_2_14 sky130_fd_sc_hd__conb_1_148/LO sky130_fd_sc_hd__clkinv_2_47/Y
+ sky130_fd_sc_hd__dfxtp_1_479/CLK sky130_fd_sc_hd__o21ai_1_909/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__a222oi_1_60 vccd1 vssd1 sky130_fd_sc_hd__and3_4_4/X sky130_fd_sc_hd__buf_4_6/X
+ sky130_fd_sc_hd__buf_4_1/X sky130_fd_sc_hd__nor2_1_61/Y sky130_fd_sc_hd__nor2_2_5/A
+ sky130_fd_sc_hd__a222oi_1_60/Y sky130_fd_sc_hd__nor2b_1_4/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_71 vccd1 vssd1 sky130_fd_sc_hd__and3_4_4/X sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__buf_4_6/X sky130_fd_sc_hd__nor2_1_61/Y sky130_fd_sc_hd__buf_4_1/X
+ sky130_fd_sc_hd__a222oi_1_71/Y sky130_fd_sc_hd__nor2b_1_4/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_82 vccd1 vssd1 sky130_fd_sc_hd__and3_4_1/X sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__buf_4_3/X sky130_fd_sc_hd__nor2_2_9/Y sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__a222oi_1_82/Y sky130_fd_sc_hd__and2b_4_3/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_93 vccd1 vssd1 sky130_fd_sc_hd__and3_4_7/X sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__buf_6_1/X sky130_fd_sc_hd__nor2_2_7/Y sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__a222oi_1_93/Y sky130_fd_sc_hd__nor2b_2_1/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__xnor2_1_40 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_40/B sky130_fd_sc_hd__inv_2_13/A
+ sky130_fd_sc_hd__xnor2_1_40/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_680 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_691 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_51 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__nor2_2_9/A
+ sky130_fd_sc_hd__xnor2_1_51/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_62 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_211/X sky130_fd_sc_hd__xnor2_1_62/Y
+ sky130_fd_sc_hd__xnor2_1_62/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_403 sky130_fd_sc_hd__xor2_1_403/B sky130_fd_sc_hd__xor2_1_403/X
+ sky130_fd_sc_hd__xor2_1_403/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_73 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_73/B sky130_fd_sc_hd__xnor2_1_73/Y
+ sky130_fd_sc_hd__xnor2_1_73/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_414 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__or2_0_50/B
+ sky130_fd_sc_hd__xor2_1_414/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_84 vssd1 vccd1 sky130_fd_sc_hd__fa_2_217/A sky130_fd_sc_hd__and3_4_13/C
+ sky130_fd_sc_hd__xnor2_1_84/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_425 sky130_fd_sc_hd__xor2_1_425/B sky130_fd_sc_hd__buf_6_3/A
+ sky130_fd_sc_hd__xor2_1_426/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_95 vssd1 vccd1 sky130_fd_sc_hd__o21ai_2_9/Y sky130_fd_sc_hd__xnor2_1_95/Y
+ sky130_fd_sc_hd__xnor2_1_95/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_436 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__xor3_1_29/A
+ sky130_fd_sc_hd__xor2_1_436/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_447 sky130_fd_sc_hd__xor2_1_447/B sky130_fd_sc_hd__inv_2_58/A
+ sky130_fd_sc_hd__xor2_1_447/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_458 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__xor2_1_458/X
+ sky130_fd_sc_hd__xor2_1_458/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_469 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__xor2_1_469/X
+ sky130_fd_sc_hd__xor2_1_469/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1690 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_2_14 sky130_fd_sc_hd__clkinv_4_9/A sky130_fd_sc_hd__clkinv_2_14/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_25 sky130_fd_sc_hd__inv_2_134/A sky130_fd_sc_hd__dfxtp_1_5/Q
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_36 sky130_fd_sc_hd__clkinv_2_36/Y sky130_fd_sc_hd__clkinv_2_36/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_47 sky130_fd_sc_hd__clkinv_2_47/Y sky130_fd_sc_hd__clkinv_8_66/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_58 sky130_fd_sc_hd__clkinv_8_45/A wb_clk_i vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__or2_1_7 sky130_fd_sc_hd__or2_1_7/A sky130_fd_sc_hd__or2_1_7/X sky130_fd_sc_hd__or2_1_7/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_1
Xsky130_fd_sc_hd__buf_12_270 sky130_fd_sc_hd__buf_6_87/X sky130_fd_sc_hd__buf_12_270/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_281 sky130_fd_sc_hd__buf_12_77/X sky130_fd_sc_hd__buf_12_664/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_140 sky130_fd_sc_hd__xor2_1_276/X sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xor2_1_63/X sky130_fd_sc_hd__o21ai_1_60/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_292 sky130_fd_sc_hd__buf_12_98/X sky130_fd_sc_hd__buf_12_292/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_151 sky130_fd_sc_hd__xnor2_1_91/Y sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xnor2_1_28/Y sky130_fd_sc_hd__o21ai_1_81/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_162 sky130_fd_sc_hd__xnor2_1_98/Y sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xnor2_1_35/Y sky130_fd_sc_hd__a22oi_1_162/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_173 sky130_fd_sc_hd__nand2_1_129/A sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xnor2_1_50/Y sky130_fd_sc_hd__a22oi_1_173/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_184 sky130_fd_sc_hd__xnor2_1_123/Y sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xnor2_1_60/Y sky130_fd_sc_hd__a22oi_1_184/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_195 sky130_fd_sc_hd__clkbuf_1_3/X sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__nor2b_1_6/Y sky130_fd_sc_hd__nor2_1_72/Y sky130_fd_sc_hd__a22oi_1_195/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_470 sky130_fd_sc_hd__nand2_1_423/A sky130_fd_sc_hd__nor2_1_137/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_481 sky130_fd_sc_hd__a21oi_1_93/B1 sky130_fd_sc_hd__nand2_1_445/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_492 sky130_fd_sc_hd__xor2_1_399/B sky130_fd_sc_hd__o21ai_1_607/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_406 vssd1 vccd1 sky130_fd_sc_hd__inv_2_33/Y sky130_fd_sc_hd__nand2b_1_14/Y
+ sky130_fd_sc_hd__o21ai_1_406/B1 sky130_fd_sc_hd__xor2_1_217/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_417 vssd1 vccd1 sky130_fd_sc_hd__buf_2_9/X sky130_fd_sc_hd__nand2b_1_13/Y
+ sky130_fd_sc_hd__o21ai_1_417/B1 sky130_fd_sc_hd__xor2_1_226/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_428 vssd1 vccd1 sky130_fd_sc_hd__inv_2_30/Y sky130_fd_sc_hd__nand2b_1_14/Y
+ sky130_fd_sc_hd__o21ai_1_428/B1 sky130_fd_sc_hd__xor2_1_235/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_439 vssd1 vccd1 sky130_fd_sc_hd__inv_2_38/Y sky130_fd_sc_hd__nand2b_1_8/Y
+ sky130_fd_sc_hd__o21ai_1_439/B1 sky130_fd_sc_hd__xor2_1_244/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2_4_15 sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__or2b_2_2/A
+ sky130_fd_sc_hd__nor2_4_15/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__xor2_1_200 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__xor2_1_200/X
+ sky130_fd_sc_hd__xor2_1_200/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_211 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__xor2_1_211/X
+ sky130_fd_sc_hd__xor2_1_211/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_222 sky130_fd_sc_hd__xor2_1_383/B sky130_fd_sc_hd__xor3_1_19/B
+ sky130_fd_sc_hd__xor2_1_222/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_233 sky130_fd_sc_hd__fa_2_239/A sky130_fd_sc_hd__fa_2_145/A
+ sky130_fd_sc_hd__xor2_1_233/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_244 sky130_fd_sc_hd__xor2_1_362/B sky130_fd_sc_hd__fa_2_155/A
+ sky130_fd_sc_hd__xor2_1_244/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_255 sky130_fd_sc_hd__xor2_1_255/B sky130_fd_sc_hd__xor2_1_255/X
+ sky130_fd_sc_hd__a21oi_2_8/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_266 sky130_fd_sc_hd__fa_2_239/A sky130_fd_sc_hd__fa_2_173/A
+ sky130_fd_sc_hd__xor2_1_266/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_277 sky130_fd_sc_hd__dfxtp_2_5/Q sky130_fd_sc_hd__fa_2_188/B
+ sky130_fd_sc_hd__xor2_1_277/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_288 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__xor2_1_288/X
+ sky130_fd_sc_hd__xor2_1_288/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_299 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__xor2_1_299/X
+ sky130_fd_sc_hd__xor2_1_299/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_204 vssd1 vccd1 sky130_fd_sc_hd__buf_8_51/A sky130_fd_sc_hd__ha_2_35/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_215 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_215/X sky130_fd_sc_hd__clkinv_1_959/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_226 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_2/A1 sky130_fd_sc_hd__clkbuf_1_226/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_237 vssd1 vccd1 sky130_fd_sc_hd__buf_8_105/A sky130_fd_sc_hd__clkbuf_1_299/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_308 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__nor2_1_73/B sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__o21ai_1_523/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_248 vssd1 vccd1 sky130_fd_sc_hd__buf_8_157/A sky130_fd_sc_hd__clkbuf_1_325/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_319 vccd1 vssd1 sky130_fd_sc_hd__and3_4_17/X sky130_fd_sc_hd__buf_4_7/X
+ sky130_fd_sc_hd__buf_4_0/X sky130_fd_sc_hd__nor2_2_20/Y sky130_fd_sc_hd__buf_2_23/X
+ sky130_fd_sc_hd__o21ai_1_536/B1 sky130_fd_sc_hd__nor2b_2_4/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_259 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_260/A sky130_fd_sc_hd__clkbuf_1_305/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_2_6 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__clkinv_4_6/Y
+ sky130_fd_sc_hd__dfxtp_2_6/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_2
Xsky130_fd_sc_hd__decap_8_0 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__buf_2_60 vccd1 vssd1 sky130_fd_sc_hd__buf_8_2/A sky130_fd_sc_hd__buf_2_60/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_71 vccd1 vssd1 sky130_fd_sc_hd__buf_2_71/X sky130_fd_sc_hd__buf_2_71/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_82 vccd1 vssd1 sky130_fd_sc_hd__buf_2_82/X sky130_fd_sc_hd__buf_2_82/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_93 vccd1 vssd1 sky130_fd_sc_hd__buf_2_93/X sky130_fd_sc_hd__buf_2_93/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_4_9 vccd1 vssd1 sky130_fd_sc_hd__buf_4_9/X sky130_fd_sc_hd__buf_4_9/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__diode_2_0 sky130_fd_sc_hd__clkinv_2_37/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__and2_0_202 vccd1 vssd1 sky130_fd_sc_hd__and2_0_202/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_81/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_213 vccd1 vssd1 sky130_fd_sc_hd__and2_0_213/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_72/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_224 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_55/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_63/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_235 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_57/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_54/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_246 vccd1 vssd1 sky130_fd_sc_hd__and2_0_246/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_246/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_257 vccd1 vssd1 sky130_fd_sc_hd__and2_0_257/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__and2_0_257/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_268 vccd1 vssd1 sky130_fd_sc_hd__and2_0_268/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__xor2_1_644/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_279 vccd1 vssd1 sky130_fd_sc_hd__and2_0_279/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__fa_2_418/SUM vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__xor3_1_11 sky130_fd_sc_hd__xor3_1_11/X sky130_fd_sc_hd__xor3_1_11/C
+ sky130_fd_sc_hd__xor3_1_12/X sky130_fd_sc_hd__xor3_1_11/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__xor3_1_22 sky130_fd_sc_hd__xor3_1_22/X sky130_fd_sc_hd__xor3_1_22/C
+ sky130_fd_sc_hd__xor3_1_23/X sky130_fd_sc_hd__xor3_1_22/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__sdlclkp_2_7 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_8_3/Y
+ sky130_fd_sc_hd__dfxtp_1_154/CLK sky130_fd_sc_hd__o21ai_1_1/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__inv_4_9 sky130_fd_sc_hd__inv_4_9/Y sky130_fd_sc_hd__inv_4_9/A vccd1
+ vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__a22o_2_1 sky130_fd_sc_hd__nand2_1_7/B sky130_fd_sc_hd__fa_2_417/A
+ sky130_fd_sc_hd__or2_0_58/A sky130_fd_sc_hd__fa_2_417/B sky130_fd_sc_hd__nand2_1_8/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_2
Xsky130_fd_sc_hd__o31ai_1_0 sky130_fd_sc_hd__o31ai_1_0/Y sky130_fd_sc_hd__o31ai_1_0/A2
+ sky130_fd_sc_hd__o31ai_1_0/A1 sky130_fd_sc_hd__nand3_1_5/Y sky130_fd_sc_hd__o31ai_1_0/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__o31ai_1
Xsky130_fd_sc_hd__clkbuf_4_10 sky130_fd_sc_hd__clkbuf_4_10/X sky130_fd_sc_hd__a22o_1_67/A2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_203 vssd1 vccd1 sky130_fd_sc_hd__inv_2_18/Y sky130_fd_sc_hd__nand2b_1_5/Y
+ sky130_fd_sc_hd__a222oi_1_77/Y sky130_fd_sc_hd__xor2_1_30/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_21 sky130_fd_sc_hd__buf_8_83/A sky130_fd_sc_hd__inv_12_0/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_214 vssd1 vccd1 sky130_fd_sc_hd__inv_2_22/Y sky130_fd_sc_hd__nand2b_1_1/Y
+ sky130_fd_sc_hd__a222oi_1_85/Y sky130_fd_sc_hd__xor2_1_39/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_32 sky130_fd_sc_hd__buf_12_83/A sky130_fd_sc_hd__buf_8_19/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_225 vssd1 vccd1 sky130_fd_sc_hd__inv_2_20/Y sky130_fd_sc_hd__nand2b_1_7/Y
+ sky130_fd_sc_hd__a222oi_1_93/Y sky130_fd_sc_hd__xor2_1_50/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_43 la_data_out[56] sky130_fd_sc_hd__dfxtp_1_489/Q vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_236 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_295/A2 sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__o21ai_1_236/B1 sky130_fd_sc_hd__xor2_1_61/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_247 vssd1 vccd1 sky130_fd_sc_hd__inv_2_12/Y sky130_fd_sc_hd__nand2b_1_1/Y
+ sky130_fd_sc_hd__o21ai_1_247/B1 sky130_fd_sc_hd__xor2_1_70/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_258 vssd1 vccd1 sky130_fd_sc_hd__buf_2_1/X sky130_fd_sc_hd__nand2b_1_6/Y
+ sky130_fd_sc_hd__o21ai_1_258/B1 sky130_fd_sc_hd__xor2_1_81/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_269 vssd1 vccd1 sky130_fd_sc_hd__inv_2_16/Y sky130_fd_sc_hd__nand2b_1_6/Y
+ sky130_fd_sc_hd__o21ai_1_269/B1 sky130_fd_sc_hd__xor2_1_91/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nand2_1_607 sky130_fd_sc_hd__xnor2_1_169/A sky130_fd_sc_hd__nand2_1_608/Y
+ sky130_fd_sc_hd__nand2_1_607/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2_4_0 sky130_fd_sc_hd__nor2_4_0/Y sky130_fd_sc_hd__nor2_4_0/A
+ sky130_fd_sc_hd__nor2_4_0/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__nand2_1_618 sky130_fd_sc_hd__nand2_1_618/Y sky130_fd_sc_hd__nor2_1_203/A
+ sky130_fd_sc_hd__nor2_1_203/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__buf_8_160 sky130_fd_sc_hd__buf_8_160/A sky130_fd_sc_hd__buf_6_88/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nand2_1_629 sky130_fd_sc_hd__xnor2_1_177/A sky130_fd_sc_hd__nand2_1_630/Y
+ sky130_fd_sc_hd__nand2_1_629/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_403 sky130_fd_sc_hd__dfxtp_1_403/Q sky130_fd_sc_hd__clkinv_4_8/Y
+ sky130_fd_sc_hd__nor2b_1_112/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_414 sky130_fd_sc_hd__dfxtp_1_414/Q sky130_fd_sc_hd__dfxtp_1_417/CLK
+ sky130_fd_sc_hd__nor2b_1_101/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_425 sky130_fd_sc_hd__dfxtp_1_425/Q sky130_fd_sc_hd__dfxtp_1_427/CLK
+ sky130_fd_sc_hd__nor2b_1_90/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_436 sky130_fd_sc_hd__dfxtp_1_436/Q sky130_fd_sc_hd__dfxtp_1_439/CLK
+ sky130_fd_sc_hd__nor2b_1_111/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_447 sky130_fd_sc_hd__dfxtp_1_447/Q sky130_fd_sc_hd__dfxtp_1_451/CLK
+ sky130_fd_sc_hd__nor2b_1_100/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_458 sky130_fd_sc_hd__dfxtp_1_458/Q sky130_fd_sc_hd__dfxtp_1_459/CLK
+ sky130_fd_sc_hd__nor2b_1_88/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_469 sky130_fd_sc_hd__ha_2_51/A sky130_fd_sc_hd__dfxtp_1_515/CLK
+ sky130_fd_sc_hd__and2_0_353/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a222oi_1_105 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__or2_0_60/A
+ sky130_fd_sc_hd__or2_0_61/A sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__or2_0_42/B
+ sky130_fd_sc_hd__o21ai_1_237/B1 sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2b_1_17 sky130_fd_sc_hd__nand2b_1_17/Y sky130_fd_sc_hd__nor2_1_167/B
+ sky130_fd_sc_hd__nor2_1_167/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a222oi_1_116 vccd1 vssd1 sky130_fd_sc_hd__and3_4_2/X sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__nor2_1_73/B sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__o21ai_1_253/B1 sky130_fd_sc_hd__and2b_4_4/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2b_1_28 sky130_fd_sc_hd__nand2b_1_28/Y sky130_fd_sc_hd__or2_0_84/A
+ sky130_fd_sc_hd__or2_0_78/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a222oi_1_127 vccd1 vssd1 sky130_fd_sc_hd__and3_4_8/X sky130_fd_sc_hd__buf_2_4/X
+ sky130_fd_sc_hd__buf_6_5/X sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__o21ai_1_267/B1 sky130_fd_sc_hd__nor2b_2_2/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_138 vccd1 vssd1 sky130_fd_sc_hd__and3_4_6/X sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__inv_6_0/Y sky130_fd_sc_hd__nor2_1_72/Y sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__o21ai_1_282/B1 sky130_fd_sc_hd__nor2b_1_6/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__o21ai_1_770 vssd1 vccd1 sky130_fd_sc_hd__inv_2_47/Y sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__o21ai_1_770/B1 sky130_fd_sc_hd__xor2_1_545/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_149 vccd1 vssd1 sky130_fd_sc_hd__and3_4_7/X sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__buf_4_6/X sky130_fd_sc_hd__nor2_2_7/Y sky130_fd_sc_hd__buf_4_1/X
+ sky130_fd_sc_hd__o21ai_1_294/B1 sky130_fd_sc_hd__nor2b_2_1/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__o21ai_1_781 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_126/A sky130_fd_sc_hd__nor2_1_187/Y
+ sky130_fd_sc_hd__nand2_1_582/Y sky130_fd_sc_hd__xnor2_1_159/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_308 sky130_fd_sc_hd__fa_2_299/A sky130_fd_sc_hd__fa_2_308/SUM
+ sky130_fd_sc_hd__fa_2_308/A sky130_fd_sc_hd__fa_2_308/B sky130_fd_sc_hd__fa_2_308/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o21ai_1_792 vssd1 vccd1 sky130_fd_sc_hd__buf_2_12/X sky130_fd_sc_hd__nand2b_2_6/Y
+ sky130_fd_sc_hd__o21ai_1_792/B1 sky130_fd_sc_hd__xor2_1_566/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_319 sky130_fd_sc_hd__fa_2_312/CIN sky130_fd_sc_hd__fa_2_321/B
+ sky130_fd_sc_hd__fa_2_319/A sky130_fd_sc_hd__fa_2_319/B sky130_fd_sc_hd__xor2_1_484/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_8_13 sky130_fd_sc_hd__clkinv_8_15/A sky130_fd_sc_hd__clkinv_8_13/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_24 sky130_fd_sc_hd__clkinv_8_24/Y sky130_fd_sc_hd__clkinv_8_24/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_35 sky130_fd_sc_hd__clkinv_8_41/A sky130_fd_sc_hd__clkinv_8_35/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_46 sky130_fd_sc_hd__clkinv_8_47/A sky130_fd_sc_hd__clkinv_8_46/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_57 sky130_fd_sc_hd__dfxtp_1_2/CLK sky130_fd_sc_hd__clkinv_8_6/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_11 sky130_fd_sc_hd__buf_12_11/A sky130_fd_sc_hd__buf_12_11/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_8_68 sky130_fd_sc_hd__clkinv_8_68/Y sky130_fd_sc_hd__clkinv_8_68/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_22 sky130_fd_sc_hd__inv_2_141/Y sky130_fd_sc_hd__buf_12_22/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_8_79 sky130_fd_sc_hd__clkinv_8_80/A sky130_fd_sc_hd__clkinv_8_79/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_33 sky130_fd_sc_hd__buf_12_33/A sky130_fd_sc_hd__buf_12_33/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_44 sky130_fd_sc_hd__buf_12_44/A sky130_fd_sc_hd__buf_12_44/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_55 sky130_fd_sc_hd__buf_12_55/A sky130_fd_sc_hd__buf_12_55/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_66 sky130_fd_sc_hd__buf_12_66/A sky130_fd_sc_hd__buf_12_66/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_77 sky130_fd_sc_hd__buf_12_77/A sky130_fd_sc_hd__buf_12_77/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_88 sky130_fd_sc_hd__buf_12_88/A sky130_fd_sc_hd__buf_12_88/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_99 sky130_fd_sc_hd__buf_8_144/X sky130_fd_sc_hd__buf_12_99/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_2_6 vccd1 vssd1 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__buf_2_6/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__inv_2_6 sky130_fd_sc_hd__inv_2_6/A sky130_fd_sc_hd__inv_2_6/Y vccd1
+ vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__nor2_1_16 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_16/Y
+ sky130_fd_sc_hd__nor2_1_16/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_27 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_27/Y
+ sky130_fd_sc_hd__nor2_1_27/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_38 sky130_fd_sc_hd__nor2_1_42/B sky130_fd_sc_hd__nor2_1_38/Y
+ sky130_fd_sc_hd__nor2_1_38/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_49 sky130_fd_sc_hd__nor2_1_49/B sky130_fd_sc_hd__nor2_1_49/Y
+ sky130_fd_sc_hd__nor2_1_49/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_12_509 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__and2_0_60 vccd1 vssd1 sky130_fd_sc_hd__and2_0_60/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__or2_0_60/B vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_71 vccd1 vssd1 sky130_fd_sc_hd__and2_0_71/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__buf_4_3/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_404 sky130_fd_sc_hd__nand2_1_404/Y sky130_fd_sc_hd__or2_0_35/A
+ sky130_fd_sc_hd__or2_0_35/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_82 vccd1 vssd1 sky130_fd_sc_hd__and2_0_82/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__buf_4_5/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_415 sky130_fd_sc_hd__nand2_1_415/Y sky130_fd_sc_hd__or2_0_37/A
+ sky130_fd_sc_hd__or2_0_37/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_93 vccd1 vssd1 sky130_fd_sc_hd__and2_0_93/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__or2_0_58/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_426 sky130_fd_sc_hd__nand2_1_426/Y sky130_fd_sc_hd__nor2_1_139/A
+ sky130_fd_sc_hd__nor2_1_139/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_437 sky130_fd_sc_hd__nand2_1_437/Y sky130_fd_sc_hd__nor2_1_145/A
+ sky130_fd_sc_hd__nor2_1_145/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_448 sky130_fd_sc_hd__xnor2_1_112/A sky130_fd_sc_hd__nand2_1_449/Y
+ sky130_fd_sc_hd__nand2_1_448/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_459 sky130_fd_sc_hd__nand2_1_459/Y sky130_fd_sc_hd__buf_2_23/X
+ sky130_fd_sc_hd__buf_2_31/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_17 sky130_fd_sc_hd__and3_4_25/C sky130_fd_sc_hd__nor2b_1_17/Y
+ sky130_fd_sc_hd__and3_4_25/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_28 sky130_fd_sc_hd__fa_2_416/A sky130_fd_sc_hd__fa_2_463/B
+ sky130_fd_sc_hd__mux2_2_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_39 sky130_fd_sc_hd__mux2_2_15/X sky130_fd_sc_hd__nor2b_1_39/Y
+ sky130_fd_sc_hd__buf_2_214/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1006 sky130_fd_sc_hd__clkinv_1_1007/A sky130_fd_sc_hd__clkinv_2_1/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1017 sky130_fd_sc_hd__clkinv_1_1017/Y sky130_fd_sc_hd__clkinv_1_1017/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1028 sky130_fd_sc_hd__buf_8_138/A sky130_fd_sc_hd__clkinv_1_1028/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_70 sky130_fd_sc_hd__buf_8_70/A sky130_fd_sc_hd__buf_8_70/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__clkinv_1_1039 sky130_fd_sc_hd__inv_4_14/A sky130_fd_sc_hd__inv_2_93/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_81 sky130_fd_sc_hd__buf_8_81/A sky130_fd_sc_hd__buf_8_81/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_200 sky130_fd_sc_hd__xor2_1_596/A sky130_fd_sc_hd__dfxtp_2_2/CLK
+ sky130_fd_sc_hd__and2_0_51/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_8_92 sky130_fd_sc_hd__buf_8_92/A sky130_fd_sc_hd__buf_8_92/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__decap_12_1508 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_211 sky130_fd_sc_hd__xor2_1_504/A sky130_fd_sc_hd__dfxtp_2_0/CLK
+ sky130_fd_sc_hd__and2_0_68/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1519 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_222 sky130_fd_sc_hd__xnor2_1_118/A sky130_fd_sc_hd__dfxtp_1_234/CLK
+ sky130_fd_sc_hd__and2_0_16/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_233 sky130_fd_sc_hd__xnor2_1_97/A sky130_fd_sc_hd__dfxtp_1_234/CLK
+ sky130_fd_sc_hd__and2_0_73/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_244 sky130_fd_sc_hd__fa_2_170/A sky130_fd_sc_hd__clkinv_4_4/Y
+ sky130_fd_sc_hd__and2_0_89/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_255 sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__dfxtp_1_266/CLK
+ sky130_fd_sc_hd__and2_0_39/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_266 sky130_fd_sc_hd__xor2_1_104/A sky130_fd_sc_hd__dfxtp_1_266/CLK
+ sky130_fd_sc_hd__and2_0_69/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_277 sky130_fd_sc_hd__dfxtp_1_277/Q sky130_fd_sc_hd__dfxtp_1_2/CLK
+ sky130_fd_sc_hd__and2_0_253/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_288 sky130_fd_sc_hd__a22oi_1_6/B2 sky130_fd_sc_hd__dfxtp_1_2/CLK
+ sky130_fd_sc_hd__and2_0_264/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_299 sky130_fd_sc_hd__dfxtp_1_299/Q sky130_fd_sc_hd__clkinv_8_6/Y
+ sky130_fd_sc_hd__and2_0_275/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o22ai_1_8 sky130_fd_sc_hd__o22ai_1_8/A2 sky130_fd_sc_hd__o22ai_1_8/B1
+ sky130_fd_sc_hd__o22ai_1_8/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__o22ai_1_9/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_105 sky130_fd_sc_hd__fa_2_101/A sky130_fd_sc_hd__fa_2_106/B
+ sky130_fd_sc_hd__fa_2_105/A sky130_fd_sc_hd__fa_2_105/B sky130_fd_sc_hd__xor2_1_140/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_116 sky130_fd_sc_hd__fa_2_114/CIN sky130_fd_sc_hd__fa_2_119/A
+ sky130_fd_sc_hd__fa_2_116/A sky130_fd_sc_hd__fa_2_116/B sky130_fd_sc_hd__xor2_1_162/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_127 sky130_fd_sc_hd__fa_2_125/B sky130_fd_sc_hd__fa_2_128/A
+ sky130_fd_sc_hd__fa_2_127/A sky130_fd_sc_hd__fa_2_127/B sky130_fd_sc_hd__fa_2_127/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_138 sky130_fd_sc_hd__nor2_1_98/A sky130_fd_sc_hd__or2_0_16/B
+ sky130_fd_sc_hd__fa_2_138/A sky130_fd_sc_hd__fa_2_138/B sky130_fd_sc_hd__fa_2_138/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_149 sky130_fd_sc_hd__xor3_1_17/B sky130_fd_sc_hd__fa_2_150/CIN
+ sky130_fd_sc_hd__fa_2_149/A sky130_fd_sc_hd__fa_2_149/B sky130_fd_sc_hd__xor2_1_224/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_100 vccd1 vssd1 sky130_fd_sc_hd__buf_2_100/X sky130_fd_sc_hd__buf_2_100/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_111 vccd1 vssd1 sky130_fd_sc_hd__buf_2_111/X sky130_fd_sc_hd__buf_2_111/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_122 vccd1 vssd1 sky130_fd_sc_hd__buf_2_122/X sky130_fd_sc_hd__buf_2_122/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_15 sky130_fd_sc_hd__o22ai_1_48/B1 sky130_fd_sc_hd__o22ai_1_15/B1
+ sky130_fd_sc_hd__o22ai_1_15/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__inv_4_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_133 vccd1 vssd1 sky130_fd_sc_hd__buf_2_133/X sky130_fd_sc_hd__inv_2_2/Y
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_26 sky130_fd_sc_hd__o22ai_1_36/B1 sky130_fd_sc_hd__o21ai_1_6/A2
+ sky130_fd_sc_hd__o22ai_1_26/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__inv_4_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_144 vccd1 vssd1 sky130_fd_sc_hd__buf_2_144/X sky130_fd_sc_hd__buf_2_144/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_37 sky130_fd_sc_hd__nor2_1_29/A sky130_fd_sc_hd__o22ai_1_37/B1
+ sky130_fd_sc_hd__o22ai_1_37/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_155 vccd1 vssd1 sky130_fd_sc_hd__mux2_8_0/A1 sky130_fd_sc_hd__buf_2_155/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_48 sky130_fd_sc_hd__nor2_1_19/A sky130_fd_sc_hd__o22ai_1_48/B1
+ sky130_fd_sc_hd__o22ai_1_48/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_166 vccd1 vssd1 sky130_fd_sc_hd__buf_2_166/X sky130_fd_sc_hd__buf_2_53/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_59 sky130_fd_sc_hd__nor2_1_8/A sky130_fd_sc_hd__o22ai_1_4/A2
+ sky130_fd_sc_hd__o22ai_1_59/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_177 vccd1 vssd1 la_data_out[60] sky130_fd_sc_hd__ha_2_23/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_188 vccd1 vssd1 sky130_fd_sc_hd__buf_2_188/X sky130_fd_sc_hd__buf_2_44/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_199 vccd1 vssd1 la_data_out[92] sky130_fd_sc_hd__nand2_2_4/Y
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__ha_2_0 vssd1 vccd1 sky130_fd_sc_hd__ha_2_0/A sky130_fd_sc_hd__xor3_1_5/C
+ sky130_fd_sc_hd__fa_2_6/A sky130_fd_sc_hd__ha_2_0/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__buf_4_17 vccd1 vssd1 sky130_fd_sc_hd__buf_4_17/X sky130_fd_sc_hd__buf_4_17/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_28 vccd1 vssd1 sky130_fd_sc_hd__buf_4_28/X sky130_fd_sc_hd__buf_8_72/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_39 vccd1 vssd1 sky130_fd_sc_hd__buf_4_39/X sky130_fd_sc_hd__buf_4_39/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__clkbuf_1_11 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_11/X sky130_fd_sc_hd__a32oi_1_0/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_480 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__buf_4_2/X sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__o21ai_1_767/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_22 vssd1 vccd1 sky130_fd_sc_hd__or2_0_61/B sky130_fd_sc_hd__or2_0_42/B
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_491 vccd1 vssd1 sky130_fd_sc_hd__and3_4_26/X sky130_fd_sc_hd__or2_0_72/A
+ sky130_fd_sc_hd__or2_0_71/B sky130_fd_sc_hd__nor2_2_31/Y sky130_fd_sc_hd__buf_2_29/X
+ sky130_fd_sc_hd__o21ai_1_782/B1 sky130_fd_sc_hd__nor2b_1_12/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_33 vssd1 vccd1 sky130_fd_sc_hd__buf_8_120/A sky130_fd_sc_hd__ha_2_35/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_44 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_44/X sky130_fd_sc_hd__inv_2_106/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_55 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_55/X sky130_fd_sc_hd__clkbuf_1_56/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_66 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_67/A sky130_fd_sc_hd__clkbuf_4_19/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_77 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_21/A1 sky130_fd_sc_hd__clkbuf_1_77/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_88 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_34/A1 sky130_fd_sc_hd__clkbuf_1_88/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_99 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_5/A1 sky130_fd_sc_hd__clkbuf_1_99/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__or2_0_13 sky130_fd_sc_hd__or2_0_66/A sky130_fd_sc_hd__or2_0_13/X
+ sky130_fd_sc_hd__or2_0_60/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_24 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__or2_0_24/X
+ sky130_fd_sc_hd__or2_0_24/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_35 sky130_fd_sc_hd__or2_0_35/A sky130_fd_sc_hd__or2_0_35/X
+ sky130_fd_sc_hd__or2_0_35/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_46 sky130_fd_sc_hd__or2_0_66/A sky130_fd_sc_hd__or2_0_46/X
+ sky130_fd_sc_hd__buf_4_5/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_57 sky130_fd_sc_hd__or2_0_58/A sky130_fd_sc_hd__or2_0_57/X
+ sky130_fd_sc_hd__or2_0_9/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_68 sky130_fd_sc_hd__or2_0_68/A sky130_fd_sc_hd__or2_0_68/X
+ sky130_fd_sc_hd__or2_0_68/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_79 sky130_fd_sc_hd__or2_0_79/A sky130_fd_sc_hd__or2_0_79/X
+ sky130_fd_sc_hd__or2_0_79/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__buf_12_0 sky130_fd_sc_hd__buf_2_25/A sky130_fd_sc_hd__or2_0_53/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_600 sky130_fd_sc_hd__buf_12_600/A sky130_fd_sc_hd__buf_12_600/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_611 sky130_fd_sc_hd__buf_12_611/A sky130_fd_sc_hd__buf_12_611/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_622 sky130_fd_sc_hd__buf_12_622/A sky130_fd_sc_hd__buf_12_622/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_633 sky130_fd_sc_hd__buf_12_633/A sky130_fd_sc_hd__buf_12_633/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_4_104 sky130_fd_sc_hd__clkinv_8_61/Y sky130_fd_sc_hd__clkinv_8_18/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_12_644 sky130_fd_sc_hd__buf_12_644/A sky130_fd_sc_hd__buf_12_644/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_4_115 sky130_fd_sc_hd__clkinv_4_115/A sky130_fd_sc_hd__clkinv_8_19/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_12_655 sky130_fd_sc_hd__buf_12_655/A sky130_fd_sc_hd__buf_12_655/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_666 sky130_fd_sc_hd__buf_12_666/A sky130_fd_sc_hd__buf_12_666/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_677 sky130_fd_sc_hd__buf_12_677/A sky130_fd_sc_hd__buf_12_677/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_306 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_317 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_201 sky130_fd_sc_hd__xnor2_1_19/A sky130_fd_sc_hd__nand2_1_202/Y
+ sky130_fd_sc_hd__or2_0_3/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_328 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_800 sky130_fd_sc_hd__and2_0_307/A sky130_fd_sc_hd__clkinv_1_800/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_212 sky130_fd_sc_hd__xnor2_1_23/A sky130_fd_sc_hd__nand2_1_213/Y
+ sky130_fd_sc_hd__or2_0_6/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_339 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_811 sky130_fd_sc_hd__nand2_1_800/A sky130_fd_sc_hd__nor2_1_256/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_223 sky130_fd_sc_hd__nand2_1_223/Y sky130_fd_sc_hd__or2_0_7/A
+ sky130_fd_sc_hd__or2_0_7/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_822 sky130_fd_sc_hd__clkinv_1_822/Y sky130_fd_sc_hd__nand2_1_823/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_234 sky130_fd_sc_hd__xnor2_1_33/A sky130_fd_sc_hd__nand2_1_235/Y
+ sky130_fd_sc_hd__nand2_1_234/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_833 sky130_fd_sc_hd__inv_2_70/A sky130_fd_sc_hd__ha_2_33/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_245 sky130_fd_sc_hd__nand2_1_245/Y sky130_fd_sc_hd__nor2_1_76/Y
+ sky130_fd_sc_hd__nand2_1_256/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_844 sky130_fd_sc_hd__inv_2_93/A la_data_out[39] vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_256 sky130_fd_sc_hd__nand2_1_256/Y sky130_fd_sc_hd__nand2_1_263/A
+ sky130_fd_sc_hd__nand2_1_256/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_855 sky130_fd_sc_hd__clkinv_1_855/Y sky130_fd_sc_hd__clkinv_8_9/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_267 sky130_fd_sc_hd__nand2_1_267/Y sky130_fd_sc_hd__nand2_1_273/A
+ sky130_fd_sc_hd__nor2_1_89/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_866 sky130_fd_sc_hd__clkinv_1_866/Y sky130_fd_sc_hd__clkinv_4_81/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_278 sky130_fd_sc_hd__nand2_1_278/Y sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__buf_2_4/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_877 sky130_fd_sc_hd__clkinv_1_877/Y sky130_fd_sc_hd__buf_4_42/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_289 sky130_fd_sc_hd__xor2_1_191/A sky130_fd_sc_hd__nand2_1_290/Y
+ sky130_fd_sc_hd__nand2_1_289/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_888 sky130_fd_sc_hd__clkinv_1_888/Y sky130_fd_sc_hd__inv_4_19/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_899 sky130_fd_sc_hd__clkinv_1_899/Y sky130_fd_sc_hd__clkinv_4_89/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__conb_1_11 sky130_fd_sc_hd__conb_1_11/LO sky130_fd_sc_hd__conb_1_11/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_22 sky130_fd_sc_hd__conb_1_22/LO sky130_fd_sc_hd__conb_1_22/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_33 sky130_fd_sc_hd__conb_1_33/LO sky130_fd_sc_hd__conb_1_33/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1305 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_44 sky130_fd_sc_hd__conb_1_44/LO sky130_fd_sc_hd__conb_1_44/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1316 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_55 sky130_fd_sc_hd__conb_1_55/LO sky130_fd_sc_hd__conb_1_55/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1327 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_66 sky130_fd_sc_hd__conb_1_66/LO sky130_fd_sc_hd__conb_1_66/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1338 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_77 sky130_fd_sc_hd__conb_1_77/LO sky130_fd_sc_hd__conb_1_77/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1349 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_88 sky130_fd_sc_hd__conb_1_88/LO sky130_fd_sc_hd__conb_1_88/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_99 sky130_fd_sc_hd__conb_1_99/LO sky130_fd_sc_hd__conb_1_99/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__mux2_2_6 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_6/A1 sky130_fd_sc_hd__buf_2_81/X
+ sky130_fd_sc_hd__mux2_8_0/S sky130_fd_sc_hd__or2_0_76/B vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__decap_12_840 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_851 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_862 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_873 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_884 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_895 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_607 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__fa_2_404/B
+ sky130_fd_sc_hd__xor2_1_607/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_790 sky130_fd_sc_hd__xnor2_1_290/A sky130_fd_sc_hd__nand2_1_791/Y
+ sky130_fd_sc_hd__or2_0_99/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_618 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__fa_2_409/B
+ sky130_fd_sc_hd__xor2_1_618/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_629 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__or2_0_67/B
+ sky130_fd_sc_hd__xor2_1_629/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1850 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1861 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1872 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o2bb2ai_1_2 sky130_fd_sc_hd__maj3_1_3/C sky130_fd_sc_hd__a21oi_1_197/Y
+ sky130_fd_sc_hd__xnor2_1_309/A sky130_fd_sc_hd__ha_2_56/B la_data_out[49] vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__fa_2_480 sky130_fd_sc_hd__nor2_1_259/B sky130_fd_sc_hd__or2_0_105/A
+ sky130_fd_sc_hd__fa_2_480/A sky130_fd_sc_hd__fa_2_480/B sky130_fd_sc_hd__nor2b_1_59/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_491 sky130_fd_sc_hd__or2_0_110/B sky130_fd_sc_hd__nor2_1_265/A
+ sky130_fd_sc_hd__fa_2_491/A sky130_fd_sc_hd__fa_2_491/B sky130_fd_sc_hd__nor2b_1_81/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_1_107 io_oeb[32] sky130_fd_sc_hd__conb_1_35/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_118 io_oeb[21] sky130_fd_sc_hd__conb_1_24/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_129 io_oeb[10] sky130_fd_sc_hd__conb_1_13/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor3b_1_1 wbs_we_i sky130_fd_sc_hd__nor3b_1_1/Y wbs_ack_o sky130_fd_sc_hd__nor4_1_1/D
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor3b_1
Xsky130_fd_sc_hd__o21ai_1_7 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_7/A2 sky130_fd_sc_hd__nor2_4_4/B
+ sky130_fd_sc_hd__o21ai_1_7/B1 sky130_fd_sc_hd__fa_2_45/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2_1_201 sky130_fd_sc_hd__nor2_1_207/Y sky130_fd_sc_hd__nor2_1_201/Y
+ sky130_fd_sc_hd__nor2_1_204/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_212 sky130_fd_sc_hd__buf_2_27/X sky130_fd_sc_hd__nor2_1_212/Y
+ sky130_fd_sc_hd__buf_2_24/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_223 sky130_fd_sc_hd__mux2_2_42/X sky130_fd_sc_hd__nor2_1_223/Y
+ sky130_fd_sc_hd__mux2_2_22/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_234 sky130_fd_sc_hd__xor2_1_659/X sky130_fd_sc_hd__nor2_1_234/Y
+ sky130_fd_sc_hd__nor2_1_234/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_245 sky130_fd_sc_hd__nor2_1_246/Y sky130_fd_sc_hd__nor2_1_245/Y
+ sky130_fd_sc_hd__nor2_1_247/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_256 sky130_fd_sc_hd__nor2_1_256/B sky130_fd_sc_hd__nor2_1_256/Y
+ sky130_fd_sc_hd__nor2_1_256/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_267 sky130_fd_sc_hd__nor2_1_267/B sky130_fd_sc_hd__nor2_1_267/Y
+ sky130_fd_sc_hd__nor2_1_278/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_278 sky130_fd_sc_hd__nor2_1_278/B sky130_fd_sc_hd__nor2_1_278/Y
+ sky130_fd_sc_hd__a21o_2_0/B1 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_430 sky130_fd_sc_hd__buf_12_430/A sky130_fd_sc_hd__buf_12_635/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_441 sky130_fd_sc_hd__buf_12_441/A sky130_fd_sc_hd__buf_12_441/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_452 sky130_fd_sc_hd__buf_12_452/A sky130_fd_sc_hd__buf_12_452/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_463 sky130_fd_sc_hd__buf_12_463/A sky130_fd_sc_hd__buf_12_510/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_474 sky130_fd_sc_hd__buf_12_474/A sky130_fd_sc_hd__buf_12_516/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_103 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_485 sky130_fd_sc_hd__buf_12_485/A sky130_fd_sc_hd__buf_12_573/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_114 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_496 sky130_fd_sc_hd__buf_12_496/A sky130_fd_sc_hd__buf_12_496/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_125 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_136 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_147 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_158 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_630 sky130_fd_sc_hd__nand2_1_672/A sky130_fd_sc_hd__nor2_1_223/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_169 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_641 sky130_fd_sc_hd__clkinv_1_641/Y sky130_fd_sc_hd__nand2_1_695/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_204 vssd1 vccd1 sky130_fd_sc_hd__or2_0_78/A sky130_fd_sc_hd__nor2b_1_25/A
+ sky130_fd_sc_hd__mux2_2_47/X vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_652 sky130_fd_sc_hd__o22ai_1_86/B1 la_data_out[79] vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_215 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_215/B sky130_fd_sc_hd__or2_0_89/B
+ sky130_fd_sc_hd__xnor2_1_215/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_663 sky130_fd_sc_hd__clkinv_1_663/Y sky130_fd_sc_hd__nand2_1_731/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_226 vssd1 vccd1 la_data_out[85] sky130_fd_sc_hd__xnor2_1_226/Y
+ la_data_out[67] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_674 sky130_fd_sc_hd__nand2_1_747/A sky130_fd_sc_hd__nor2_1_240/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_237 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_4/B sky130_fd_sc_hd__xnor2_1_237/Y
+ la_data_out[67] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_685 sky130_fd_sc_hd__nand2_1_760/A sky130_fd_sc_hd__nor2_1_247/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_248 vssd1 vccd1 la_data_out[77] sky130_fd_sc_hd__xnor2_1_248/Y
+ la_data_out[71] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_696 sky130_fd_sc_hd__clkinv_1_696/Y sky130_fd_sc_hd__nand2_1_783/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_259 vssd1 vccd1 la_data_out[77] sky130_fd_sc_hd__xnor2_1_259/Y
+ sky130_fd_sc_hd__or2_0_79/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_1102 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1113 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1124 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1135 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1146 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1157 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand3_1_3 sky130_fd_sc_hd__nor2_4_7/B sky130_fd_sc_hd__nand3_1_3/A
+ sky130_fd_sc_hd__nand3_1_3/C sky130_fd_sc_hd__nor2_1_42/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__decap_12_1168 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1179 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__fah_1_8 sky130_fd_sc_hd__nor2_1_196/A sky130_fd_sc_hd__fah_1_8/B
+ sky130_fd_sc_hd__fah_1_8/A sky130_fd_sc_hd__nor2_2_30/B sky130_fd_sc_hd__fah_1_8/CI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__fah_1
Xsky130_fd_sc_hd__a222oi_1_50 vccd1 vssd1 sky130_fd_sc_hd__and3_4_4/X sky130_fd_sc_hd__buf_4_1/X
+ sky130_fd_sc_hd__nor2_2_5/A sky130_fd_sc_hd__nor2_1_61/Y sky130_fd_sc_hd__nor2_2_5/B
+ sky130_fd_sc_hd__a222oi_1_50/Y sky130_fd_sc_hd__nor2b_1_4/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__sdlclkp_2_15 sky130_fd_sc_hd__conb_1_148/LO sky130_fd_sc_hd__clkinv_2_47/Y
+ sky130_fd_sc_hd__dfxtp_1_480/CLK sky130_fd_sc_hd__o21ai_1_909/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__a222oi_1_61 vccd1 vssd1 sky130_fd_sc_hd__and3_4_5/X sky130_fd_sc_hd__nor2_2_5/B
+ sky130_fd_sc_hd__nor2_2_4/B sky130_fd_sc_hd__nor2_1_68/Y sky130_fd_sc_hd__buf_2_4/X
+ sky130_fd_sc_hd__a222oi_1_61/Y sky130_fd_sc_hd__nor2b_1_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_72 vccd1 vssd1 sky130_fd_sc_hd__and3_4_2/X sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__or2_0_66/A sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__or2_0_60/B
+ sky130_fd_sc_hd__a222oi_1_72/Y sky130_fd_sc_hd__and2b_4_4/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_83 vccd1 vssd1 sky130_fd_sc_hd__and3_4_5/X sky130_fd_sc_hd__buf_4_1/X
+ sky130_fd_sc_hd__nor2_2_5/A sky130_fd_sc_hd__nor2_1_68/Y sky130_fd_sc_hd__nor2_2_5/B
+ sky130_fd_sc_hd__a222oi_1_83/Y sky130_fd_sc_hd__nor2b_1_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_670 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_30 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_30/B sky130_fd_sc_hd__inv_2_23/A
+ sky130_fd_sc_hd__xnor2_1_30/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__a222oi_1_94 vccd1 vssd1 sky130_fd_sc_hd__and3_4_8/X sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__nor2_2_10/B sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__buf_6_4/X
+ sky130_fd_sc_hd__a222oi_1_94/Y sky130_fd_sc_hd__nor2b_2_2/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__xnor2_1_41 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_41/B sky130_fd_sc_hd__xnor2_1_41/Y
+ sky130_fd_sc_hd__xnor2_1_41/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_681 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_692 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_52 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_52/B sky130_fd_sc_hd__inv_2_18/A
+ sky130_fd_sc_hd__xnor2_1_52/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_63 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_63/B sky130_fd_sc_hd__buf_2_8/A
+ sky130_fd_sc_hd__xnor2_1_63/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_404 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__xor2_1_404/X
+ sky130_fd_sc_hd__xor2_1_404/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_74 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_74/B sky130_fd_sc_hd__xnor2_1_74/Y
+ sky130_fd_sc_hd__xnor2_1_74/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_415 sky130_fd_sc_hd__fa_2_281/A sky130_fd_sc_hd__fa_2_280/B
+ sky130_fd_sc_hd__xor2_1_415/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_85 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_85/B sky130_fd_sc_hd__xnor2_1_85/Y
+ sky130_fd_sc_hd__xnor2_1_85/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_426 sky130_fd_sc_hd__xor2_1_426/B sky130_fd_sc_hd__xor2_1_426/X
+ sky130_fd_sc_hd__xor3_1_20/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_96 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_96/B sky130_fd_sc_hd__inv_2_40/A
+ sky130_fd_sc_hd__xnor2_1_96/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_437 sky130_fd_sc_hd__xor2_1_548/B sky130_fd_sc_hd__xor2_1_437/X
+ sky130_fd_sc_hd__xor2_1_437/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_448 sky130_fd_sc_hd__fa_2_379/A sky130_fd_sc_hd__xor2_1_448/X
+ sky130_fd_sc_hd__xor2_1_448/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_459 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__fa_2_302/B
+ sky130_fd_sc_hd__xor2_1_459/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1680 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1691 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_0 sky130_fd_sc_hd__buf_12_459/A sky130_fd_sc_hd__clkbuf_16_0/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__nor4_1_0 sky130_fd_sc_hd__ha_2_4/A sky130_fd_sc_hd__ha_2_3/A sky130_fd_sc_hd__nor4_1_0/Y
+ sky130_fd_sc_hd__ha_2_6/A sky130_fd_sc_hd__ha_2_5/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor4_1
Xsky130_fd_sc_hd__decap_12_4 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_2_15 sky130_fd_sc_hd__inv_2_79/A sky130_fd_sc_hd__clkinv_2_15/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_26 sky130_fd_sc_hd__inv_2_136/A sky130_fd_sc_hd__buf_8_92/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_37 sky130_fd_sc_hd__clkinv_2_37/Y sky130_fd_sc_hd__buf_4_26/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_48 sky130_fd_sc_hd__clkinv_2_48/Y sky130_fd_sc_hd__clkinv_8_19/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_59 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkinv_8_56/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__or2_1_8 sky130_fd_sc_hd__or2_1_8/A sky130_fd_sc_hd__or2_1_8/X sky130_fd_sc_hd__or2_1_8/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_1
Xsky130_fd_sc_hd__buf_12_260 sky130_fd_sc_hd__buf_6_59/X sky130_fd_sc_hd__buf_12_483/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_271 sky130_fd_sc_hd__buf_6_86/X sky130_fd_sc_hd__buf_12_326/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_130 sky130_fd_sc_hd__xnor2_2_1/Y sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__o2bb2ai_1_0/Y sky130_fd_sc_hd__o21ai_1_40/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_282 sky130_fd_sc_hd__buf_12_87/X sky130_fd_sc_hd__buf_12_282/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_141 sky130_fd_sc_hd__xor2_1_276/X sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xor2_1_63/X sky130_fd_sc_hd__o21ai_1_61/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_293 sky130_fd_sc_hd__buf_12_293/A sky130_fd_sc_hd__buf_12_293/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_152 sky130_fd_sc_hd__xor2_1_330/X sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xor2_1_117/X sky130_fd_sc_hd__o21ai_1_84/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_163 sky130_fd_sc_hd__xnor2_1_98/Y sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xnor2_1_35/Y sky130_fd_sc_hd__a22oi_1_163/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_174 sky130_fd_sc_hd__nand2_1_131/A sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xor2_1_187/X sky130_fd_sc_hd__a22oi_1_174/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_185 sky130_fd_sc_hd__xnor2_1_123/Y sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xnor2_1_60/Y sky130_fd_sc_hd__a22oi_1_185/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_196 sky130_fd_sc_hd__clkbuf_1_3/X sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__nor2b_2_1/Y sky130_fd_sc_hd__nor2_2_7/Y sky130_fd_sc_hd__a22oi_1_196/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_460 sky130_fd_sc_hd__o21ai_1_535/B1 sky130_fd_sc_hd__nand2_1_400/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_471 sky130_fd_sc_hd__nand2_1_425/A sky130_fd_sc_hd__nor2_1_139/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_482 sky130_fd_sc_hd__nand2_1_439/A sky130_fd_sc_hd__nor2_1_146/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_493 sky130_fd_sc_hd__nand2_1_456/A sky130_fd_sc_hd__nor2_1_154/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_407 vssd1 vccd1 sky130_fd_sc_hd__inv_2_31/Y sky130_fd_sc_hd__nand2b_1_13/Y
+ sky130_fd_sc_hd__o21ai_1_407/B1 sky130_fd_sc_hd__xor2_1_218/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_418 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_454/A2 sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_418/B1 sky130_fd_sc_hd__xor2_1_227/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_429 vssd1 vccd1 sky130_fd_sc_hd__buf_2_7/X sky130_fd_sc_hd__nand2b_1_11/Y
+ sky130_fd_sc_hd__o21ai_1_429/B1 sky130_fd_sc_hd__xor2_1_236/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2_4_16 sky130_fd_sc_hd__nor2_4_16/Y sky130_fd_sc_hd__nor2_4_16/A
+ sky130_fd_sc_hd__nor2_4_16/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__xor2_1_201 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__or2_0_23/A
+ sky130_fd_sc_hd__xor2_1_201/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_212 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__nor2_4_8/B
+ sky130_fd_sc_hd__xor2_1_212/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_223 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__xor3_1_19/A
+ sky130_fd_sc_hd__xor2_1_223/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_234 sky130_fd_sc_hd__xor2_1_234/B sky130_fd_sc_hd__xor2_1_234/X
+ sky130_fd_sc_hd__a21oi_2_7/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_245 sky130_fd_sc_hd__dfxtp_2_5/Q sky130_fd_sc_hd__xor2_1_245/X
+ sky130_fd_sc_hd__xor2_1_245/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_256 sky130_fd_sc_hd__dfxtp_2_5/Q sky130_fd_sc_hd__xor2_1_256/X
+ sky130_fd_sc_hd__xor2_1_256/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_267 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__xor2_1_267/X
+ sky130_fd_sc_hd__xor2_1_267/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_278 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__fa_2_188/A
+ sky130_fd_sc_hd__xor2_1_278/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_289 sky130_fd_sc_hd__fa_2_217/A sky130_fd_sc_hd__fa_2_200/B
+ sky130_fd_sc_hd__xor2_1_289/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_205 vssd1 vccd1 sky130_fd_sc_hd__buf_8_43/A sky130_fd_sc_hd__clkbuf_1_56/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_216 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2_15/A la_data_out[48]
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_227 vssd1 vccd1 sky130_fd_sc_hd__buf_12_15/A sky130_fd_sc_hd__inv_2_150/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_238 vssd1 vccd1 sky130_fd_sc_hd__buf_2_165/A sky130_fd_sc_hd__inv_4_14/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_309 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__and2_0_87/A
+ sky130_fd_sc_hd__buf_6_0/X sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__o21ai_1_524/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_249 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_249/X sky130_fd_sc_hd__clkinv_1_959/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_2_7 sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__dfxtp_2_7/CLK
+ la_data_out[56] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_2
Xsky130_fd_sc_hd__decap_8_1 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__buf_2_50 vccd1 vssd1 sky130_fd_sc_hd__buf_2_50/X sky130_fd_sc_hd__buf_2_50/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_61 vccd1 vssd1 sky130_fd_sc_hd__buf_2_61/X sky130_fd_sc_hd__buf_2_61/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_72 vccd1 vssd1 sky130_fd_sc_hd__buf_2_72/X sky130_fd_sc_hd__buf_2_72/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_83 vccd1 vssd1 sky130_fd_sc_hd__buf_2_83/X sky130_fd_sc_hd__buf_2_83/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_94 vccd1 vssd1 sky130_fd_sc_hd__buf_2_94/X sky130_fd_sc_hd__buf_2_94/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__diode_2_1 sky130_fd_sc_hd__clkbuf_4_20/X vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__and2_0_203 vccd1 vssd1 sky130_fd_sc_hd__and2_0_203/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_80/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_214 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_85/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_71/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_225 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_87/D sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__o21ai_1_62/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_236 vccd1 vssd1 sky130_fd_sc_hd__and2_0_236/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_236/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_247 vccd1 vssd1 sky130_fd_sc_hd__and2_0_247/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__o21ai_1_44/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_258 vccd1 vssd1 sky130_fd_sc_hd__and2_0_258/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__xor2_1_649/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_269 vccd1 vssd1 sky130_fd_sc_hd__and2_0_269/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__and2_0_269/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__xor3_1_12 sky130_fd_sc_hd__xor3_1_12/X sky130_fd_sc_hd__xor3_1_12/C
+ sky130_fd_sc_hd__xor3_1_13/X sky130_fd_sc_hd__xor3_1_12/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__xor3_1_23 sky130_fd_sc_hd__xor3_1_23/X sky130_fd_sc_hd__xor3_1_23/C
+ sky130_fd_sc_hd__xor3_1_24/X sky130_fd_sc_hd__xor3_1_23/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__sdlclkp_2_8 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_8_3/Y
+ sky130_fd_sc_hd__dfxtp_1_152/CLK sky130_fd_sc_hd__o21ai_1_1/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__a22o_2_2 sky130_fd_sc_hd__nand2_1_7/B sky130_fd_sc_hd__mux2_2_9/X
+ sky130_fd_sc_hd__or2_0_58/B sky130_fd_sc_hd__fa_2_418/A sky130_fd_sc_hd__nand2_1_8/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_2
Xsky130_fd_sc_hd__o31ai_1_1 sky130_fd_sc_hd__o31ai_1_1/Y sky130_fd_sc_hd__nand3_1_5/B
+ sky130_fd_sc_hd__o31ai_1_1/A1 sky130_fd_sc_hd__a21o_2_0/X sky130_fd_sc_hd__o31ai_1_1/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__o31ai_1
Xsky130_fd_sc_hd__clkinv_1_290 sky130_fd_sc_hd__and2_0_185/A sky130_fd_sc_hd__a222oi_1_34/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkbuf_4_11 sky130_fd_sc_hd__clkbuf_4_11/X sky130_fd_sc_hd__and2_0_352/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_204 vssd1 vccd1 sky130_fd_sc_hd__inv_2_13/Y sky130_fd_sc_hd__nand2b_1_7/Y
+ sky130_fd_sc_hd__a222oi_1_78/Y sky130_fd_sc_hd__xor2_1_31/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_22 sky130_fd_sc_hd__clkbuf_4_22/X sky130_fd_sc_hd__buf_6_10/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_215 vssd1 vccd1 sky130_fd_sc_hd__inv_2_12/Y sky130_fd_sc_hd__nand2b_1_7/Y
+ sky130_fd_sc_hd__a222oi_1_86/Y sky130_fd_sc_hd__xor2_1_40/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_33 sky130_fd_sc_hd__buf_12_88/A sky130_fd_sc_hd__buf_8_152/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_226 vssd1 vccd1 sky130_fd_sc_hd__inv_2_21/Y sky130_fd_sc_hd__nand2b_1_1/Y
+ sky130_fd_sc_hd__a222oi_1_94/Y sky130_fd_sc_hd__xor2_1_51/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_44 sky130_fd_sc_hd__buf_2_16/A sky130_fd_sc_hd__buf_6_91/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_237 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_237/A2 sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__o21ai_1_237/B1 sky130_fd_sc_hd__xor2_1_62/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_248 vssd1 vccd1 sky130_fd_sc_hd__inv_2_17/Y sky130_fd_sc_hd__nand2b_1_7/Y
+ sky130_fd_sc_hd__o21ai_1_248/B1 sky130_fd_sc_hd__xor2_1_71/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_259 vssd1 vccd1 sky130_fd_sc_hd__inv_2_19/Y sky130_fd_sc_hd__nand2b_1_7/Y
+ sky130_fd_sc_hd__o21ai_1_259/B1 sky130_fd_sc_hd__xor2_1_82/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nand2_1_608 sky130_fd_sc_hd__nand2_1_608/Y sky130_fd_sc_hd__nor2_2_30/A
+ sky130_fd_sc_hd__nor2_2_30/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2_4_1 sky130_fd_sc_hd__nor2_4_1/Y sky130_fd_sc_hd__inv_4_7/A
+ sky130_fd_sc_hd__nor2_4_1/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__buf_8_150 sky130_fd_sc_hd__buf_8_150/A sky130_fd_sc_hd__buf_8_150/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nand2_1_619 sky130_fd_sc_hd__xnor2_1_174/A sky130_fd_sc_hd__nand2_1_620/Y
+ sky130_fd_sc_hd__nand2_1_619/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__buf_8_161 sky130_fd_sc_hd__buf_8_161/A sky130_fd_sc_hd__buf_4_34/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_404 sky130_fd_sc_hd__dfxtp_1_404/Q sky130_fd_sc_hd__clkinv_4_8/Y
+ sky130_fd_sc_hd__nor2b_1_111/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_415 sky130_fd_sc_hd__dfxtp_1_415/Q sky130_fd_sc_hd__dfxtp_1_423/CLK
+ sky130_fd_sc_hd__nor2b_1_100/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_426 sky130_fd_sc_hd__dfxtp_1_426/Q sky130_fd_sc_hd__dfxtp_1_427/CLK
+ sky130_fd_sc_hd__nor2b_1_88/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_437 sky130_fd_sc_hd__dfxtp_1_437/Q sky130_fd_sc_hd__dfxtp_1_439/CLK
+ sky130_fd_sc_hd__nor2b_1_110/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_448 sky130_fd_sc_hd__dfxtp_1_448/Q sky130_fd_sc_hd__dfxtp_1_451/CLK
+ sky130_fd_sc_hd__nor2b_1_99/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_459 sky130_fd_sc_hd__dfxtp_1_459/Q sky130_fd_sc_hd__dfxtp_1_459/CLK
+ sky130_fd_sc_hd__nor2b_1_89/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a222oi_1_106 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__buf_4_5/X sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__o21ai_1_240/B1 sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2b_1_18 sky130_fd_sc_hd__nand2b_1_18/Y sky130_fd_sc_hd__and3_1_2/C
+ sky130_fd_sc_hd__and3_1_2/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a222oi_1_117 vccd1 vssd1 sky130_fd_sc_hd__and3_4_5/X sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__inv_6_0/Y sky130_fd_sc_hd__nor2_1_68/Y sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__o21ai_1_254/B1 sky130_fd_sc_hd__nor2b_1_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2b_1_29 sky130_fd_sc_hd__nand2b_1_29/Y sky130_fd_sc_hd__or2_0_84/A
+ sky130_fd_sc_hd__or2_0_77/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a222oi_1_128 vccd1 vssd1 sky130_fd_sc_hd__and3_4_5/X sky130_fd_sc_hd__clkbuf_1_3/X
+ sky130_fd_sc_hd__or2_0_53/A sky130_fd_sc_hd__nor2_1_68/Y sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__o21ai_1_268/B1 sky130_fd_sc_hd__nor2b_1_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__o21ai_1_760 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_780/A2 sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_760/B1 sky130_fd_sc_hd__xor2_1_535/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_139 vccd1 vssd1 sky130_fd_sc_hd__and3_4_1/X sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__buf_6_1/X sky130_fd_sc_hd__nor2_2_9/Y sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__o21ai_1_284/B1 sky130_fd_sc_hd__and2b_4_3/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__o21ai_1_771 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_771/A2 sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_771/B1 sky130_fd_sc_hd__xor2_1_546/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_782 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_2/Y sky130_fd_sc_hd__nand2b_1_15/Y
+ sky130_fd_sc_hd__o21ai_1_782/B1 sky130_fd_sc_hd__xor2_1_555/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_309 sky130_fd_sc_hd__fa_2_308/CIN sky130_fd_sc_hd__fa_2_316/B
+ sky130_fd_sc_hd__fa_2_309/A sky130_fd_sc_hd__fa_2_309/B sky130_fd_sc_hd__xor2_1_469/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o21ai_1_793 vssd1 vccd1 sky130_fd_sc_hd__inv_2_46/Y sky130_fd_sc_hd__nand2b_1_16/Y
+ sky130_fd_sc_hd__o21ai_1_793/B1 sky130_fd_sc_hd__xor2_1_567/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkinv_8_14 sky130_fd_sc_hd__clkinv_8_14/Y sky130_fd_sc_hd__clkinv_8_15/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_25 sky130_fd_sc_hd__clkinv_8_28/A sky130_fd_sc_hd__clkinv_8_25/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_36 sky130_fd_sc_hd__clkinv_8_39/A sky130_fd_sc_hd__clkinv_8_41/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_47 sky130_fd_sc_hd__clkinv_8_47/Y sky130_fd_sc_hd__clkinv_8_47/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_58 sky130_fd_sc_hd__clkinv_8_62/A sky130_fd_sc_hd__clkinv_8_58/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_12 sky130_fd_sc_hd__buf_12_12/A sky130_fd_sc_hd__buf_12_12/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_8_69 sky130_fd_sc_hd__clkinv_8_70/A sky130_fd_sc_hd__clkinv_8_69/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_23 sky130_fd_sc_hd__inv_2_144/Y sky130_fd_sc_hd__buf_12_23/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_34 sky130_fd_sc_hd__buf_12_34/A sky130_fd_sc_hd__buf_12_34/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_45 sky130_fd_sc_hd__buf_12_45/A sky130_fd_sc_hd__buf_12_45/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_56 sky130_fd_sc_hd__buf_12_56/A sky130_fd_sc_hd__buf_12_56/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_67 sky130_fd_sc_hd__buf_8_16/X sky130_fd_sc_hd__buf_12_67/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_78 sky130_fd_sc_hd__buf_12_78/A sky130_fd_sc_hd__buf_12_78/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_89 sky130_fd_sc_hd__buf_8_139/X sky130_fd_sc_hd__buf_12_89/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_2_7 vccd1 vssd1 sky130_fd_sc_hd__buf_2_7/X sky130_fd_sc_hd__buf_2_7/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o21ai_2_10 sky130_fd_sc_hd__a21oi_1_85/Y sky130_fd_sc_hd__xnor2_1_98/B
+ sky130_fd_sc_hd__a21oi_1_91/Y sky130_fd_sc_hd__o21ai_2_10/A1 vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__o21ai_2
Xsky130_fd_sc_hd__inv_2_7 sky130_fd_sc_hd__inv_2_7/A sky130_fd_sc_hd__inv_2_7/Y vccd1
+ vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__nor2_1_17 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_17/Y
+ sky130_fd_sc_hd__nor2_1_17/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_28 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_28/Y
+ sky130_fd_sc_hd__nor2_1_28/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_39 sky130_fd_sc_hd__nor3_1_0/C sky130_fd_sc_hd__nor2_1_39/Y
+ sky130_fd_sc_hd__nor2_1_39/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__and2_0_50 vccd1 vssd1 sky130_fd_sc_hd__and2_0_50/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__nor2_1_73/B vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_61 vccd1 vssd1 sky130_fd_sc_hd__and2_0_61/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__or2_0_60/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_72 vccd1 vssd1 sky130_fd_sc_hd__and2_0_72/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__buf_4_2/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_405 sky130_fd_sc_hd__xnor2_1_96/A sky130_fd_sc_hd__nand2_1_406/Y
+ sky130_fd_sc_hd__nand2_1_405/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_83 vccd1 vssd1 sky130_fd_sc_hd__and2_0_83/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__buf_4_4/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_416 sky130_fd_sc_hd__nand2_1_416/Y sky130_fd_sc_hd__nor2_1_134/Y
+ sky130_fd_sc_hd__nand2_1_427/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_94 vccd1 vssd1 sky130_fd_sc_hd__and2_0_94/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__or2_0_58/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_427 sky130_fd_sc_hd__nand2_1_427/Y sky130_fd_sc_hd__nand2_1_434/A
+ sky130_fd_sc_hd__nand2_1_427/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_438 sky130_fd_sc_hd__nand2_1_438/Y sky130_fd_sc_hd__nand2_1_444/A
+ sky130_fd_sc_hd__nor2_1_105/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_449 sky130_fd_sc_hd__nand2_1_449/Y sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__buf_2_19/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_18 sky130_fd_sc_hd__or2_0_84/A sky130_fd_sc_hd__or2_0_85/B
+ sky130_fd_sc_hd__inv_2_65/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_29 sky130_fd_sc_hd__fa_2_416/B sky130_fd_sc_hd__nor2b_1_29/Y
+ sky130_fd_sc_hd__buf_2_214/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1007 sky130_fd_sc_hd__clkinv_1_1007/Y sky130_fd_sc_hd__clkinv_1_1007/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1018 sky130_fd_sc_hd__clkinv_1_1019/A sky130_fd_sc_hd__buf_4_40/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_60 sky130_fd_sc_hd__buf_8_60/A sky130_fd_sc_hd__buf_8_60/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__clkinv_1_1029 sky130_fd_sc_hd__buf_8_8/A sky130_fd_sc_hd__inv_4_10/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_71 sky130_fd_sc_hd__buf_8_71/A sky130_fd_sc_hd__buf_8_71/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_82 sky130_fd_sc_hd__buf_8_82/A sky130_fd_sc_hd__buf_8_82/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_201 sky130_fd_sc_hd__xnor2_1_164/A sky130_fd_sc_hd__dfxtp_2_2/CLK
+ sky130_fd_sc_hd__and2_0_79/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_8_93 sky130_fd_sc_hd__buf_8_93/A sky130_fd_sc_hd__buf_8_93/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__decap_12_1509 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_212 sky130_fd_sc_hd__fa_2_338/A sky130_fd_sc_hd__dfxtp_2_0/CLK
+ sky130_fd_sc_hd__and2_0_98/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_223 sky130_fd_sc_hd__xor2_1_409/A sky130_fd_sc_hd__dfxtp_1_234/CLK
+ sky130_fd_sc_hd__and2_0_30/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_234 sky130_fd_sc_hd__xor2_1_344/A sky130_fd_sc_hd__dfxtp_1_234/CLK
+ sky130_fd_sc_hd__and2_0_74/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_245 sky130_fd_sc_hd__xnor2_1_71/A sky130_fd_sc_hd__clkinv_4_4/Y
+ sky130_fd_sc_hd__and2_0_101/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_256 sky130_fd_sc_hd__xnor2_1_46/A sky130_fd_sc_hd__dfxtp_1_269/CLK
+ sky130_fd_sc_hd__and2_0_37/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_267 sky130_fd_sc_hd__fa_2_75/A sky130_fd_sc_hd__dfxtp_1_269/CLK
+ sky130_fd_sc_hd__and2_0_70/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_278 sky130_fd_sc_hd__dfxtp_1_278/Q sky130_fd_sc_hd__dfxtp_1_2/CLK
+ sky130_fd_sc_hd__and2_0_254/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_289 sky130_fd_sc_hd__a22oi_1_4/B2 sky130_fd_sc_hd__clkinv_8_6/Y
+ sky130_fd_sc_hd__and2_0_265/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o22ai_1_9 sky130_fd_sc_hd__o22ai_1_9/A2 sky130_fd_sc_hd__o22ai_1_9/B1
+ sky130_fd_sc_hd__o22ai_1_9/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__o22ai_1_9/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_106 sky130_fd_sc_hd__fa_2_103/B sky130_fd_sc_hd__fa_2_108/CIN
+ sky130_fd_sc_hd__fa_2_106/A sky130_fd_sc_hd__fa_2_106/B sky130_fd_sc_hd__fa_2_106/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o21ai_1_590 vssd1 vccd1 sky130_fd_sc_hd__inv_2_30/Y sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_590/B1 sky130_fd_sc_hd__xor2_1_385/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_117 sky130_fd_sc_hd__fa_2_115/B sky130_fd_sc_hd__fa_2_119/CIN
+ sky130_fd_sc_hd__fa_2_117/A sky130_fd_sc_hd__fa_2_117/B sky130_fd_sc_hd__xor2_1_160/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_128 sky130_fd_sc_hd__fa_2_126/B sky130_fd_sc_hd__fa_2_129/CIN
+ sky130_fd_sc_hd__fa_2_128/A sky130_fd_sc_hd__fa_2_128/B sky130_fd_sc_hd__xor2_1_177/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_139 sky130_fd_sc_hd__fa_2_138/CIN sky130_fd_sc_hd__or2_0_23/B
+ sky130_fd_sc_hd__fa_2_139/A sky130_fd_sc_hd__fa_2_139/B sky130_fd_sc_hd__xor2_1_200/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_101 vccd1 vssd1 sky130_fd_sc_hd__buf_2_101/X sky130_fd_sc_hd__buf_2_101/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_112 vccd1 vssd1 sky130_fd_sc_hd__buf_2_112/X sky130_fd_sc_hd__buf_2_112/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_123 vccd1 vssd1 sky130_fd_sc_hd__buf_2_123/X sky130_fd_sc_hd__buf_2_123/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_16 sky130_fd_sc_hd__o22ai_1_47/B1 sky130_fd_sc_hd__o22ai_1_16/B1
+ sky130_fd_sc_hd__o22ai_1_16/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__inv_4_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_134 vccd1 vssd1 sky130_fd_sc_hd__buf_2_134/X sky130_fd_sc_hd__inv_2_1/Y
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_27 sky130_fd_sc_hd__o22ai_1_34/B1 sky130_fd_sc_hd__o21ai_1_4/A2
+ sky130_fd_sc_hd__o22ai_1_27/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__inv_4_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_145 vccd1 vssd1 sky130_fd_sc_hd__buf_2_145/X sky130_fd_sc_hd__buf_2_145/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_38 sky130_fd_sc_hd__nor2_1_28/A sky130_fd_sc_hd__o22ai_1_38/B1
+ sky130_fd_sc_hd__o22ai_1_38/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_156 vccd1 vssd1 sky130_fd_sc_hd__buf_8_97/A sky130_fd_sc_hd__buf_2_156/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_49 sky130_fd_sc_hd__nor2_1_18/A sky130_fd_sc_hd__o22ai_1_49/B1
+ sky130_fd_sc_hd__o22ai_1_49/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_167 vccd1 vssd1 sky130_fd_sc_hd__buf_2_167/X sky130_fd_sc_hd__buf_2_167/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_178 vccd1 vssd1 la_data_out[59] sky130_fd_sc_hd__ha_2_24/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_189 vccd1 vssd1 sky130_fd_sc_hd__nand2_1_8/B sky130_fd_sc_hd__buf_2_189/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__ha_2_1 vssd1 vccd1 sky130_fd_sc_hd__ha_2_1/A sky130_fd_sc_hd__xor3_1_15/C
+ sky130_fd_sc_hd__ha_2_1/SUM sky130_fd_sc_hd__ha_2_1/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__buf_4_18 vccd1 vssd1 sky130_fd_sc_hd__buf_4_18/X sky130_fd_sc_hd__buf_4_18/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_29 vccd1 vssd1 sky130_fd_sc_hd__buf_4_29/X sky130_fd_sc_hd__buf_4_29/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__a222oi_1_470 vccd1 vssd1 sky130_fd_sc_hd__and3_4_21/X sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__nor2_2_10/B sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__buf_6_4/X
+ sky130_fd_sc_hd__o21ai_1_757/B1 sky130_fd_sc_hd__and2b_4_12/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_12 vssd1 vccd1 sky130_fd_sc_hd__o21ai_2_0/B1 sky130_fd_sc_hd__and2_0_9/B
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_481 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__nor2_2_10/B
+ sky130_fd_sc_hd__buf_6_4/X sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__o21ai_1_769/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_23 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_23/X sky130_fd_sc_hd__nor2_4_5/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_492 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__nor2_2_10/B sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__buf_6_4/X
+ sky130_fd_sc_hd__o21ai_1_784/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_34 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_34/X sky130_fd_sc_hd__ha_2_36/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_45 vssd1 vccd1 sky130_fd_sc_hd__inv_2_108/A wbs_dat_i[1]
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_56 vssd1 vccd1 sky130_fd_sc_hd__buf_2_60/A sky130_fd_sc_hd__clkbuf_1_56/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_67 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4_16/A sky130_fd_sc_hd__clkbuf_1_67/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_78 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_22/A1 sky130_fd_sc_hd__clkbuf_1_78/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_89 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_0/A1 sky130_fd_sc_hd__clkbuf_1_89/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__and2_4_0 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__and2_4_0/B
+ la_data_out[32] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__and2_4
Xsky130_fd_sc_hd__or2_0_14 sky130_fd_sc_hd__or2_0_60/A sky130_fd_sc_hd__or2_0_14/X
+ sky130_fd_sc_hd__or2_0_60/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_25 sky130_fd_sc_hd__or2_0_53/A sky130_fd_sc_hd__or2_0_25/X
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_36 sky130_fd_sc_hd__or2_0_9/A sky130_fd_sc_hd__or2_0_36/X
+ sky130_fd_sc_hd__or2_0_9/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_47 sky130_fd_sc_hd__buf_4_5/X sky130_fd_sc_hd__or2_0_47/X
+ sky130_fd_sc_hd__buf_4_4/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_58 sky130_fd_sc_hd__or2_0_58/A sky130_fd_sc_hd__or2_0_58/X
+ sky130_fd_sc_hd__or2_0_58/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_69 sky130_fd_sc_hd__or2_0_69/A sky130_fd_sc_hd__or2_0_69/X
+ sky130_fd_sc_hd__or2_0_69/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__buf_12_1 sky130_fd_sc_hd__buf_2_68/A sky130_fd_sc_hd__buf_12_1/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_601 sky130_fd_sc_hd__buf_12_601/A sky130_fd_sc_hd__buf_12_601/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_612 sky130_fd_sc_hd__buf_12_612/A sky130_fd_sc_hd__buf_12_612/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_623 sky130_fd_sc_hd__buf_12_623/A sky130_fd_sc_hd__buf_12_623/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_634 sky130_fd_sc_hd__buf_12_634/A sky130_fd_sc_hd__buf_12_634/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_4_105 sky130_fd_sc_hd__clkinv_8_18/A sky130_fd_sc_hd__dfxtp_1_8/CLK
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_12_645 sky130_fd_sc_hd__buf_12_645/A sky130_fd_sc_hd__buf_12_645/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_4_116 sky130_fd_sc_hd__clkinv_8_73/Y sky130_fd_sc_hd__clkinv_4_117/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_12_656 sky130_fd_sc_hd__buf_12_656/A sky130_fd_sc_hd__buf_12_656/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_667 sky130_fd_sc_hd__buf_12_667/A sky130_fd_sc_hd__buf_12_667/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_678 sky130_fd_sc_hd__buf_12_678/A sky130_fd_sc_hd__buf_12_679/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_307 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_318 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_202 sky130_fd_sc_hd__nand2_1_202/Y sky130_fd_sc_hd__or2_0_3/A
+ sky130_fd_sc_hd__or2_0_3/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_329 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_801 sky130_fd_sc_hd__and2_0_306/A sky130_fd_sc_hd__clkinv_1_801/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_213 sky130_fd_sc_hd__nand2_1_213/Y sky130_fd_sc_hd__or2_0_6/A
+ sky130_fd_sc_hd__or2_0_6/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_812 sky130_fd_sc_hd__clkinv_1_812/Y sky130_fd_sc_hd__nand2_1_803/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_224 sky130_fd_sc_hd__nand2_1_224/Y sky130_fd_sc_hd__or2_0_18/X
+ sky130_fd_sc_hd__nor2_1_70/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_823 sky130_fd_sc_hd__nand2_1_824/A sky130_fd_sc_hd__nor2_1_262/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_235 sky130_fd_sc_hd__nand2_1_235/Y sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__nor2_1_73/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_834 sky130_fd_sc_hd__buf_8_100/A sky130_fd_sc_hd__inv_2_70/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_246 sky130_fd_sc_hd__xnor2_1_37/A sky130_fd_sc_hd__nand2_1_247/Y
+ sky130_fd_sc_hd__nand2_1_246/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_845 sky130_fd_sc_hd__clkinv_1_845/Y sky130_fd_sc_hd__clkinv_1_846/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_257 sky130_fd_sc_hd__xnor2_1_40/A sky130_fd_sc_hd__nand2_1_258/Y
+ sky130_fd_sc_hd__nand2_1_257/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_856 sky130_fd_sc_hd__clkinv_1_856/Y sky130_fd_sc_hd__clkinv_8_9/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_268 sky130_fd_sc_hd__xnor2_1_45/A sky130_fd_sc_hd__nand2_1_269/Y
+ sky130_fd_sc_hd__nand2_1_268/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_867 sky130_fd_sc_hd__clkinv_1_867/Y sky130_fd_sc_hd__inv_2_95/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_279 sky130_fd_sc_hd__xnor2_1_50/A sky130_fd_sc_hd__nand2_1_280/Y
+ sky130_fd_sc_hd__nand2_1_279/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_878 sky130_fd_sc_hd__clkinv_1_878/Y sky130_fd_sc_hd__buf_4_42/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_889 sky130_fd_sc_hd__clkinv_1_889/Y sky130_fd_sc_hd__inv_4_20/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__conb_1_12 sky130_fd_sc_hd__conb_1_12/LO sky130_fd_sc_hd__conb_1_12/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_23 sky130_fd_sc_hd__conb_1_23/LO sky130_fd_sc_hd__conb_1_23/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_34 sky130_fd_sc_hd__conb_1_34/LO sky130_fd_sc_hd__conb_1_34/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1306 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_45 sky130_fd_sc_hd__conb_1_45/LO sky130_fd_sc_hd__conb_1_45/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1317 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_56 sky130_fd_sc_hd__conb_1_56/LO sky130_fd_sc_hd__conb_1_56/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1328 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_67 sky130_fd_sc_hd__conb_1_67/LO sky130_fd_sc_hd__conb_1_67/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1339 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_78 sky130_fd_sc_hd__conb_1_78/LO sky130_fd_sc_hd__conb_1_78/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_89 sky130_fd_sc_hd__conb_1_89/LO sky130_fd_sc_hd__conb_1_89/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__mux2_2_7 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_7/A1 sky130_fd_sc_hd__buf_2_88/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__or2_0_73/A vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__decap_12_830 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_841 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_852 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_863 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_874 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_885 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_896 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_780 sky130_fd_sc_hd__nand2_1_780/Y sky130_fd_sc_hd__nor2_1_251/A
+ sky130_fd_sc_hd__nor2_1_251/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_608 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__fah_1_15/CI
+ sky130_fd_sc_hd__xor2_1_608/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_791 sky130_fd_sc_hd__nand2_1_791/Y sky130_fd_sc_hd__or2_0_99/A
+ sky130_fd_sc_hd__or2_0_99/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_619 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__fa_2_408/B
+ sky130_fd_sc_hd__xor2_1_619/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1840 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1851 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1862 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__fa_2_470 sky130_fd_sc_hd__nor2_1_254/B sky130_fd_sc_hd__or2_0_100/A
+ sky130_fd_sc_hd__fa_2_470/A sky130_fd_sc_hd__fa_2_470/B sky130_fd_sc_hd__nor2b_1_39/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_481 sky130_fd_sc_hd__or2_0_105/B sky130_fd_sc_hd__nor2_1_260/A
+ sky130_fd_sc_hd__fa_2_481/A sky130_fd_sc_hd__fa_2_481/B sky130_fd_sc_hd__nor2b_1_61/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_492 sky130_fd_sc_hd__nor2_1_265/B sky130_fd_sc_hd__or2_0_111/B
+ sky130_fd_sc_hd__fa_2_492/A sky130_fd_sc_hd__fa_2_492/B sky130_fd_sc_hd__nor2b_1_83/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_1_108 io_oeb[31] sky130_fd_sc_hd__conb_1_34/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_119 io_oeb[20] sky130_fd_sc_hd__conb_1_23/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_8 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_8/A2 sky130_fd_sc_hd__nor2_4_4/B
+ sky130_fd_sc_hd__o21ai_1_8/B1 sky130_fd_sc_hd__fa_2_56/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2_1_202 sky130_fd_sc_hd__buf_2_21/X sky130_fd_sc_hd__nor2_1_202/Y
+ sky130_fd_sc_hd__buf_2_20/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_213 sky130_fd_sc_hd__nor2_1_216/Y sky130_fd_sc_hd__nor2_1_213/Y
+ sky130_fd_sc_hd__nor2_1_214/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_224 sky130_fd_sc_hd__mux2_2_39/X sky130_fd_sc_hd__nor2_1_224/Y
+ sky130_fd_sc_hd__mux2_2_8/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_235 sky130_fd_sc_hd__xor2_1_660/X sky130_fd_sc_hd__nor2_1_235/Y
+ sky130_fd_sc_hd__nor2_1_235/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_246 sky130_fd_sc_hd__nor2_1_246/B sky130_fd_sc_hd__nor2_1_246/Y
+ sky130_fd_sc_hd__nor2_1_246/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_257 sky130_fd_sc_hd__nor2_1_257/B sky130_fd_sc_hd__nor2_1_257/Y
+ sky130_fd_sc_hd__nor2_1_257/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_268 sky130_fd_sc_hd__nor2_1_268/B sky130_fd_sc_hd__o31ai_1_0/A2
+ sky130_fd_sc_hd__nor2_1_275/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_279 sky130_fd_sc_hd__maj3_1_1/X sky130_fd_sc_hd__nor2_1_279/Y
+ sky130_fd_sc_hd__ha_2_49/SUM vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_420 sky130_fd_sc_hd__buf_12_420/A sky130_fd_sc_hd__buf_12_466/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_431 sky130_fd_sc_hd__buf_12_431/A sky130_fd_sc_hd__buf_12_473/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_442 sky130_fd_sc_hd__buf_12_442/A sky130_fd_sc_hd__buf_12_442/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_453 sky130_fd_sc_hd__buf_12_453/A sky130_fd_sc_hd__buf_12_453/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_464 sky130_fd_sc_hd__buf_12_464/A sky130_fd_sc_hd__buf_12_464/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_475 sky130_fd_sc_hd__buf_12_475/A sky130_fd_sc_hd__buf_12_521/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_104 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_486 sky130_fd_sc_hd__buf_12_486/A sky130_fd_sc_hd__buf_12_525/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_115 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_497 sky130_fd_sc_hd__buf_12_497/A sky130_fd_sc_hd__buf_12_606/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_126 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_137 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_148 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_620 sky130_fd_sc_hd__nand2_1_652/A sky130_fd_sc_hd__nor2_1_218/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_159 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_631 sky130_fd_sc_hd__clkinv_1_631/Y sky130_fd_sc_hd__nand2_1_675/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_642 sky130_fd_sc_hd__nand2_1_696/A sky130_fd_sc_hd__nor2_1_229/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_205 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_205/B sky130_fd_sc_hd__a22o_1_21/B1
+ sky130_fd_sc_hd__xnor2_1_205/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_653 sky130_fd_sc_hd__o22ai_1_101/B1 la_data_out[81] vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_216 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_216/B sky130_fd_sc_hd__or2_0_88/B
+ sky130_fd_sc_hd__xnor2_1_216/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_664 sky130_fd_sc_hd__xnor2_1_206/B sky130_fd_sc_hd__a21oi_1_153/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_227 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_4/B sky130_fd_sc_hd__xnor2_1_227/Y
+ sky130_fd_sc_hd__or2_1_10/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_675 sky130_fd_sc_hd__clkinv_1_675/Y sky130_fd_sc_hd__nand2_1_750/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_238 vssd1 vccd1 la_data_out[77] sky130_fd_sc_hd__xnor2_1_238/Y
+ sky130_fd_sc_hd__or2_0_82/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_686 sky130_fd_sc_hd__xor2_1_662/A sky130_fd_sc_hd__o21ai_1_887/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_249 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_4/B sky130_fd_sc_hd__xnor2_1_249/Y
+ la_data_out[68] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_697 sky130_fd_sc_hd__clkinv_1_697/Y sky130_fd_sc_hd__nand2_1_785/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1103 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1114 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1125 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1136 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1147 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1158 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand3_1_4 sky130_fd_sc_hd__nor2_1_42/A sky130_fd_sc_hd__nand3_1_4/A
+ sky130_fd_sc_hd__nand3_1_4/C sky130_fd_sc_hd__nor3_1_0/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__decap_12_1169 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__fah_1_9 sky130_fd_sc_hd__nor2_2_29/A sky130_fd_sc_hd__fah_1_9/B
+ sky130_fd_sc_hd__fah_1_9/A sky130_fd_sc_hd__fah_1_9/SUM sky130_fd_sc_hd__fah_1_9/CI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__fah_1
Xsky130_fd_sc_hd__a222oi_1_40 vccd1 vssd1 sky130_fd_sc_hd__xor2_1_255/X sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__inv_2_59/A sky130_fd_sc_hd__xor2_1_42/X sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_40/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_51 vccd1 vssd1 sky130_fd_sc_hd__and3_1_0/X sky130_fd_sc_hd__buf_2_32/X
+ sky130_fd_sc_hd__buf_8_0/X sky130_fd_sc_hd__nor2_1_56/Y sky130_fd_sc_hd__buf_4_6/X
+ sky130_fd_sc_hd__a222oi_1_51/Y sky130_fd_sc_hd__nor2b_1_3/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__sdlclkp_2_16 sky130_fd_sc_hd__conb_1_149/LO sky130_fd_sc_hd__clkinv_4_119/A
+ sky130_fd_sc_hd__dfxtp_1_533/CLK sky130_fd_sc_hd__or2_0_113/X vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__a222oi_1_62 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__or2_0_61/A
+ sky130_fd_sc_hd__or2_0_42/B sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__or2_0_58/B
+ sky130_fd_sc_hd__a222oi_1_62/Y sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_73 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__or2_0_60/A
+ sky130_fd_sc_hd__or2_0_61/A sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__or2_0_42/B
+ sky130_fd_sc_hd__a222oi_1_73/Y sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__xnor2_1_20 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_20/B sky130_fd_sc_hd__xnor2_1_20/Y
+ sky130_fd_sc_hd__xnor2_1_20/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_660 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_84 vccd1 vssd1 sky130_fd_sc_hd__and3_4_4/X sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__buf_8_0/X sky130_fd_sc_hd__nor2_1_61/Y sky130_fd_sc_hd__buf_4_6/X
+ sky130_fd_sc_hd__a222oi_1_84/Y sky130_fd_sc_hd__nor2b_1_4/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_671 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_95 vccd1 vssd1 sky130_fd_sc_hd__and3_4_5/X sky130_fd_sc_hd__buf_4_6/X
+ sky130_fd_sc_hd__buf_4_1/X sky130_fd_sc_hd__nor2_1_68/Y sky130_fd_sc_hd__nor2_2_5/A
+ sky130_fd_sc_hd__a222oi_1_95/Y sky130_fd_sc_hd__nor2b_1_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__xnor2_1_31 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_131/A sky130_fd_sc_hd__and3_4_6/B
+ sky130_fd_sc_hd__xnor2_1_34/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_682 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_42 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_42/B sky130_fd_sc_hd__inv_2_12/A
+ sky130_fd_sc_hd__xnor2_1_42/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_693 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_53 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_55/A sky130_fd_sc_hd__and3_4_2/C
+ sky130_fd_sc_hd__xor2_1_197/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_64 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_64/B sky130_fd_sc_hd__buf_2_9/A
+ sky130_fd_sc_hd__inv_2_42/Y vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_405 sky130_fd_sc_hd__fa_2_281/A sky130_fd_sc_hd__fa_2_276/B
+ sky130_fd_sc_hd__xor2_1_405/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_75 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_77/B sky130_fd_sc_hd__and3_1_1/A
+ sky130_fd_sc_hd__xor2_1_262/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_416 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__or2_0_48/B
+ sky130_fd_sc_hd__xor2_1_416/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_86 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_86/B sky130_fd_sc_hd__xnor2_1_86/Y
+ sky130_fd_sc_hd__xnor2_1_86/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_427 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__xor3_1_23/C
+ sky130_fd_sc_hd__xor2_1_427/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_97 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_362/B sky130_fd_sc_hd__and3_4_15/C
+ sky130_fd_sc_hd__xnor2_1_97/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_438 sky130_fd_sc_hd__fa_2_338/A sky130_fd_sc_hd__fa_2_289/B
+ sky130_fd_sc_hd__xor2_1_438/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_449 sky130_fd_sc_hd__fa_2_310/A sky130_fd_sc_hd__xor2_1_449/X
+ sky130_fd_sc_hd__xor2_1_449/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1670 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a211oi_1_0 sky130_fd_sc_hd__nor2_4_1/B sky130_fd_sc_hd__ha_2_9/A
+ sky130_fd_sc_hd__inv_2_8/A sky130_fd_sc_hd__buf_2_18/A sky130_fd_sc_hd__nor2_1_40/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__decap_12_1681 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1692 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_1 sky130_fd_sc_hd__buf_12_461/A sky130_fd_sc_hd__buf_8_162/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__nor4_1_1 sky130_fd_sc_hd__nor4_1_1/D wbs_adr_i[11] sky130_fd_sc_hd__nor4_1_1/Y
+ wbs_adr_i[19] wbs_adr_i[17] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor4_1
Xsky130_fd_sc_hd__a22oi_1_0 sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__a22oi_1_0/B2 sky130_fd_sc_hd__a22oi_1_0/A2 sky130_fd_sc_hd__nand2_1_9/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__decap_12_5 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_2_16 sky130_fd_sc_hd__clkinv_2_16/Y sky130_fd_sc_hd__clkinv_4_81/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_27 sky130_fd_sc_hd__inv_2_140/A sky130_fd_sc_hd__buf_8_84/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_38 sky130_fd_sc_hd__clkinv_2_38/Y sky130_fd_sc_hd__inv_2_132/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_49 sky130_fd_sc_hd__inv_2_92/A sky130_fd_sc_hd__ha_2_32/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__or2_1_9 sky130_fd_sc_hd__or2_1_9/A sky130_fd_sc_hd__or2_1_9/X sky130_fd_sc_hd__or2_1_9/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_1
Xsky130_fd_sc_hd__buf_12_250 sky130_fd_sc_hd__buf_6_44/X sky130_fd_sc_hd__buf_12_417/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_261 sky130_fd_sc_hd__buf_12_67/X sky130_fd_sc_hd__buf_12_330/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_120 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_166/Q sky130_fd_sc_hd__dfxtp_1_134/Q sky130_fd_sc_hd__o21ai_1_26/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_272 sky130_fd_sc_hd__buf_6_88/X sky130_fd_sc_hd__buf_12_368/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_131 sky130_fd_sc_hd__xnor2_2_1/Y sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__o2bb2ai_1_0/Y sky130_fd_sc_hd__o21ai_1_41/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_283 sky130_fd_sc_hd__buf_12_283/A sky130_fd_sc_hd__buf_12_572/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_142 sky130_fd_sc_hd__xnor2_1_82/Y sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xnor2_1_19/Y sky130_fd_sc_hd__o21ai_1_64/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_294 sky130_fd_sc_hd__buf_12_294/A sky130_fd_sc_hd__buf_12_494/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_153 sky130_fd_sc_hd__xor2_1_330/X sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xor2_1_117/X sky130_fd_sc_hd__o21ai_1_85/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_164 sky130_fd_sc_hd__xnor2_1_104/Y sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xnor2_1_41/Y sky130_fd_sc_hd__a22oi_1_164/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_175 sky130_fd_sc_hd__nand2_1_131/A sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xor2_1_187/X sky130_fd_sc_hd__a22oi_1_175/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_186 sky130_fd_sc_hd__xor2_1_419/X sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xor2_1_207/X sky130_fd_sc_hd__a22oi_1_186/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_197 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__nor2b_2_2/Y sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__a22oi_1_197/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_450 sky130_fd_sc_hd__a21oi_2_10/B1 sky130_fd_sc_hd__nand2_1_384/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_461 sky130_fd_sc_hd__nor2_1_126/B sky130_fd_sc_hd__nor2_1_128/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_472 sky130_fd_sc_hd__a21oi_1_89/B1 sky130_fd_sc_hd__nand2_1_435/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_483 sky130_fd_sc_hd__nand2_1_441/A sky130_fd_sc_hd__nor2_1_147/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_494 sky130_fd_sc_hd__a21oi_1_96/B1 sky130_fd_sc_hd__nand2_1_466/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_408 vssd1 vccd1 sky130_fd_sc_hd__inv_2_36/Y sky130_fd_sc_hd__nand2b_1_8/Y
+ sky130_fd_sc_hd__o21ai_1_408/B1 sky130_fd_sc_hd__xor2_1_219/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_419 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_486/A2 sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_419/B1 sky130_fd_sc_hd__xor2_1_228/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2_4_17 sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__nor2_4_17/A
+ sky130_fd_sc_hd__nor2_4_17/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__nand2_2_10 sky130_fd_sc_hd__nor2_4_4/B sky130_fd_sc_hd__nor2_1_40/A
+ sky130_fd_sc_hd__nand2_2_11/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__decap_12_490 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_202 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__or2_0_22/B
+ sky130_fd_sc_hd__xor2_1_202/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_213 sky130_fd_sc_hd__xor2_1_213/B sky130_fd_sc_hd__xor2_2_1/A
+ sky130_fd_sc_hd__xor3_1_10/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_224 sky130_fd_sc_hd__xor2_1_362/B sky130_fd_sc_hd__xor2_1_224/X
+ sky130_fd_sc_hd__xor2_1_224/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_235 sky130_fd_sc_hd__fa_2_239/A sky130_fd_sc_hd__xor2_1_235/X
+ sky130_fd_sc_hd__xor2_1_235/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_246 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__fa_2_162/B
+ sky130_fd_sc_hd__xor2_1_246/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_257 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__fa_2_169/B
+ sky130_fd_sc_hd__xor2_1_257/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_268 sky130_fd_sc_hd__fa_2_239/A sky130_fd_sc_hd__fa_2_180/B
+ sky130_fd_sc_hd__xor2_1_268/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_279 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__xor2_1_279/X
+ sky130_fd_sc_hd__xor2_1_279/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_206 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_254/A sky130_fd_sc_hd__clkbuf_1_53/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_217 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_43/A sky130_fd_sc_hd__clkinv_1_902/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_228 vssd1 vccd1 sky130_fd_sc_hd__buf_8_61/A sky130_fd_sc_hd__clkbuf_4_34/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o21ai_1_920 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_280/Y la_data_out[51]
+ sky130_fd_sc_hd__a21oi_1_196/Y sky130_fd_sc_hd__o21ai_1_920/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_1_239 vssd1 vccd1 sky130_fd_sc_hd__buf_8_107/A sky130_fd_sc_hd__clkbuf_1_296/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_8_2 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__buf_2_40 vccd1 vssd1 sky130_fd_sc_hd__buf_2_40/X sky130_fd_sc_hd__buf_2_40/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_51 vccd1 vssd1 sky130_fd_sc_hd__buf_2_51/X sky130_fd_sc_hd__buf_2_51/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_62 vccd1 vssd1 sky130_fd_sc_hd__mux2_8_1/S sky130_fd_sc_hd__mux2_8_0/S
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_73 vccd1 vssd1 sky130_fd_sc_hd__buf_2_73/X sky130_fd_sc_hd__buf_2_73/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_84 vccd1 vssd1 sky130_fd_sc_hd__buf_2_84/X sky130_fd_sc_hd__buf_2_84/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_95 vccd1 vssd1 sky130_fd_sc_hd__buf_2_95/X sky130_fd_sc_hd__buf_2_95/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__diode_2_2 sky130_fd_sc_hd__clkbuf_4_20/X vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__and2_0_204 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_83/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_79/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_215 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_53/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_70/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_226 vccd1 vssd1 sky130_fd_sc_hd__and2_0_226/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_226/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_237 vccd1 vssd1 sky130_fd_sc_hd__and2_0_237/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_53/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_248 vccd1 vssd1 sky130_fd_sc_hd__and2_0_248/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_248/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_259 vccd1 vssd1 sky130_fd_sc_hd__and2_0_259/X sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__and2_0_259/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__xor3_1_13 sky130_fd_sc_hd__xor3_1_13/X sky130_fd_sc_hd__xor3_1_13/C
+ sky130_fd_sc_hd__xor3_1_14/X sky130_fd_sc_hd__xor3_1_13/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__xor3_1_24 sky130_fd_sc_hd__xor3_1_24/X sky130_fd_sc_hd__xor3_1_24/C
+ sky130_fd_sc_hd__xor3_1_24/B sky130_fd_sc_hd__xor3_1_25/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__sdlclkp_2_9 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_8_1/Y
+ sky130_fd_sc_hd__dfxtp_1_217/CLK sky130_fd_sc_hd__o21ai_2_2/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__a22o_2_3 sky130_fd_sc_hd__nand2_1_7/B sky130_fd_sc_hd__fa_2_419/A
+ sky130_fd_sc_hd__or2_0_42/B sky130_fd_sc_hd__fa_2_419/B sky130_fd_sc_hd__nand2_1_8/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_2
Xsky130_fd_sc_hd__clkinv_1_280 sky130_fd_sc_hd__and2_0_115/A sky130_fd_sc_hd__a222oi_1_24/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_291 sky130_fd_sc_hd__and2_0_184/A sky130_fd_sc_hd__a222oi_1_35/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkbuf_4_12 sky130_fd_sc_hd__buf_2_67/A sky130_fd_sc_hd__buf_6_7/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_205 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_241/A2 sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__a222oi_1_79/Y sky130_fd_sc_hd__xor2_1_32/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_23 sky130_fd_sc_hd__buf_2_52/A sky130_fd_sc_hd__inv_8_0/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_216 vssd1 vccd1 sky130_fd_sc_hd__inv_2_17/Y sky130_fd_sc_hd__nand2b_1_6/Y
+ sky130_fd_sc_hd__a222oi_1_87/Y sky130_fd_sc_hd__xor2_1_41/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_34 sky130_fd_sc_hd__clkbuf_4_34/X sky130_fd_sc_hd__buf_8_55/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_227 vssd1 vccd1 sky130_fd_sc_hd__buf_2_1/X sky130_fd_sc_hd__nand2b_1_5/Y
+ sky130_fd_sc_hd__a222oi_1_95/Y sky130_fd_sc_hd__xor2_1_52/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_45 sky130_fd_sc_hd__buf_2_45/A wbs_dat_i[10] vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_238 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_2/X sky130_fd_sc_hd__nand2_1_192/Y
+ sky130_fd_sc_hd__a21oi_1_43/Y sky130_fd_sc_hd__xnor2_1_16/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_249 vssd1 vccd1 sky130_fd_sc_hd__inv_2_22/Y sky130_fd_sc_hd__nand2b_2_0/Y
+ sky130_fd_sc_hd__o21ai_1_249/B1 sky130_fd_sc_hd__xor2_1_72/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__buf_8_140 sky130_fd_sc_hd__inv_2_112/Y sky130_fd_sc_hd__buf_8_140/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nand2_1_609 sky130_fd_sc_hd__nand2_1_609/Y sky130_fd_sc_hd__nand2_1_615/A
+ sky130_fd_sc_hd__nor2_1_201/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__buf_8_151 sky130_fd_sc_hd__buf_8_151/A sky130_fd_sc_hd__buf_8_151/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nor2_4_2 sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__ha_2_8/A sky130_fd_sc_hd__nor2_4_2/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__buf_8_162 sky130_fd_sc_hd__buf_8_162/A sky130_fd_sc_hd__buf_8_162/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_405 sky130_fd_sc_hd__dfxtp_1_405/Q sky130_fd_sc_hd__dfxtp_1_410/CLK
+ sky130_fd_sc_hd__nor2b_1_110/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_416 sky130_fd_sc_hd__dfxtp_1_416/Q sky130_fd_sc_hd__dfxtp_1_417/CLK
+ sky130_fd_sc_hd__nor2b_1_99/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_427 sky130_fd_sc_hd__dfxtp_1_427/Q sky130_fd_sc_hd__dfxtp_1_427/CLK
+ sky130_fd_sc_hd__nor2b_1_89/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_438 sky130_fd_sc_hd__dfxtp_1_438/Q sky130_fd_sc_hd__dfxtp_1_439/CLK
+ sky130_fd_sc_hd__nor2b_1_109/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_449 sky130_fd_sc_hd__dfxtp_1_449/Q sky130_fd_sc_hd__dfxtp_1_451/CLK
+ sky130_fd_sc_hd__nor2b_1_98/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a222oi_1_107 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__or2_0_60/B
+ sky130_fd_sc_hd__or2_0_60/A sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__or2_0_61/A
+ sky130_fd_sc_hd__o21ai_1_241/B1 sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2b_1_19 sky130_fd_sc_hd__nand2b_1_19/Y sky130_fd_sc_hd__and3_4_23/C
+ sky130_fd_sc_hd__and3_4_23/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a222oi_1_118 vccd1 vssd1 sky130_fd_sc_hd__and3_4_8/X sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__buf_6_1/X sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__o21ai_1_256/B1 sky130_fd_sc_hd__nor2b_2_2/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__o21ai_1_750 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_771/A2 sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_750/B1 sky130_fd_sc_hd__xor2_1_525/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_129 vccd1 vssd1 sky130_fd_sc_hd__and3_4_6/X sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__buf_4_6/X sky130_fd_sc_hd__nor2_1_72/Y sky130_fd_sc_hd__buf_4_1/X
+ sky130_fd_sc_hd__o21ai_1_269/B1 sky130_fd_sc_hd__nor2b_1_6/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__o21ai_1_761 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_126/Y sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_761/B1 sky130_fd_sc_hd__xor2_1_536/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_772 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_10/X sky130_fd_sc_hd__nor2_1_182/B
+ sky130_fd_sc_hd__o21ai_1_772/B1 sky130_fd_sc_hd__xnor2_1_156/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_783 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_861/A2 sky130_fd_sc_hd__nand2b_1_21/Y
+ sky130_fd_sc_hd__nand2_1_496/Y sky130_fd_sc_hd__xor2_1_556/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_794 vssd1 vccd1 sky130_fd_sc_hd__nand2_2_13/Y sky130_fd_sc_hd__nand2b_1_15/Y
+ sky130_fd_sc_hd__a22oi_1_218/Y sky130_fd_sc_hd__xor2_1_568/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkinv_8_15 sky130_fd_sc_hd__clkinv_8_17/A sky130_fd_sc_hd__clkinv_8_15/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_26 sky130_fd_sc_hd__clkinv_8_26/Y sky130_fd_sc_hd__clkinv_8_28/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_37 sky130_fd_sc_hd__clkinv_8_38/A sky130_fd_sc_hd__clkinv_8_39/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_48 sky130_fd_sc_hd__clkinv_8_49/A sky130_fd_sc_hd__clkinv_8_48/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_59 sky130_fd_sc_hd__clkinv_8_2/A sky130_fd_sc_hd__clkinv_8_62/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_13 sky130_fd_sc_hd__buf_12_13/A sky130_fd_sc_hd__buf_12_13/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_24 sky130_fd_sc_hd__inv_2_125/Y sky130_fd_sc_hd__buf_12_24/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_35 sky130_fd_sc_hd__inv_2_170/Y sky130_fd_sc_hd__buf_12_35/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_90 sky130_fd_sc_hd__fa_2_75/A sky130_fd_sc_hd__xor2_1_90/X
+ sky130_fd_sc_hd__xor2_1_90/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_46 sky130_fd_sc_hd__buf_12_46/A sky130_fd_sc_hd__buf_12_46/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_57 sky130_fd_sc_hd__buf_12_57/A sky130_fd_sc_hd__buf_12_57/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_68 sky130_fd_sc_hd__buf_8_100/X sky130_fd_sc_hd__buf_12_68/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_79 sky130_fd_sc_hd__buf_6_19/X sky130_fd_sc_hd__buf_12_79/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_2_8 vccd1 vssd1 sky130_fd_sc_hd__buf_2_8/X sky130_fd_sc_hd__buf_2_8/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o21ai_2_11 sky130_fd_sc_hd__o21ai_2_11/B1 sky130_fd_sc_hd__xnor2_1_73/B
+ sky130_fd_sc_hd__a21oi_2_8/Y sky130_fd_sc_hd__nor2_2_11/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__o21ai_2
Xsky130_fd_sc_hd__inv_2_8 sky130_fd_sc_hd__inv_2_8/A sky130_fd_sc_hd__inv_2_8/Y vccd1
+ vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__nor2_1_18 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_18/Y
+ sky130_fd_sc_hd__nor2_1_18/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_29 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_29/Y
+ sky130_fd_sc_hd__nor2_1_29/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__and2_0_40 vccd1 vssd1 sky130_fd_sc_hd__and2_0_40/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__nor2_2_10/B vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_51 vccd1 vssd1 sky130_fd_sc_hd__and2_0_51/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__nor2_1_85/B vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_62 vccd1 vssd1 sky130_fd_sc_hd__and2_0_62/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__or2_0_66/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_73 vccd1 vssd1 sky130_fd_sc_hd__and2_0_73/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__buf_4_3/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_406 sky130_fd_sc_hd__nand2_1_406/Y sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__nor2_1_73/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_84 vccd1 vssd1 sky130_fd_sc_hd__and2_0_84/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__buf_4_2/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_417 sky130_fd_sc_hd__xnor2_1_100/A sky130_fd_sc_hd__nand2_1_418/Y
+ sky130_fd_sc_hd__nand2_1_417/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_95 vccd1 vssd1 sky130_fd_sc_hd__and2_0_95/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__or2_0_58/B vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_428 sky130_fd_sc_hd__xnor2_1_103/A sky130_fd_sc_hd__nand2_1_429/Y
+ sky130_fd_sc_hd__nand2_1_428/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_439 sky130_fd_sc_hd__xnor2_1_108/A sky130_fd_sc_hd__nand2_1_440/Y
+ sky130_fd_sc_hd__nand2_1_439/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_19 sky130_fd_sc_hd__or2_0_84/A sky130_fd_sc_hd__fa_2_432/A
+ sky130_fd_sc_hd__nor2b_1_19/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1008 sky130_fd_sc_hd__clkinv_1_1009/A sky130_fd_sc_hd__inv_2_1/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_50 sky130_fd_sc_hd__buf_8_50/A sky130_fd_sc_hd__buf_8_50/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__clkinv_1_1019 sky130_fd_sc_hd__clkinv_1_1019/Y sky130_fd_sc_hd__clkinv_1_1019/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_61 sky130_fd_sc_hd__buf_8_61/A sky130_fd_sc_hd__buf_8_61/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_72 sky130_fd_sc_hd__buf_8_72/A sky130_fd_sc_hd__buf_8_72/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_83 sky130_fd_sc_hd__buf_8_83/A sky130_fd_sc_hd__buf_8_83/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_202 sky130_fd_sc_hd__xor2_1_575/A sky130_fd_sc_hd__dfxtp_2_2/CLK
+ sky130_fd_sc_hd__and2_0_78/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_8_94 sky130_fd_sc_hd__buf_8_94/A sky130_fd_sc_hd__buf_8_94/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_213 sky130_fd_sc_hd__xnor2_1_140/B sky130_fd_sc_hd__dfxtp_1_217/CLK
+ sky130_fd_sc_hd__and2_0_95/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_224 sky130_fd_sc_hd__xnor2_1_114/A sky130_fd_sc_hd__dfxtp_2_4/CLK
+ sky130_fd_sc_hd__and2_0_56/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_235 sky130_fd_sc_hd__fa_2_239/A sky130_fd_sc_hd__dfxtp_2_5/CLK
+ sky130_fd_sc_hd__and2_0_75/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_246 sky130_fd_sc_hd__xnor2_1_68/A sky130_fd_sc_hd__clkinv_4_4/Y
+ sky130_fd_sc_hd__and2_0_58/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_257 sky130_fd_sc_hd__xor2_1_170/A sky130_fd_sc_hd__dfxtp_1_269/CLK
+ sky130_fd_sc_hd__and2_0_47/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_268 sky130_fd_sc_hd__xnor2_1_21/A sky130_fd_sc_hd__dfxtp_1_269/CLK
+ sky130_fd_sc_hd__and2_0_67/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_279 sky130_fd_sc_hd__dfxtp_1_279/Q sky130_fd_sc_hd__dfxtp_1_2/CLK
+ sky130_fd_sc_hd__and2_0_255/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_580 vssd1 vccd1 sky130_fd_sc_hd__buf_2_8/X sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_580/B1 sky130_fd_sc_hd__xor2_1_375/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_107 sky130_fd_sc_hd__fa_2_103/A sky130_fd_sc_hd__fa_2_108/A
+ sky130_fd_sc_hd__fa_2_107/A sky130_fd_sc_hd__fa_2_107/B sky130_fd_sc_hd__xor2_1_144/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o21ai_1_591 vssd1 vccd1 sky130_fd_sc_hd__inv_2_42/Y sky130_fd_sc_hd__o21ai_1_591/A1
+ sky130_fd_sc_hd__o21ai_1_591/B1 sky130_fd_sc_hd__xnor2_1_110/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_118 sky130_fd_sc_hd__fa_2_113/B sky130_fd_sc_hd__fa_2_116/A
+ sky130_fd_sc_hd__fa_2_118/A sky130_fd_sc_hd__fa_2_118/B sky130_fd_sc_hd__fa_2_118/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_129 sky130_fd_sc_hd__nor2_1_88/A sky130_fd_sc_hd__nor2_1_91/B
+ sky130_fd_sc_hd__fa_2_129/A sky130_fd_sc_hd__fa_2_129/B sky130_fd_sc_hd__fa_2_129/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_102 vccd1 vssd1 sky130_fd_sc_hd__buf_2_102/X sky130_fd_sc_hd__buf_2_102/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_113 vccd1 vssd1 sky130_fd_sc_hd__buf_2_113/X sky130_fd_sc_hd__buf_2_113/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_124 vccd1 vssd1 sky130_fd_sc_hd__buf_2_124/X sky130_fd_sc_hd__buf_2_124/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_17 sky130_fd_sc_hd__o22ai_1_46/B1 sky130_fd_sc_hd__o22ai_1_17/B1
+ sky130_fd_sc_hd__o22ai_1_17/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__inv_4_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_135 vccd1 vssd1 sky130_fd_sc_hd__buf_2_135/X sky130_fd_sc_hd__inv_2_0/Y
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_28 sky130_fd_sc_hd__o22ai_1_33/B1 sky130_fd_sc_hd__o21ai_1_3/A2
+ sky130_fd_sc_hd__o22ai_1_28/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__inv_4_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_146 vccd1 vssd1 sky130_fd_sc_hd__buf_2_146/X sky130_fd_sc_hd__buf_2_146/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_39 sky130_fd_sc_hd__nor2_1_35/A sky130_fd_sc_hd__o22ai_1_39/B1
+ sky130_fd_sc_hd__o22ai_1_39/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__nor2_4_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_157 vccd1 vssd1 sky130_fd_sc_hd__buf_2_157/X sky130_fd_sc_hd__buf_2_157/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_168 vccd1 vssd1 la_data_out[55] sky130_fd_sc_hd__ha_2_33/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_179 vccd1 vssd1 la_data_out[32] sky130_fd_sc_hd__nor4b_2_0/Y
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__ha_2_2 vssd1 vccd1 sky130_fd_sc_hd__ha_2_2/A sky130_fd_sc_hd__xor3_1_25/C
+ sky130_fd_sc_hd__ha_2_2/SUM sky130_fd_sc_hd__ha_2_2/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__buf_4_19 vccd1 vssd1 sky130_fd_sc_hd__buf_4_19/X sky130_fd_sc_hd__buf_4_19/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__a222oi_1_460 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__buf_4_5/X sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__o21ai_1_742/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_471 vccd1 vssd1 sky130_fd_sc_hd__and3_4_26/X sky130_fd_sc_hd__buf_2_30/X
+ sky130_fd_sc_hd__buf_2_26/X sky130_fd_sc_hd__nor2_2_31/Y sky130_fd_sc_hd__buf_2_24/X
+ sky130_fd_sc_hd__o21ai_1_758/B1 sky130_fd_sc_hd__nor2b_1_12/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_13 vssd1 vccd1 sky130_fd_sc_hd__nand2_1_135/A sky130_fd_sc_hd__xnor2_1_117/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_482 vccd1 vssd1 sky130_fd_sc_hd__and3_4_21/X sky130_fd_sc_hd__buf_2_21/X
+ sky130_fd_sc_hd__nor2_1_87/A sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__o21ai_1_770/B1 sky130_fd_sc_hd__and2b_4_12/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_24 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_24/X sky130_fd_sc_hd__nor2_4_2/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_493 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__buf_6_4/X
+ sky130_fd_sc_hd__buf_6_0/X sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__o21ai_1_785/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_35 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_35/X la_data_out[44]
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_46 vssd1 vccd1 sky130_fd_sc_hd__nand2_2_14/A sky130_fd_sc_hd__clkbuf_1_46/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_57 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_57/X sky130_fd_sc_hd__clkbuf_1_60/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_68 vssd1 vccd1 sky130_fd_sc_hd__mux2_4_5/A1 sky130_fd_sc_hd__clkbuf_1_68/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_79 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_6/A1 sky130_fd_sc_hd__clkbuf_1_79/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__or2_0_15 sky130_fd_sc_hd__or2_0_61/A sky130_fd_sc_hd__or2_0_15/X
+ sky130_fd_sc_hd__or2_0_42/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_26 sky130_fd_sc_hd__or2_0_53/A sky130_fd_sc_hd__or2_0_26/X
+ sky130_fd_sc_hd__inv_6_0/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_37 sky130_fd_sc_hd__or2_0_37/A sky130_fd_sc_hd__or2_0_37/X
+ sky130_fd_sc_hd__or2_0_37/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_48 sky130_fd_sc_hd__or2_0_48/A sky130_fd_sc_hd__or2_0_48/X
+ sky130_fd_sc_hd__or2_0_48/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_59 sky130_fd_sc_hd__or2_0_66/A sky130_fd_sc_hd__or2_0_59/X
+ sky130_fd_sc_hd__or2_0_60/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__buf_12_2 sky130_fd_sc_hd__buf_12_2/A sky130_fd_sc_hd__buf_12_2/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_602 sky130_fd_sc_hd__buf_12_602/A sky130_fd_sc_hd__buf_12_602/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_613 sky130_fd_sc_hd__buf_12_613/A sky130_fd_sc_hd__buf_12_613/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_624 sky130_fd_sc_hd__buf_12_624/A sky130_fd_sc_hd__buf_12_624/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_635 sky130_fd_sc_hd__buf_12_635/A sky130_fd_sc_hd__buf_12_635/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_4_106 sky130_fd_sc_hd__clkinv_8_65/Y sky130_fd_sc_hd__clkinv_2_60/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_12_646 sky130_fd_sc_hd__buf_12_646/A sky130_fd_sc_hd__buf_12_646/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_4_117 sky130_fd_sc_hd__clkinv_4_117/A sky130_fd_sc_hd__clkinv_8_74/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_12_657 sky130_fd_sc_hd__buf_12_657/A sky130_fd_sc_hd__buf_12_657/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_668 sky130_fd_sc_hd__buf_12_668/A sky130_fd_sc_hd__buf_12_668/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_679 sky130_fd_sc_hd__buf_12_679/A sky130_fd_sc_hd__buf_12_679/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_308 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_319 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_203 sky130_fd_sc_hd__nand2_1_203/Y sky130_fd_sc_hd__or2_0_13/X
+ sky130_fd_sc_hd__nand2_1_203/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_802 sky130_fd_sc_hd__and2_0_305/A sky130_fd_sc_hd__clkinv_1_802/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_214 sky130_fd_sc_hd__nand2_1_214/Y sky130_fd_sc_hd__or2_0_17/X
+ sky130_fd_sc_hd__nor2_1_67/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_813 sky130_fd_sc_hd__nand2_1_804/A sky130_fd_sc_hd__nor2_1_257/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_225 sky130_fd_sc_hd__xnor2_1_29/A sky130_fd_sc_hd__nand2_1_226/Y
+ sky130_fd_sc_hd__or2_0_19/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_824 sky130_fd_sc_hd__clkinv_1_824/Y sky130_fd_sc_hd__nand2_1_827/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_236 sky130_fd_sc_hd__xor2_1_133/B sky130_fd_sc_hd__nand2_1_237/Y
+ sky130_fd_sc_hd__nand2_1_236/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_835 sky130_fd_sc_hd__inv_2_72/A sky130_fd_sc_hd__ha_2_35/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_247 sky130_fd_sc_hd__nand2_1_247/Y sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__buf_6_4/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_846 sky130_fd_sc_hd__buf_2_36/A sky130_fd_sc_hd__clkinv_1_846/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_258 sky130_fd_sc_hd__nand2_1_258/Y sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__nor2_2_10/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_857 sky130_fd_sc_hd__clkinv_1_857/Y sky130_fd_sc_hd__inv_2_195/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_269 sky130_fd_sc_hd__nand2_1_269/Y sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__buf_6_1/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_868 sky130_fd_sc_hd__clkinv_1_868/Y sky130_fd_sc_hd__inv_2_95/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_879 sky130_fd_sc_hd__clkinv_1_879/Y sky130_fd_sc_hd__inv_4_15/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__conb_1_13 sky130_fd_sc_hd__conb_1_13/LO sky130_fd_sc_hd__conb_1_13/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_24 sky130_fd_sc_hd__conb_1_24/LO sky130_fd_sc_hd__conb_1_24/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_35 sky130_fd_sc_hd__conb_1_35/LO sky130_fd_sc_hd__conb_1_35/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1307 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_46 sky130_fd_sc_hd__conb_1_46/LO sky130_fd_sc_hd__conb_1_46/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1318 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_57 sky130_fd_sc_hd__conb_1_57/LO sky130_fd_sc_hd__conb_1_57/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1329 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_68 sky130_fd_sc_hd__conb_1_68/LO sky130_fd_sc_hd__conb_1_68/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_79 sky130_fd_sc_hd__conb_1_79/LO sky130_fd_sc_hd__conb_1_79/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__mux2_2_8 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_8/A1 sky130_fd_sc_hd__buf_2_82/X
+ sky130_fd_sc_hd__mux2_8_0/S sky130_fd_sc_hd__mux2_2_8/X vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__decap_12_820 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_831 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_842 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_853 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_864 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_875 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_886 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_770 sky130_fd_sc_hd__nand2_1_770/Y sky130_fd_sc_hd__nor2_1_253/A
+ sky130_fd_sc_hd__nor2_1_253/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_897 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_781 sky130_fd_sc_hd__nand2_1_781/Y sky130_fd_sc_hd__nor2_1_252/A
+ sky130_fd_sc_hd__nor2_1_252/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_609 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__nor2_4_16/B
+ sky130_fd_sc_hd__xor2_1_609/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_792 sky130_fd_sc_hd__xor2_1_676/B sky130_fd_sc_hd__nand2_1_793/Y
+ sky130_fd_sc_hd__nand2_1_792/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_1830 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1841 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1852 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1863 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_290 vccd1 vssd1 sky130_fd_sc_hd__and3_4_16/X sky130_fd_sc_hd__buf_4_0/X
+ sky130_fd_sc_hd__buf_2_23/X sky130_fd_sc_hd__nor2_2_19/Y sky130_fd_sc_hd__buf_2_31/X
+ sky130_fd_sc_hd__o21ai_1_500/B1 sky130_fd_sc_hd__nor2b_2_3/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_460 sky130_fd_sc_hd__xor2_1_674/B sky130_fd_sc_hd__fa_2_460/SUM
+ sky130_fd_sc_hd__fa_2_460/A sky130_fd_sc_hd__fa_2_460/B sky130_fd_sc_hd__fa_2_460/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_471 sky130_fd_sc_hd__or2_0_100/B sky130_fd_sc_hd__nor2_1_255/A
+ sky130_fd_sc_hd__fa_2_471/A sky130_fd_sc_hd__fa_2_471/B sky130_fd_sc_hd__nor2b_1_41/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_482 sky130_fd_sc_hd__nor2_1_260/B sky130_fd_sc_hd__or2_0_106/A
+ sky130_fd_sc_hd__fa_2_482/A sky130_fd_sc_hd__fa_2_482/B sky130_fd_sc_hd__nor2b_1_63/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_1_109 io_oeb[30] sky130_fd_sc_hd__conb_1_33/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_9 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_9/A2 sky130_fd_sc_hd__nor2_4_4/B
+ sky130_fd_sc_hd__o21ai_1_9/B1 sky130_fd_sc_hd__xor3_1_5/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_8_10 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__nor2_1_203 sky130_fd_sc_hd__nor2_1_203/B sky130_fd_sc_hd__nor2_1_203/Y
+ sky130_fd_sc_hd__nor2_1_203/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_214 sky130_fd_sc_hd__buf_2_26/X sky130_fd_sc_hd__nor2_1_214/Y
+ sky130_fd_sc_hd__buf_2_24/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_225 sky130_fd_sc_hd__mux2_2_37/X sky130_fd_sc_hd__nor2_1_225/Y
+ sky130_fd_sc_hd__mux2_2_18/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_236 sky130_fd_sc_hd__nor2_1_237/Y sky130_fd_sc_hd__nor2_1_236/Y
+ sky130_fd_sc_hd__nor2_1_238/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_247 sky130_fd_sc_hd__nor2_1_247/B sky130_fd_sc_hd__nor2_1_247/Y
+ sky130_fd_sc_hd__nor2_1_247/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_258 sky130_fd_sc_hd__nor2_1_258/B sky130_fd_sc_hd__nor2_1_258/Y
+ sky130_fd_sc_hd__nor2_1_258/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_269 sky130_fd_sc_hd__nor2_1_271/Y sky130_fd_sc_hd__nor2_1_269/Y
+ sky130_fd_sc_hd__and2_4_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_410 sky130_fd_sc_hd__buf_12_93/X sky130_fd_sc_hd__buf_12_486/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_421 sky130_fd_sc_hd__buf_12_421/A sky130_fd_sc_hd__buf_12_495/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_432 sky130_fd_sc_hd__buf_12_432/A sky130_fd_sc_hd__buf_12_643/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_443 sky130_fd_sc_hd__buf_12_443/A sky130_fd_sc_hd__buf_12_443/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_454 sky130_fd_sc_hd__buf_12_454/A sky130_fd_sc_hd__buf_12_454/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_465 sky130_fd_sc_hd__buf_12_465/A sky130_fd_sc_hd__buf_12_665/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_476 sky130_fd_sc_hd__buf_12_476/A sky130_fd_sc_hd__buf_12_476/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_105 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_487 sky130_fd_sc_hd__buf_12_487/A sky130_fd_sc_hd__buf_12_552/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_116 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_498 sky130_fd_sc_hd__buf_12_498/A sky130_fd_sc_hd__buf_12_668/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_127 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_138 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_610 sky130_fd_sc_hd__nand2_1_654/A sky130_fd_sc_hd__nor2_1_219/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_149 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_621 sky130_fd_sc_hd__o21ai_1_41/A2 sky130_fd_sc_hd__buf_2_22/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_632 sky130_fd_sc_hd__nand2_1_676/A sky130_fd_sc_hd__nor2_1_224/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_643 sky130_fd_sc_hd__clkinv_1_643/Y sky130_fd_sc_hd__nand2_1_699/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_206 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_206/B sky130_fd_sc_hd__a22o_1_18/B1
+ sky130_fd_sc_hd__xnor2_1_206/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_654 sky130_fd_sc_hd__o22ai_1_92/B1 sky130_fd_sc_hd__buf_2_207/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_217 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_217/B sky130_fd_sc_hd__nor2_1_240/B
+ sky130_fd_sc_hd__xnor2_1_217/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_665 sky130_fd_sc_hd__nand2_1_732/A sky130_fd_sc_hd__nor2_1_237/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_228 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_5/B sky130_fd_sc_hd__xnor2_1_228/Y
+ la_data_out[71] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_676 sky130_fd_sc_hd__clkinv_1_676/Y sky130_fd_sc_hd__nand2_1_754/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_239 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_5/B sky130_fd_sc_hd__xnor2_1_239/Y
+ sky130_fd_sc_hd__or2_0_82/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_687 sky130_fd_sc_hd__xnor2_1_215/B sky130_fd_sc_hd__a21oi_1_166/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_698 sky130_fd_sc_hd__xnor2_1_218/A sky130_fd_sc_hd__and2_0_302/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1104 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1115 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1126 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1137 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1148 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1159 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand3_1_5 sky130_fd_sc_hd__nand3_1_5/Y la_data_out[36] sky130_fd_sc_hd__nand3_1_5/C
+ sky130_fd_sc_hd__nand3_1_5/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__a222oi_1_30 vccd1 vssd1 sky130_fd_sc_hd__xor2_1_330/X sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__xor2_1_543/X sky130_fd_sc_hd__xor2_1_117/X sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_30/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_41 vccd1 vssd1 sky130_fd_sc_hd__xnor2_1_78/Y sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__xnor2_1_141/Y sky130_fd_sc_hd__xnor2_1_15/Y sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_41/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_52 vccd1 vssd1 sky130_fd_sc_hd__and3_4_6/X sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__nor2_1_87/A sky130_fd_sc_hd__nor2_1_72/Y sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__a222oi_1_52/Y sky130_fd_sc_hd__nor2b_1_6/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_63 vccd1 vssd1 sky130_fd_sc_hd__and3_4_2/X sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__or2_0_60/B sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__or2_0_60/A
+ sky130_fd_sc_hd__a222oi_1_63/Y sky130_fd_sc_hd__and2b_4_4/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_650 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_74 vccd1 vssd1 sky130_fd_sc_hd__and3_4_1/X sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__buf_4_2/X sky130_fd_sc_hd__nor2_2_9/Y sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__a222oi_1_74/Y sky130_fd_sc_hd__and2b_4_3/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__xnor2_1_10 vssd1 vccd1 sky130_fd_sc_hd__o21ai_2_5/Y sky130_fd_sc_hd__xnor2_1_10/Y
+ sky130_fd_sc_hd__xnor2_1_10/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_661 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_85 vccd1 vssd1 sky130_fd_sc_hd__and3_4_8/X sky130_fd_sc_hd__nor2_2_10/B
+ sky130_fd_sc_hd__buf_6_4/X sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__a222oi_1_85/Y sky130_fd_sc_hd__nor2b_2_2/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__xnor2_1_21 vssd1 vccd1 sky130_fd_sc_hd__fa_2_75/A sky130_fd_sc_hd__and3_4_4/C
+ sky130_fd_sc_hd__xnor2_1_21/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_672 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_96 vccd1 vssd1 sky130_fd_sc_hd__and3_4_6/X sky130_fd_sc_hd__nor2_2_5/B
+ sky130_fd_sc_hd__nor2_2_4/B sky130_fd_sc_hd__nor2_1_72/Y sky130_fd_sc_hd__buf_2_4/X
+ sky130_fd_sc_hd__a222oi_1_96/Y sky130_fd_sc_hd__nor2b_1_6/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__xnor2_1_32 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_32/B sky130_fd_sc_hd__xnor2_1_32/Y
+ sky130_fd_sc_hd__xnor2_1_32/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_683 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_43 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_170/A sky130_fd_sc_hd__and3_4_8/B
+ sky130_fd_sc_hd__xnor2_1_46/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_54 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_54/B sky130_fd_sc_hd__xnor2_1_54/Y
+ sky130_fd_sc_hd__xnor2_1_54/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_694 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_65 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_65/B sky130_fd_sc_hd__buf_2_11/A
+ sky130_fd_sc_hd__xnor2_1_65/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_406 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__fa_2_275/B
+ sky130_fd_sc_hd__xor2_1_406/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_76 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_76/B sky130_fd_sc_hd__xnor2_1_76/Y
+ sky130_fd_sc_hd__xnor2_1_76/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_417 sky130_fd_sc_hd__fa_2_281/A sky130_fd_sc_hd__xor2_1_417/X
+ sky130_fd_sc_hd__xor2_1_417/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_87 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_87/B sky130_fd_sc_hd__xnor2_1_87/Y
+ sky130_fd_sc_hd__xnor2_1_87/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_428 sky130_fd_sc_hd__fa_2_338/A sky130_fd_sc_hd__xor3_1_24/C
+ sky130_fd_sc_hd__xor2_1_428/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_98 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_98/B sky130_fd_sc_hd__xnor2_1_98/Y
+ sky130_fd_sc_hd__xnor2_1_98/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_439 sky130_fd_sc_hd__fa_2_357/A sky130_fd_sc_hd__fa_2_289/A
+ sky130_fd_sc_hd__xor2_1_439/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1660 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1671 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1682 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1693 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_2 sky130_fd_sc_hd__buf_12_460/A sky130_fd_sc_hd__buf_4_32/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__fa_2_290 sky130_fd_sc_hd__xor3_1_26/B sky130_fd_sc_hd__fa_2_290/SUM
+ sky130_fd_sc_hd__fa_2_290/A sky130_fd_sc_hd__fa_2_290/B sky130_fd_sc_hd__fa_2_290/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor4_1_2 wbs_adr_i[1] wbs_adr_i[13] sky130_fd_sc_hd__nor4_1_2/Y
+ wbs_adr_i[30] wbs_adr_i[31] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor4_1
Xsky130_fd_sc_hd__a22oi_1_1 sky130_fd_sc_hd__nor2_4_0/Y sky130_fd_sc_hd__nor2_2_0/Y
+ sky130_fd_sc_hd__a22oi_1_1/B2 sky130_fd_sc_hd__nor2_1_234/A sky130_fd_sc_hd__nand2_1_9/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__decap_12_6 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_2_17 sky130_fd_sc_hd__clkinv_2_17/Y sky130_fd_sc_hd__clkinv_4_88/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_28 sky130_fd_sc_hd__inv_2_141/A sky130_fd_sc_hd__buf_8_26/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_39 sky130_fd_sc_hd__clkinv_2_39/Y sky130_fd_sc_hd__inv_2_144/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__buf_12_240 sky130_fd_sc_hd__buf_6_29/X sky130_fd_sc_hd__buf_12_405/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_251 sky130_fd_sc_hd__buf_6_76/X sky130_fd_sc_hd__buf_12_343/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_110 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_176/Q sky130_fd_sc_hd__dfxtp_1_144/Q sky130_fd_sc_hd__o21ai_1_16/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_262 sky130_fd_sc_hd__buf_8_159/X sky130_fd_sc_hd__buf_12_301/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_121 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_165/Q sky130_fd_sc_hd__dfxtp_1_133/Q sky130_fd_sc_hd__o21ai_1_27/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_273 sky130_fd_sc_hd__buf_6_90/X sky130_fd_sc_hd__buf_12_315/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_132 sky130_fd_sc_hd__xor2_1_234/X sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xor2_1_21/X sky130_fd_sc_hd__o21ai_1_44/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_284 sky130_fd_sc_hd__buf_12_284/A sky130_fd_sc_hd__buf_12_653/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_143 sky130_fd_sc_hd__xnor2_1_82/Y sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xnor2_1_19/Y sky130_fd_sc_hd__o21ai_1_65/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_295 sky130_fd_sc_hd__buf_12_295/A sky130_fd_sc_hd__buf_12_542/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_154 sky130_fd_sc_hd__xnor2_1_95/Y sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xnor2_1_32/Y sky130_fd_sc_hd__o21ai_1_88/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_165 sky130_fd_sc_hd__xnor2_1_104/Y sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xnor2_1_41/Y sky130_fd_sc_hd__a22oi_1_165/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_176 sky130_fd_sc_hd__nand2_1_133/A sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xor2_1_191/X sky130_fd_sc_hd__a22oi_1_176/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_187 sky130_fd_sc_hd__xor2_1_419/X sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xor2_1_207/X sky130_fd_sc_hd__a22oi_1_187/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_198 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__and2b_4_3/X sky130_fd_sc_hd__nor2_2_9/Y sky130_fd_sc_hd__a22oi_1_198/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_440 sky130_fd_sc_hd__nand2_1_368/B sky130_fd_sc_hd__nor2_1_118/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_451 sky130_fd_sc_hd__o21ai_1_505/A2 sky130_fd_sc_hd__xnor2_1_87/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_462 sky130_fd_sc_hd__a21oi_2_11/B1 sky130_fd_sc_hd__nand2_1_404/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_473 sky130_fd_sc_hd__a21oi_1_89/A1 sky130_fd_sc_hd__a21oi_1_92/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_484 sky130_fd_sc_hd__o21ai_1_591/B1 sky130_fd_sc_hd__nand2_1_443/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_495 sky130_fd_sc_hd__nand2_1_460/A sky130_fd_sc_hd__nor2_1_155/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_409 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_442/A2 sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_409/B1 sky130_fd_sc_hd__xor2_1_220/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2_4_18 sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__nor2_4_18/A
+ sky130_fd_sc_hd__nor2_4_18/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__nand2_2_11 sky130_fd_sc_hd__inv_4_7/A sky130_fd_sc_hd__nand2_2_11/A
+ sky130_fd_sc_hd__ha_2_9/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__decap_12_480 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_491 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_203 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__fa_2_140/B
+ sky130_fd_sc_hd__xor2_1_203/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_214 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__xor3_1_13/C
+ sky130_fd_sc_hd__xor2_1_214/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_225 sky130_fd_sc_hd__fa_2_198/A sky130_fd_sc_hd__fa_2_149/B
+ sky130_fd_sc_hd__xor2_1_225/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_236 sky130_fd_sc_hd__fa_2_170/A sky130_fd_sc_hd__xor2_1_236/X
+ sky130_fd_sc_hd__xor2_1_236/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_247 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__fa_2_162/A
+ sky130_fd_sc_hd__xor2_1_247/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_258 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__fa_2_169/A
+ sky130_fd_sc_hd__xor2_1_258/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_269 sky130_fd_sc_hd__xor2_1_383/B sky130_fd_sc_hd__fa_2_180/A
+ sky130_fd_sc_hd__xor2_1_269/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_207 vssd1 vccd1 sky130_fd_sc_hd__buf_8_31/A sky130_fd_sc_hd__buf_8_34/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_218 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_218/X sky130_fd_sc_hd__clkinv_1_884/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o21ai_1_910 vssd1 vccd1 sky130_fd_sc_hd__nor2_2_1/B sky130_fd_sc_hd__o21ai_1_912/B1
+ sky130_fd_sc_hd__and2_0_401/B sky130_fd_sc_hd__o21ai_1_910/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1490 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_229 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_37/A1 sky130_fd_sc_hd__clkbuf_1_229/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o21ai_1_921 vssd1 vccd1 sky130_fd_sc_hd__nand2_1_861/B la_data_out[52]
+ sky130_fd_sc_hd__a21oi_1_199/Y sky130_fd_sc_hd__nor4b_1_0/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_8_3 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__buf_2_30 vccd1 vssd1 sky130_fd_sc_hd__buf_2_30/X sky130_fd_sc_hd__buf_6_2/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_41 vccd1 vssd1 sky130_fd_sc_hd__buf_2_41/X sky130_fd_sc_hd__buf_2_41/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_52 vccd1 vssd1 sky130_fd_sc_hd__buf_2_53/A sky130_fd_sc_hd__buf_2_52/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_63 vccd1 vssd1 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__buf_2_63/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_74 vccd1 vssd1 sky130_fd_sc_hd__buf_2_74/X sky130_fd_sc_hd__buf_2_74/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_85 vccd1 vssd1 sky130_fd_sc_hd__buf_2_85/X sky130_fd_sc_hd__buf_2_85/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_96 vccd1 vssd1 sky130_fd_sc_hd__buf_2_96/X sky130_fd_sc_hd__buf_2_96/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__diode_2_3 sky130_fd_sc_hd__clkbuf_4_20/X vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__and2_0_205 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_51/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_78/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_216 vccd1 vssd1 sky130_fd_sc_hd__and2_0_216/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_216/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_227 vccd1 vssd1 sky130_fd_sc_hd__and2_0_227/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__o21ai_1_61/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_238 vccd1 vssd1 sky130_fd_sc_hd__and2_0_238/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_52/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_249 vccd1 vssd1 sky130_fd_sc_hd__and2_0_249/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_249/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__xor3_1_14 sky130_fd_sc_hd__xor3_1_14/X sky130_fd_sc_hd__xor3_1_14/C
+ sky130_fd_sc_hd__xor3_1_14/B sky130_fd_sc_hd__xor3_1_15/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__xor3_1_25 sky130_fd_sc_hd__xor3_1_25/X sky130_fd_sc_hd__xor3_1_25/C
+ sky130_fd_sc_hd__xor3_1_25/B sky130_fd_sc_hd__xor3_1_25/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__clkinv_1_270 sky130_fd_sc_hd__nand3_1_2/A sky130_fd_sc_hd__nor3_1_0/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_2_4 sky130_fd_sc_hd__nand2_1_7/B sky130_fd_sc_hd__fa_2_415/A
+ sky130_fd_sc_hd__or2_0_9/A sky130_fd_sc_hd__fa_2_415/B sky130_fd_sc_hd__nand2_1_8/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_2
Xsky130_fd_sc_hd__clkinv_1_281 sky130_fd_sc_hd__and2_0_106/A sky130_fd_sc_hd__a222oi_1_25/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_292 sky130_fd_sc_hd__and2_0_175/A sky130_fd_sc_hd__a222oi_1_36/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_0 sky130_fd_sc_hd__ha_2_9/B sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__a21oi_1_0/Y sky130_fd_sc_hd__nor2b_1_1/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkbuf_4_13 sky130_fd_sc_hd__buf_2_138/A sky130_fd_sc_hd__buf_2_139/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_206 vssd1 vccd1 sky130_fd_sc_hd__inv_2_14/Y sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__a222oi_1_80/Y sky130_fd_sc_hd__xor2_1_33/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_24 sky130_fd_sc_hd__inv_2_190/A sky130_fd_sc_hd__inv_2_189/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_217 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_251/A2 sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__a222oi_1_88/Y sky130_fd_sc_hd__xor2_1_43/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_35 sky130_fd_sc_hd__buf_6_74/A sky130_fd_sc_hd__buf_12_263/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_228 vssd1 vccd1 sky130_fd_sc_hd__inv_2_19/Y sky130_fd_sc_hd__nand2b_1_6/Y
+ sky130_fd_sc_hd__a222oi_1_96/Y sky130_fd_sc_hd__xor2_1_53/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_46 sky130_fd_sc_hd__buf_2_49/A sky130_fd_sc_hd__buf_6_93/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_239 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_59/Y sky130_fd_sc_hd__nor2_1_60/Y
+ sky130_fd_sc_hd__nand2_1_200/Y sky130_fd_sc_hd__o21ai_1_239/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__buf_8_130 sky130_fd_sc_hd__buf_8_130/A sky130_fd_sc_hd__buf_8_162/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_141 sky130_fd_sc_hd__inv_2_83/Y sky130_fd_sc_hd__buf_8_160/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nor2_4_3 sky130_fd_sc_hd__nor2_4_3/Y sky130_fd_sc_hd__nor2_4_3/A
+ sky130_fd_sc_hd__nor2_4_4/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__buf_8_152 sky130_fd_sc_hd__inv_2_187/Y sky130_fd_sc_hd__buf_8_152/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_163 sky130_fd_sc_hd__buf_6_20/X sky130_fd_sc_hd__buf_8_163/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_406 sky130_fd_sc_hd__dfxtp_1_406/Q sky130_fd_sc_hd__dfxtp_1_410/CLK
+ sky130_fd_sc_hd__nor2b_1_109/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_417 sky130_fd_sc_hd__dfxtp_1_417/Q sky130_fd_sc_hd__dfxtp_1_417/CLK
+ sky130_fd_sc_hd__nor2b_1_98/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_428 sky130_fd_sc_hd__dfxtp_1_428/Q sky130_fd_sc_hd__clkinv_4_9/Y
+ sky130_fd_sc_hd__nor2b_1_119/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_439 sky130_fd_sc_hd__dfxtp_1_439/Q sky130_fd_sc_hd__dfxtp_1_439/CLK
+ sky130_fd_sc_hd__nor2b_1_108/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a222oi_1_108 vccd1 vssd1 sky130_fd_sc_hd__and3_4_2/X sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__buf_4_3/X sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__o21ai_1_243/B1 sky130_fd_sc_hd__and2b_4_4/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__o21ai_1_740 vssd1 vccd1 sky130_fd_sc_hd__buf_2_13/X sky130_fd_sc_hd__nand2b_1_20/Y
+ sky130_fd_sc_hd__o21ai_1_740/B1 sky130_fd_sc_hd__xor2_1_516/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_119 vccd1 vssd1 sky130_fd_sc_hd__and3_4_1/X sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__nor2_2_10/B sky130_fd_sc_hd__nor2_2_9/Y sky130_fd_sc_hd__buf_6_4/X
+ sky130_fd_sc_hd__o21ai_1_257/B1 sky130_fd_sc_hd__and2b_4_3/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__o21ai_1_751 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_751/A2 sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_751/B1 sky130_fd_sc_hd__xor2_1_527/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_762 vssd1 vccd1 sky130_fd_sc_hd__inv_2_49/Y sky130_fd_sc_hd__nand2b_1_16/Y
+ sky130_fd_sc_hd__o21ai_1_762/B1 sky130_fd_sc_hd__xor2_1_537/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_773 vssd1 vccd1 sky130_fd_sc_hd__buf_2_12/X sky130_fd_sc_hd__nand2b_1_16/Y
+ sky130_fd_sc_hd__o21ai_1_773/B1 sky130_fd_sc_hd__xor2_1_547/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_6_0 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__o21ai_1_784 vssd1 vccd1 sky130_fd_sc_hd__inv_2_51/Y sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_784/B1 sky130_fd_sc_hd__xor2_1_558/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_795 vssd1 vccd1 sky130_fd_sc_hd__inv_2_47/Y sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_795/B1 sky130_fd_sc_hd__xor2_1_569/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkinv_8_16 sky130_fd_sc_hd__clkinv_8_16/Y sky130_fd_sc_hd__clkinv_8_17/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_27 sky130_fd_sc_hd__clkinv_8_27/Y sky130_fd_sc_hd__clkinv_8_28/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_38 sky130_fd_sc_hd__clkinv_8_38/Y sky130_fd_sc_hd__clkinv_8_38/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_49 sky130_fd_sc_hd__clkinv_8_76/A sky130_fd_sc_hd__clkinv_8_49/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_14 sky130_fd_sc_hd__buf_12_14/A sky130_fd_sc_hd__buf_12_14/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_25 sky130_fd_sc_hd__inv_2_136/Y sky130_fd_sc_hd__buf_12_25/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_80 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__xor2_1_80/X
+ sky130_fd_sc_hd__xor2_1_80/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_36 sky130_fd_sc_hd__buf_12_36/A sky130_fd_sc_hd__buf_12_36/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_91 sky130_fd_sc_hd__fa_2_97/A sky130_fd_sc_hd__fa_2_61/A
+ sky130_fd_sc_hd__xor2_1_91/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_47 sky130_fd_sc_hd__inv_2_174/Y sky130_fd_sc_hd__buf_12_47/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_58 sky130_fd_sc_hd__inv_2_184/Y sky130_fd_sc_hd__buf_12_58/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_69 sky130_fd_sc_hd__buf_8_28/X sky130_fd_sc_hd__buf_12_69/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_2_9 vccd1 vssd1 sky130_fd_sc_hd__buf_2_9/X sky130_fd_sc_hd__buf_2_9/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o21ai_2_12 sky130_fd_sc_hd__o21ai_2_12/B1 sky130_fd_sc_hd__o21ai_2_12/Y
+ sky130_fd_sc_hd__xor2_1_468/A sky130_fd_sc_hd__nor2_2_21/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__o21ai_2
Xsky130_fd_sc_hd__inv_2_9 sky130_fd_sc_hd__inv_2_9/A sky130_fd_sc_hd__inv_2_9/Y vccd1
+ vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__nor2_1_19 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_1_19/Y
+ sky130_fd_sc_hd__nor2_1_19/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__and2_0_30 vccd1 vssd1 sky130_fd_sc_hd__and2_0_30/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__buf_2_23/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_41 vccd1 vssd1 sky130_fd_sc_hd__and2_0_41/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__nor2_1_87/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_52 vccd1 vssd1 sky130_fd_sc_hd__and2_0_52/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__buf_6_5/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_63 vccd1 vssd1 sky130_fd_sc_hd__and2_0_63/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__or2_0_60/B vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_74 vccd1 vssd1 sky130_fd_sc_hd__and2_0_74/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__buf_4_2/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_407 sky130_fd_sc_hd__xor2_1_346/B sky130_fd_sc_hd__o21ai_2_9/B1
+ sky130_fd_sc_hd__nand2_1_407/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2_2_0 sky130_fd_sc_hd__nor2_2_0/B sky130_fd_sc_hd__nor2_2_0/Y
+ sky130_fd_sc_hd__nor2_4_0/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__and2_0_85 vccd1 vssd1 sky130_fd_sc_hd__and2_0_85/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__buf_4_3/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_418 sky130_fd_sc_hd__nand2_1_418/Y sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__buf_6_4/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_96 vccd1 vssd1 sky130_fd_sc_hd__and2_0_96/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__or2_0_39/B vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_429 sky130_fd_sc_hd__nand2_1_429/Y sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__nor2_2_10/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__buf_8_40 sky130_fd_sc_hd__buf_8_40/A sky130_fd_sc_hd__buf_8_40/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__clkinv_1_1009 sky130_fd_sc_hd__clkinv_1_1009/Y sky130_fd_sc_hd__clkinv_1_1009/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_51 sky130_fd_sc_hd__buf_8_51/A sky130_fd_sc_hd__buf_8_51/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_62 sky130_fd_sc_hd__buf_8_62/A sky130_fd_sc_hd__buf_8_62/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_73 sky130_fd_sc_hd__buf_8_73/A sky130_fd_sc_hd__buf_8_73/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_84 sky130_fd_sc_hd__buf_8_84/A sky130_fd_sc_hd__buf_8_84/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_203 sky130_fd_sc_hd__fa_2_389/A sky130_fd_sc_hd__dfxtp_2_0/CLK
+ sky130_fd_sc_hd__and2_0_50/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_8_95 sky130_fd_sc_hd__inv_4_13/Y sky130_fd_sc_hd__buf_8_95/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_214 sky130_fd_sc_hd__xor2_1_475/A sky130_fd_sc_hd__dfxtp_1_217/CLK
+ sky130_fd_sc_hd__and2_0_93/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_225 sky130_fd_sc_hd__xor2_1_396/A sky130_fd_sc_hd__dfxtp_2_4/CLK
+ sky130_fd_sc_hd__and2_0_52/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_236 sky130_fd_sc_hd__xnor2_1_90/A sky130_fd_sc_hd__dfxtp_2_5/CLK
+ sky130_fd_sc_hd__and2_0_76/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_247 sky130_fd_sc_hd__dfxtp_1_247/Q sky130_fd_sc_hd__clkinv_4_6/Y
+ sky130_fd_sc_hd__and2_0_10/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_258 sky130_fd_sc_hd__fa_2_122/A sky130_fd_sc_hd__dfxtp_1_266/CLK
+ sky130_fd_sc_hd__and2_0_40/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_269 sky130_fd_sc_hd__xor2_1_78/A sky130_fd_sc_hd__dfxtp_1_269/CLK
+ sky130_fd_sc_hd__and2_0_66/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_570 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_139/Y sky130_fd_sc_hd__nand2_1_431/Y
+ sky130_fd_sc_hd__nand2_1_426/Y sky130_fd_sc_hd__o21ai_1_570/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_581 vssd1 vccd1 sky130_fd_sc_hd__inv_2_28/Y sky130_fd_sc_hd__nand2b_2_3/Y
+ sky130_fd_sc_hd__o21ai_1_581/B1 sky130_fd_sc_hd__xor2_1_376/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_108 sky130_fd_sc_hd__nor2_2_3/A sky130_fd_sc_hd__or2_0_11/B
+ sky130_fd_sc_hd__fa_2_108/A sky130_fd_sc_hd__fa_2_108/B sky130_fd_sc_hd__fa_2_108/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o21ai_1_592 vssd1 vccd1 sky130_fd_sc_hd__buf_2_7/X sky130_fd_sc_hd__nand2b_2_3/Y
+ sky130_fd_sc_hd__o21ai_1_592/B1 sky130_fd_sc_hd__xor2_1_386/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_119 sky130_fd_sc_hd__nor2_1_80/A sky130_fd_sc_hd__nor2_1_83/B
+ sky130_fd_sc_hd__fa_2_119/A sky130_fd_sc_hd__fa_2_119/B sky130_fd_sc_hd__fa_2_119/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_103 vccd1 vssd1 sky130_fd_sc_hd__buf_2_103/X sky130_fd_sc_hd__buf_2_103/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_114 vccd1 vssd1 sky130_fd_sc_hd__buf_2_114/X sky130_fd_sc_hd__buf_2_114/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_125 vccd1 vssd1 sky130_fd_sc_hd__buf_2_125/X sky130_fd_sc_hd__buf_2_125/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_18 sky130_fd_sc_hd__o22ai_1_45/B1 sky130_fd_sc_hd__o22ai_1_18/B1
+ sky130_fd_sc_hd__o22ai_1_18/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__inv_4_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_136 vccd1 vssd1 sky130_fd_sc_hd__buf_2_136/X sky130_fd_sc_hd__buf_2_136/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_29 sky130_fd_sc_hd__o22ai_1_32/B1 sky130_fd_sc_hd__o21ai_1_2/A2
+ sky130_fd_sc_hd__o22ai_1_29/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__inv_4_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_147 vccd1 vssd1 sky130_fd_sc_hd__buf_2_147/X sky130_fd_sc_hd__buf_2_147/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_158 vccd1 vssd1 sky130_fd_sc_hd__buf_2_158/X sky130_fd_sc_hd__buf_2_188/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_169 vccd1 vssd1 la_data_out[53] sky130_fd_sc_hd__ha_2_35/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__ha_2_3 vssd1 vccd1 sky130_fd_sc_hd__ha_2_3/A sky130_fd_sc_hd__ha_2_10/B
+ sky130_fd_sc_hd__ha_2_3/SUM sky130_fd_sc_hd__ha_2_3/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__a222oi_1_450 vccd1 vssd1 sky130_fd_sc_hd__and3_4_25/X sky130_fd_sc_hd__buf_2_30/X
+ sky130_fd_sc_hd__buf_2_26/X sky130_fd_sc_hd__nor2_1_186/Y sky130_fd_sc_hd__buf_2_24/X
+ sky130_fd_sc_hd__o21ai_1_730/B1 sky130_fd_sc_hd__nor2b_1_17/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_461 vccd1 vssd1 sky130_fd_sc_hd__and3_4_26/X sky130_fd_sc_hd__buf_2_26/X
+ sky130_fd_sc_hd__buf_2_24/X sky130_fd_sc_hd__nor2_2_31/Y sky130_fd_sc_hd__buf_2_27/X
+ sky130_fd_sc_hd__o21ai_1_744/B1 sky130_fd_sc_hd__nor2b_1_12/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_472 vccd1 vssd1 sky130_fd_sc_hd__and3_4_18/X sky130_fd_sc_hd__buf_2_27/X
+ sky130_fd_sc_hd__buf_2_15/X sky130_fd_sc_hd__nor2_2_32/Y sky130_fd_sc_hd__buf_2_4/A
+ sky130_fd_sc_hd__o21ai_1_759/B1 sky130_fd_sc_hd__nor2b_2_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_14 vssd1 vccd1 sky130_fd_sc_hd__nand2_1_133/A sky130_fd_sc_hd__xor2_1_403/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_483 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__buf_4_3/X sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__o21ai_1_771/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_25 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_25/X sky130_fd_sc_hd__nor2_4_3/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_494 vccd1 vssd1 sky130_fd_sc_hd__and3_4_20/X sky130_fd_sc_hd__buf_2_24/X
+ sky130_fd_sc_hd__buf_2_27/X sky130_fd_sc_hd__nor2_4_16/Y sky130_fd_sc_hd__buf_2_15/X
+ sky130_fd_sc_hd__o21ai_1_787/B1 sky130_fd_sc_hd__and2b_4_11/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_36 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_36/X sky130_fd_sc_hd__clkbuf_1_36/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_47 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_47/X sky130_fd_sc_hd__buf_8_26/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_58 vssd1 vccd1 sky130_fd_sc_hd__buf_2_61/A sky130_fd_sc_hd__clkbuf_1_60/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_69 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_13/A1 sky130_fd_sc_hd__clkbuf_1_69/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__or2_0_16 sky130_fd_sc_hd__or2_0_16/A sky130_fd_sc_hd__or2_0_16/X
+ sky130_fd_sc_hd__or2_0_16/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_27 sky130_fd_sc_hd__or2_0_27/A sky130_fd_sc_hd__or2_0_27/X
+ sky130_fd_sc_hd__or2_0_27/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_38 sky130_fd_sc_hd__or2_0_58/A sky130_fd_sc_hd__or2_0_38/X
+ sky130_fd_sc_hd__or2_0_9/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_49 sky130_fd_sc_hd__or2_0_49/A sky130_fd_sc_hd__or2_0_49/X
+ sky130_fd_sc_hd__or2_0_49/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__buf_12_3 sky130_fd_sc_hd__buf_12_3/A sky130_fd_sc_hd__buf_12_3/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_603 sky130_fd_sc_hd__buf_12_603/A sky130_fd_sc_hd__buf_12_603/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_614 sky130_fd_sc_hd__buf_12_614/A sky130_fd_sc_hd__buf_12_614/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_625 sky130_fd_sc_hd__buf_12_625/A sky130_fd_sc_hd__buf_12_625/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_636 sky130_fd_sc_hd__buf_12_636/A sky130_fd_sc_hd__buf_12_636/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_4_107 sky130_fd_sc_hd__clkinv_2_60/Y sky130_fd_sc_hd__dfxtp_1_20/CLK
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_12_647 sky130_fd_sc_hd__buf_12_647/A sky130_fd_sc_hd__buf_12_647/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_4_118 sky130_fd_sc_hd__clkinv_8_73/Y sky130_fd_sc_hd__clkinv_4_119/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_12_658 sky130_fd_sc_hd__buf_12_658/A sky130_fd_sc_hd__buf_12_658/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_669 sky130_fd_sc_hd__buf_12_669/A sky130_fd_sc_hd__buf_12_669/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_309 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_204 sky130_fd_sc_hd__xnor2_1_20/A sky130_fd_sc_hd__nand2_1_205/Y
+ sky130_fd_sc_hd__or2_0_14/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_803 sky130_fd_sc_hd__and2_0_304/A sky130_fd_sc_hd__clkinv_1_803/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_215 sky130_fd_sc_hd__xnor2_1_24/A sky130_fd_sc_hd__nand2_1_216/Y
+ sky130_fd_sc_hd__or2_0_20/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_814 sky130_fd_sc_hd__clkinv_1_814/Y sky130_fd_sc_hd__nand2_1_807/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_226 sky130_fd_sc_hd__nand2_1_226/Y sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__buf_4_4/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_825 sky130_fd_sc_hd__nand2_1_828/A sky130_fd_sc_hd__nor2_1_263/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_237 sky130_fd_sc_hd__nand2_1_237/Y sky130_fd_sc_hd__nor2_2_3/A
+ sky130_fd_sc_hd__nor2_2_3/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_836 sky130_fd_sc_hd__inv_2_73/A sky130_fd_sc_hd__ha_2_36/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_248 sky130_fd_sc_hd__xor2_1_146/B sky130_fd_sc_hd__nand2_1_249/Y
+ sky130_fd_sc_hd__nand2_1_248/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_847 sky130_fd_sc_hd__clkinv_1_847/Y sky130_fd_sc_hd__clkinv_4_13/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_259 sky130_fd_sc_hd__xnor2_1_41/A sky130_fd_sc_hd__nand2_1_260/Y
+ sky130_fd_sc_hd__nand2_1_259/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_858 sky130_fd_sc_hd__clkinv_1_858/Y sky130_fd_sc_hd__inv_2_195/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_869 sky130_fd_sc_hd__clkinv_1_869/Y sky130_fd_sc_hd__clkinv_4_83/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__conb_1_14 sky130_fd_sc_hd__conb_1_14/LO sky130_fd_sc_hd__conb_1_14/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_25 sky130_fd_sc_hd__conb_1_25/LO sky130_fd_sc_hd__conb_1_25/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_36 sky130_fd_sc_hd__conb_1_36/LO sky130_fd_sc_hd__conb_1_36/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1308 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_47 sky130_fd_sc_hd__conb_1_47/LO sky130_fd_sc_hd__conb_1_47/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1319 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_58 sky130_fd_sc_hd__conb_1_58/LO sky130_fd_sc_hd__conb_1_58/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_69 sky130_fd_sc_hd__conb_1_69/LO sky130_fd_sc_hd__conb_1_69/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__mux2_2_9 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_9/A1 sky130_fd_sc_hd__buf_2_73/X
+ sky130_fd_sc_hd__mux2_8_0/S sky130_fd_sc_hd__mux2_2_9/X vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__decap_12_810 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_821 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_832 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_843 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_854 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_865 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_876 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_760 sky130_fd_sc_hd__xor2_1_662/B sky130_fd_sc_hd__nand2_1_776/Y
+ sky130_fd_sc_hd__nand2_1_760/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_887 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_771 sky130_fd_sc_hd__nand2_1_771/Y sky130_fd_sc_hd__or2_1_12/A
+ sky130_fd_sc_hd__or2_1_12/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_898 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_782 sky130_fd_sc_hd__nand2_1_782/Y sky130_fd_sc_hd__nor2_1_249/A
+ sky130_fd_sc_hd__nor2_1_249/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_793 sky130_fd_sc_hd__nand2_1_793/Y sky130_fd_sc_hd__nor2_1_254/A
+ sky130_fd_sc_hd__nor2_1_254/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_1820 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1831 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1842 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1853 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1864 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_280 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__or2_0_60/B sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__or2_0_60/A
+ sky130_fd_sc_hd__o21ai_1_486/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_291 vccd1 vssd1 sky130_fd_sc_hd__and3_4_10/X sky130_fd_sc_hd__and2_0_38/A
+ sky130_fd_sc_hd__and2_0_49/A sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__and2_0_45/A
+ sky130_fd_sc_hd__o21ai_1_501/B1 sky130_fd_sc_hd__and2b_4_7/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_450 sky130_fd_sc_hd__fa_2_459/CIN sky130_fd_sc_hd__fa_2_450/SUM
+ sky130_fd_sc_hd__fa_2_450/A sky130_fd_sc_hd__fa_2_450/B sky130_fd_sc_hd__fa_2_450/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_461 sky130_fd_sc_hd__xor2_1_675/A sky130_fd_sc_hd__fa_2_460/A
+ sky130_fd_sc_hd__fa_2_461/A sky130_fd_sc_hd__fa_2_461/B sky130_fd_sc_hd__nor2b_1_27/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_472 sky130_fd_sc_hd__nor2_1_255/B sky130_fd_sc_hd__or2_0_101/A
+ sky130_fd_sc_hd__fa_2_472/A sky130_fd_sc_hd__fa_2_472/B sky130_fd_sc_hd__nor2b_1_43/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_483 sky130_fd_sc_hd__or2_0_106/B sky130_fd_sc_hd__nor2_1_261/A
+ sky130_fd_sc_hd__fa_2_483/A sky130_fd_sc_hd__fa_2_483/B sky130_fd_sc_hd__nor2b_1_65/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__decap_8_11 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__nor2_1_204 sky130_fd_sc_hd__buf_2_4/A sky130_fd_sc_hd__nor2_1_204/Y
+ sky130_fd_sc_hd__buf_2_20/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_215 sky130_fd_sc_hd__nor2_1_218/Y sky130_fd_sc_hd__nor2_1_215/Y
+ sky130_fd_sc_hd__nor2_1_217/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_226 sky130_fd_sc_hd__mux2_2_47/X sky130_fd_sc_hd__nor2_1_226/Y
+ sky130_fd_sc_hd__mux2_2_27/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_237 sky130_fd_sc_hd__nor2_1_237/B sky130_fd_sc_hd__nor2_1_237/Y
+ sky130_fd_sc_hd__nor2_1_237/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_248 sky130_fd_sc_hd__ha_2_14/SUM sky130_fd_sc_hd__nor2_1_248/Y
+ sky130_fd_sc_hd__o22ai_1_86/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_259 sky130_fd_sc_hd__nor2_1_259/B sky130_fd_sc_hd__nor2_1_259/Y
+ sky130_fd_sc_hd__nor2_1_259/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_400 sky130_fd_sc_hd__buf_12_400/A sky130_fd_sc_hd__buf_12_655/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_411 sky130_fd_sc_hd__buf_12_411/A sky130_fd_sc_hd__buf_12_584/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_422 sky130_fd_sc_hd__buf_12_422/A sky130_fd_sc_hd__buf_12_594/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_433 sky130_fd_sc_hd__buf_12_433/A sky130_fd_sc_hd__buf_12_614/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_444 sky130_fd_sc_hd__buf_12_444/A sky130_fd_sc_hd__buf_12_444/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_455 sky130_fd_sc_hd__buf_12_455/A sky130_fd_sc_hd__buf_12_561/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_466 sky130_fd_sc_hd__buf_12_466/A sky130_fd_sc_hd__buf_12_466/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_477 sky130_fd_sc_hd__buf_12_477/A sky130_fd_sc_hd__buf_12_477/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_106 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_488 sky130_fd_sc_hd__buf_12_488/A sky130_fd_sc_hd__buf_12_593/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_117 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_499 sky130_fd_sc_hd__buf_12_499/A sky130_fd_sc_hd__buf_12_589/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_128 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_600 sky130_fd_sc_hd__nand2_1_631/A sky130_fd_sc_hd__nor2_1_211/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_139 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_611 sky130_fd_sc_hd__clkinv_1_611/Y sky130_fd_sc_hd__nand2_1_661/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_622 sky130_fd_sc_hd__buf_2_28/A sky130_fd_sc_hd__inv_4_8/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_633 sky130_fd_sc_hd__clkinv_1_633/Y sky130_fd_sc_hd__nand2_1_679/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_644 sky130_fd_sc_hd__nand2_1_700/A sky130_fd_sc_hd__nor2_1_230/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_207 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_207/B sky130_fd_sc_hd__a22o_1_17/B1
+ sky130_fd_sc_hd__xnor2_1_207/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_655 sky130_fd_sc_hd__o22ai_1_78/B1 la_data_out[85] vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_218 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_218/B sky130_fd_sc_hd__a22o_1_8/A2
+ sky130_fd_sc_hd__xnor2_1_218/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_666 sky130_fd_sc_hd__nand2_1_734/A sky130_fd_sc_hd__nor2_1_238/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_229 vssd1 vccd1 sky130_fd_sc_hd__buf_2_207/X sky130_fd_sc_hd__xnor2_1_229/Y
+ sky130_fd_sc_hd__or2_0_82/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_677 sky130_fd_sc_hd__nand2_1_751/A sky130_fd_sc_hd__nor2_1_241/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_688 sky130_fd_sc_hd__nand2_1_763/A sky130_fd_sc_hd__nor2_1_251/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_699 sky130_fd_sc_hd__nand2_1_755/A sky130_fd_sc_hd__nor2_1_253/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1105 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1116 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1127 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1138 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1149 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_20 vccd1 vssd1 sky130_fd_sc_hd__xor2_1_411/X sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__xor2_1_624/X sky130_fd_sc_hd__xor2_1_199/X sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_20/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_31 vccd1 vssd1 sky130_fd_sc_hd__xnor2_1_95/Y sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__xnor2_1_158/Y sky130_fd_sc_hd__xnor2_1_32/Y sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_31/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_42 vccd1 vssd1 sky130_fd_sc_hd__xor2_1_276/X sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__inv_2_60/A sky130_fd_sc_hd__xor2_1_63/X sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_42/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_53 vccd1 vssd1 sky130_fd_sc_hd__and3_4_5/X sky130_fd_sc_hd__nor2_2_4/B
+ sky130_fd_sc_hd__buf_2_4/X sky130_fd_sc_hd__nor2_1_68/Y sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__a222oi_1_53/Y sky130_fd_sc_hd__nor2b_1_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_640 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_64 vccd1 vssd1 sky130_fd_sc_hd__and3_4_8/X sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__nor2_1_73/B sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__a222oi_1_64/Y sky130_fd_sc_hd__nor2b_2_2/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_651 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_11 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_11/B sky130_fd_sc_hd__xnor2_1_11/Y
+ sky130_fd_sc_hd__xnor2_1_11/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__a222oi_1_75 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__or2_0_58/B
+ sky130_fd_sc_hd__or2_0_58/A sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__or2_0_9/B
+ sky130_fd_sc_hd__a222oi_1_75/Y sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_662 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_22 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_22/B sky130_fd_sc_hd__xnor2_1_22/Y
+ sky130_fd_sc_hd__xnor2_1_22/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__a222oi_1_86 vccd1 vssd1 sky130_fd_sc_hd__and3_4_7/X sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__nor2_1_87/A sky130_fd_sc_hd__nor2_2_7/Y sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__a222oi_1_86/Y sky130_fd_sc_hd__nor2b_2_1/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__xnor2_1_33 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_33/B sky130_fd_sc_hd__inv_2_24/A
+ sky130_fd_sc_hd__xnor2_1_33/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_673 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_97 vccd1 vssd1 sky130_fd_sc_hd__and3_4_1/X sky130_fd_sc_hd__buf_6_4/X
+ sky130_fd_sc_hd__buf_6_0/X sky130_fd_sc_hd__nor2_2_9/Y sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__a222oi_1_97/Y sky130_fd_sc_hd__and2b_4_3/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_684 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_44 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_44/B sky130_fd_sc_hd__xnor2_1_44/Y
+ sky130_fd_sc_hd__xnor2_1_44/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_695 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_55 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__nor2_4_9/A
+ sky130_fd_sc_hd__xnor2_1_55/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_66 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_66/B sky130_fd_sc_hd__buf_2_10/A
+ sky130_fd_sc_hd__xnor2_1_66/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_407 sky130_fd_sc_hd__fa_2_281/A sky130_fd_sc_hd__fa_2_278/B
+ sky130_fd_sc_hd__xor2_1_407/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_590 sky130_fd_sc_hd__nand2_1_590/Y sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__buf_6_4/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_77 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_77/B sky130_fd_sc_hd__and3_1_1/C
+ sky130_fd_sc_hd__fa_2_198/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_418 sky130_fd_sc_hd__dfxtp_2_5/Q sky130_fd_sc_hd__nor2_4_14/B
+ sky130_fd_sc_hd__xor2_1_418/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_88 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_317/A sky130_fd_sc_hd__and3_4_14/B
+ sky130_fd_sc_hd__xnor2_1_90/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_429 sky130_fd_sc_hd__fa_2_310/A sky130_fd_sc_hd__xor3_1_24/B
+ sky130_fd_sc_hd__xor2_1_429/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_99 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_362/A sky130_fd_sc_hd__nor2b_2_3/A
+ sky130_fd_sc_hd__xnor2_1_99/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_2_0 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_0/Y sky130_fd_sc_hd__xnor2_2_0/A
+ sky130_fd_sc_hd__xnor2_2_0/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_2
Xsky130_fd_sc_hd__decap_12_1650 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1661 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1672 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1683 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1694 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_3 sky130_fd_sc_hd__buf_12_674/A sky130_fd_sc_hd__buf_12_137/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__fa_2_280 sky130_fd_sc_hd__fa_2_279/B sky130_fd_sc_hd__or2_0_50/A
+ sky130_fd_sc_hd__fa_2_280/A sky130_fd_sc_hd__fa_2_280/B sky130_fd_sc_hd__fa_2_280/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_291 sky130_fd_sc_hd__fa_2_290/B sky130_fd_sc_hd__fa_2_292/CIN
+ sky130_fd_sc_hd__fa_2_291/A sky130_fd_sc_hd__fa_2_291/B sky130_fd_sc_hd__xor2_1_448/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor4_1_3 wbs_adr_i[15] wbs_adr_i[14] sky130_fd_sc_hd__nor4_1_3/Y
+ wbs_adr_i[12] wbs_adr_i[16] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor4_1
Xsky130_fd_sc_hd__a22oi_1_2 sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__a22oi_1_2/B2 sky130_fd_sc_hd__a22oi_1_2/A2 sky130_fd_sc_hd__a22oi_1_2/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__decap_12_7 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_2_18 sky130_fd_sc_hd__clkinv_2_18/Y sky130_fd_sc_hd__inv_2_105/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_29 sky130_fd_sc_hd__clkinv_2_29/Y sky130_fd_sc_hd__clkinv_2_29/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__buf_12_230 sky130_fd_sc_hd__buf_6_52/X sky130_fd_sc_hd__buf_12_452/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_241 sky130_fd_sc_hd__buf_6_77/X sky130_fd_sc_hd__buf_12_317/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_100 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_185/Q sky130_fd_sc_hd__dfxtp_1_153/Q sky130_fd_sc_hd__o21ai_1_6/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_252 sky130_fd_sc_hd__buf_8_163/X sky130_fd_sc_hd__buf_12_362/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_111 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_175/Q sky130_fd_sc_hd__dfxtp_1_143/Q sky130_fd_sc_hd__o21ai_1_17/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_263 sky130_fd_sc_hd__buf_12_263/A sky130_fd_sc_hd__buf_12_356/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_122 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_164/Q sky130_fd_sc_hd__dfxtp_1_132/Q sky130_fd_sc_hd__o21ai_1_28/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_274 sky130_fd_sc_hd__buf_12_6/X sky130_fd_sc_hd__buf_12_670/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_133 sky130_fd_sc_hd__xor2_1_234/X sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xor2_1_21/X sky130_fd_sc_hd__o21ai_1_45/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_285 sky130_fd_sc_hd__buf_12_5/X sky130_fd_sc_hd__buf_12_603/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_144 sky130_fd_sc_hd__xor2_1_296/X sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xor2_1_83/X sky130_fd_sc_hd__o21ai_1_68/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_296 sky130_fd_sc_hd__buf_12_296/A sky130_fd_sc_hd__buf_12_462/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_155 sky130_fd_sc_hd__xnor2_1_95/Y sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xnor2_1_32/Y sky130_fd_sc_hd__o21ai_1_89/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_166 sky130_fd_sc_hd__nand2_1_123/A sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xnor2_1_44/Y sky130_fd_sc_hd__a22oi_1_166/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_177 sky130_fd_sc_hd__nand2_1_133/A sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xor2_1_191/X sky130_fd_sc_hd__a22oi_1_177/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_188 sky130_fd_sc_hd__xor2_1_421/X sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xor2_1_209/X sky130_fd_sc_hd__a22oi_1_188/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_430 sky130_fd_sc_hd__o21ai_1_454/A2 sky130_fd_sc_hd__xnor2_1_76/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22oi_1_199 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__and2b_4_4/X sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__a22oi_1_199/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_441 sky130_fd_sc_hd__nand2_1_370/A sky130_fd_sc_hd__nor2_1_120/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_452 sky130_fd_sc_hd__nor2_1_122/A sky130_fd_sc_hd__nand2_1_392/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_463 sky130_fd_sc_hd__nand2_1_405/A sky130_fd_sc_hd__nor2_1_129/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_474 sky130_fd_sc_hd__nand2_1_427/A sky130_fd_sc_hd__nor2_1_132/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_485 sky130_fd_sc_hd__o21ai_1_591/A1 sky130_fd_sc_hd__nor2_1_105/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_496 sky130_fd_sc_hd__nand2_1_467/A sky130_fd_sc_hd__nor2_1_157/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_4_19 sky130_fd_sc_hd__nor2_4_19/Y sky130_fd_sc_hd__nor2_4_19/A
+ sky130_fd_sc_hd__nor2_4_19/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__nand2_2_12 sky130_fd_sc_hd__nand2_2_12/Y sky130_fd_sc_hd__or2_0_52/X
+ sky130_fd_sc_hd__xnor2_1_67/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__decap_12_470 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_481 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_492 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_204 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__or2_0_21/B
+ sky130_fd_sc_hd__xor2_1_204/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_215 sky130_fd_sc_hd__fa_2_198/A sky130_fd_sc_hd__xor3_1_14/C
+ sky130_fd_sc_hd__xor2_1_215/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_226 sky130_fd_sc_hd__fa_2_217/A sky130_fd_sc_hd__fa_2_149/A
+ sky130_fd_sc_hd__xor2_1_226/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_237 sky130_fd_sc_hd__fa_2_198/A sky130_fd_sc_hd__fa_2_151/A
+ sky130_fd_sc_hd__xor2_1_237/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_248 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__xor2_1_248/X
+ sky130_fd_sc_hd__xor2_1_248/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_259 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__xor2_1_259/X
+ sky130_fd_sc_hd__xor2_1_259/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_208 vssd1 vccd1 sky130_fd_sc_hd__buf_8_96/A sky130_fd_sc_hd__clkbuf_1_280/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o21ai_1_900 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_683/A sky130_fd_sc_hd__nor2_1_261/Y
+ sky130_fd_sc_hd__nand2_1_821/Y sky130_fd_sc_hd__xnor2_1_297/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1480 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_219 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_219/X sky130_fd_sc_hd__clkinv_1_864/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o21ai_1_911 vssd1 vccd1 sky130_fd_sc_hd__nand3_1_5/Y sky130_fd_sc_hd__nor2_1_275/Y
+ sky130_fd_sc_hd__a31oi_1_1/Y sky130_fd_sc_hd__o21ai_1_911/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1491 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_922 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_922/A2 la_data_out[56]
+ sky130_fd_sc_hd__a21oi_1_200/Y sky130_fd_sc_hd__nor4b_1_0/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_8_4 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__buf_2_20 vccd1 vssd1 sky130_fd_sc_hd__buf_2_20/X sky130_fd_sc_hd__buf_6_5/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_31 vccd1 vssd1 sky130_fd_sc_hd__buf_2_31/X sky130_fd_sc_hd__buf_2_31/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_42 vccd1 vssd1 sky130_fd_sc_hd__buf_2_42/X sky130_fd_sc_hd__buf_2_42/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_53 vccd1 vssd1 sky130_fd_sc_hd__buf_8_81/A sky130_fd_sc_hd__buf_2_53/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_64 vccd1 vssd1 sky130_fd_sc_hd__buf_2_66/A sky130_fd_sc_hd__buf_6_7/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_75 vccd1 vssd1 sky130_fd_sc_hd__buf_2_75/X sky130_fd_sc_hd__buf_2_75/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_86 vccd1 vssd1 sky130_fd_sc_hd__buf_2_86/X sky130_fd_sc_hd__buf_2_86/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_97 vccd1 vssd1 sky130_fd_sc_hd__buf_2_97/X sky130_fd_sc_hd__buf_2_97/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__diode_2_4 sky130_fd_sc_hd__clkbuf_4_20/X vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__and2_0_206 vccd1 vssd1 sky130_fd_sc_hd__and2_0_206/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_206/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_217 vccd1 vssd1 sky130_fd_sc_hd__and2_0_217/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__o21ai_1_69/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_228 vccd1 vssd1 sky130_fd_sc_hd__and2_0_228/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__o21ai_1_60/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_239 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_90/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_51/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__xor3_1_15 sky130_fd_sc_hd__xor3_1_15/X sky130_fd_sc_hd__xor3_1_15/C
+ sky130_fd_sc_hd__xor3_1_15/B sky130_fd_sc_hd__xor3_1_15/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__xor3_1_26 sky130_fd_sc_hd__xor3_1_26/X sky130_fd_sc_hd__xor3_1_27/X
+ sky130_fd_sc_hd__xor3_1_26/B sky130_fd_sc_hd__xor3_1_29/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__clkinv_1_260 sky130_fd_sc_hd__o21ai_1_129/A2 sky130_fd_sc_hd__xor2_1_612/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_271 sky130_fd_sc_hd__o21ai_1_160/A1 sky130_fd_sc_hd__xnor2_1_187/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_2_5 sky130_fd_sc_hd__nand2_1_7/B sky130_fd_sc_hd__mux2_4_5/X
+ sky130_fd_sc_hd__or2_0_4/B sky130_fd_sc_hd__mux2_2_0/X sky130_fd_sc_hd__nand2_1_8/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22o_2
Xsky130_fd_sc_hd__clkinv_1_282 sky130_fd_sc_hd__and2_0_105/A sky130_fd_sc_hd__a222oi_1_26/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_293 sky130_fd_sc_hd__and2_0_168/A sky130_fd_sc_hd__a222oi_1_37/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xor3_1_0 sky130_fd_sc_hd__xor3_1_0/X sky130_fd_sc_hd__xor3_1_1/X
+ sky130_fd_sc_hd__xor3_1_0/B sky130_fd_sc_hd__xor3_1_6/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__a21oi_1_1 sky130_fd_sc_hd__nor3_2_0/Y sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__a21oi_1_1/Y sky130_fd_sc_hd__nor2_4_3/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkbuf_4_14 sky130_fd_sc_hd__buf_2_137/A sky130_fd_sc_hd__clkbuf_4_18/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_207 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_207/A2 sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__a222oi_1_81/Y sky130_fd_sc_hd__xor2_1_34/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_25 sky130_fd_sc_hd__clkbuf_4_25/X sky130_fd_sc_hd__buf_12_66/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_218 vssd1 vccd1 sky130_fd_sc_hd__inv_2_10/Y sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__a222oi_1_89/Y sky130_fd_sc_hd__xor2_1_44/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_36 sky130_fd_sc_hd__buf_8_117/A sky130_fd_sc_hd__buf_12_256/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_229 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_0/Y sky130_fd_sc_hd__nand2b_2_0/Y
+ sky130_fd_sc_hd__a222oi_1_97/Y sky130_fd_sc_hd__xor2_1_54/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_47 sky130_fd_sc_hd__buf_2_50/A wbs_dat_i[1] vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__a21oi_1_190 sky130_fd_sc_hd__maj3_1_1/X sky130_fd_sc_hd__nor3_1_3/A
+ sky130_fd_sc_hd__a21oi_1_190/Y sky130_fd_sc_hd__ha_2_49/SUM vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_120 sky130_fd_sc_hd__buf_8_120/A sky130_fd_sc_hd__buf_6_42/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_131 sky130_fd_sc_hd__inv_2_89/Y sky130_fd_sc_hd__buf_8_131/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_142 sky130_fd_sc_hd__buf_8_142/A sky130_fd_sc_hd__buf_8_142/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nor2_4_4 sky130_fd_sc_hd__nor2_4_4/Y sky130_fd_sc_hd__ha_2_8/A sky130_fd_sc_hd__nor2_4_4/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__buf_8_153 sky130_fd_sc_hd__inv_2_186/Y sky130_fd_sc_hd__buf_8_153/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_164 sky130_fd_sc_hd__buf_6_23/X sky130_fd_sc_hd__buf_8_164/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_407 sky130_fd_sc_hd__dfxtp_1_407/Q sky130_fd_sc_hd__clkinv_4_8/Y
+ sky130_fd_sc_hd__nor2b_1_108/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_418 sky130_fd_sc_hd__dfxtp_1_418/Q sky130_fd_sc_hd__dfxtp_1_427/CLK
+ sky130_fd_sc_hd__nor2b_1_97/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_429 sky130_fd_sc_hd__dfxtp_1_429/Q sky130_fd_sc_hd__dfxtp_1_439/CLK
+ sky130_fd_sc_hd__nor2b_1_118/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_730 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_9/X sky130_fd_sc_hd__nand2b_1_21/Y
+ sky130_fd_sc_hd__o21ai_1_730/B1 sky130_fd_sc_hd__xor2_1_507/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_109 vccd1 vssd1 sky130_fd_sc_hd__and3_4_6/X sky130_fd_sc_hd__buf_4_1/X
+ sky130_fd_sc_hd__nor2_2_5/A sky130_fd_sc_hd__nor2_1_72/Y sky130_fd_sc_hd__nor2_2_5/B
+ sky130_fd_sc_hd__o21ai_1_244/B1 sky130_fd_sc_hd__nor2b_1_6/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__o21ai_1_741 vssd1 vccd1 sky130_fd_sc_hd__inv_2_48/Y sky130_fd_sc_hd__nand2b_1_21/Y
+ sky130_fd_sc_hd__o21ai_1_741/B1 sky130_fd_sc_hd__xor2_1_517/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_752 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_10/X sky130_fd_sc_hd__o21ai_1_752/A1
+ sky130_fd_sc_hd__o21ai_1_752/B1 sky130_fd_sc_hd__xnor2_1_152/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_763 vssd1 vccd1 sky130_fd_sc_hd__inv_2_43/Y sky130_fd_sc_hd__nand2b_2_6/Y
+ sky130_fd_sc_hd__o21ai_1_763/B1 sky130_fd_sc_hd__xor2_1_538/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_774 vssd1 vccd1 sky130_fd_sc_hd__inv_2_46/Y sky130_fd_sc_hd__nand2b_1_15/Y
+ sky130_fd_sc_hd__o21ai_1_774/B1 sky130_fd_sc_hd__xor2_1_548/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_6_1 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__o21ai_1_785 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_126/Y sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_785/B1 sky130_fd_sc_hd__xor2_1_560/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_796 vssd1 vccd1 sky130_fd_sc_hd__inv_2_44/Y sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__o21ai_1_796/B1 sky130_fd_sc_hd__xor2_1_570/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkinv_8_17 sky130_fd_sc_hd__clkinv_8_17/Y sky130_fd_sc_hd__clkinv_8_17/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_28 sky130_fd_sc_hd__clkinv_8_28/Y sky130_fd_sc_hd__clkinv_8_28/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_39 sky130_fd_sc_hd__clkinv_8_40/A sky130_fd_sc_hd__clkinv_8_39/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_15 sky130_fd_sc_hd__buf_12_15/A sky130_fd_sc_hd__buf_12_15/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_70 sky130_fd_sc_hd__xor2_1_9/B sky130_fd_sc_hd__fa_2_48/A
+ sky130_fd_sc_hd__xor2_1_70/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_26 sky130_fd_sc_hd__inv_2_132/Y sky130_fd_sc_hd__buf_12_26/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_81 sky130_fd_sc_hd__fa_2_97/A sky130_fd_sc_hd__fa_2_53/B
+ sky130_fd_sc_hd__xor2_1_81/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_37 sky130_fd_sc_hd__inv_2_169/A sky130_fd_sc_hd__buf_12_37/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_92 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__xor2_1_92/X
+ sky130_fd_sc_hd__xor2_1_92/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_48 sky130_fd_sc_hd__inv_2_181/Y sky130_fd_sc_hd__buf_12_48/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_59 sky130_fd_sc_hd__buf_12_59/A sky130_fd_sc_hd__buf_12_64/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__o21ai_2_13 sky130_fd_sc_hd__o21ai_2_13/B1 sky130_fd_sc_hd__o21ai_2_13/Y
+ sky130_fd_sc_hd__xor2_1_489/A sky130_fd_sc_hd__nor2_2_24/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__o21ai_2
Xsky130_fd_sc_hd__xor2_1_590 sky130_fd_sc_hd__fah_1_14/A sky130_fd_sc_hd__fah_1_13/B
+ sky130_fd_sc_hd__xor2_1_590/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__maj3_1_0 sky130_fd_sc_hd__maj3_1_0/C sky130_fd_sc_hd__maj3_1_0/X
+ sky130_fd_sc_hd__maj3_1_0/B la_data_out[46] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__and2_0_20 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_4_1/D sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__buf_2_32/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_31 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_2_5/D sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__buf_4_7/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_42 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_2_1/D sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__buf_2_21/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_53 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_2_4/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__buf_2_31/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_64 vccd1 vssd1 sky130_fd_sc_hd__and2_0_64/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__or2_0_60/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_75 vccd1 vssd1 sky130_fd_sc_hd__and2_0_75/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__buf_4_4/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_408 sky130_fd_sc_hd__o21ai_2_9/B1 sky130_fd_sc_hd__nor2_2_14/A
+ sky130_fd_sc_hd__nor2_2_14/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2_2_1 sky130_fd_sc_hd__nor2_2_1/B sky130_fd_sc_hd__nor2_2_1/Y
+ sky130_fd_sc_hd__nor2_2_1/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__and2_0_86 vccd1 vssd1 sky130_fd_sc_hd__and2_0_86/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__buf_6_0/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_419 sky130_fd_sc_hd__xor2_1_359/B sky130_fd_sc_hd__nand2_1_420/Y
+ sky130_fd_sc_hd__or2_1_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_97 vccd1 vssd1 sky130_fd_sc_hd__and2_0_97/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__or2_0_42/B vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_8_30 sky130_fd_sc_hd__buf_8_30/A sky130_fd_sc_hd__buf_8_30/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_41 sky130_fd_sc_hd__buf_8_41/A sky130_fd_sc_hd__buf_8_41/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_52 sky130_fd_sc_hd__buf_8_52/A sky130_fd_sc_hd__buf_8_52/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_63 sky130_fd_sc_hd__buf_8_63/A sky130_fd_sc_hd__buf_8_63/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_74 sky130_fd_sc_hd__inv_2_72/Y sky130_fd_sc_hd__buf_8_74/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_85 sky130_fd_sc_hd__ha_2_30/A sky130_fd_sc_hd__buf_8_85/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_204 sky130_fd_sc_hd__xnor2_1_160/A sky130_fd_sc_hd__dfxtp_2_2/CLK
+ sky130_fd_sc_hd__and2_0_71/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_8_96 sky130_fd_sc_hd__buf_8_96/A sky130_fd_sc_hd__buf_8_96/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_215 sky130_fd_sc_hd__fa_2_310/A sky130_fd_sc_hd__dfxtp_1_217/CLK
+ sky130_fd_sc_hd__and2_0_91/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_226 sky130_fd_sc_hd__buf_2_6/A sky130_fd_sc_hd__dfxtp_1_230/CLK
+ sky130_fd_sc_hd__and2_0_48/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_237 sky130_fd_sc_hd__xor2_1_317/A sky130_fd_sc_hd__dfxtp_2_5/CLK
+ sky130_fd_sc_hd__and2_0_62/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_248 sky130_fd_sc_hd__xor2_1_212/A sky130_fd_sc_hd__clkinv_4_6/Y
+ sky130_fd_sc_hd__and2_0_34/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_259 sky130_fd_sc_hd__xnor2_1_38/A sky130_fd_sc_hd__dfxtp_1_269/CLK
+ sky130_fd_sc_hd__and2_0_88/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_560 vssd1 vccd1 sky130_fd_sc_hd__inv_2_36/Y sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_560/B1 sky130_fd_sc_hd__xor2_1_358/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_571 vssd1 vccd1 sky130_fd_sc_hd__inv_2_34/Y sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_571/B1 sky130_fd_sc_hd__xor2_1_368/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_582 vssd1 vccd1 sky130_fd_sc_hd__nand2_2_12/Y sky130_fd_sc_hd__nand2b_1_9/Y
+ sky130_fd_sc_hd__a22oi_1_209/Y sky130_fd_sc_hd__xor2_1_377/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_109 sky130_fd_sc_hd__fa_2_106/CIN sky130_fd_sc_hd__fah_1_0/A
+ sky130_fd_sc_hd__fa_2_109/A sky130_fd_sc_hd__fa_2_109/B sky130_fd_sc_hd__xor2_1_151/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o21ai_1_593 vssd1 vccd1 sky130_fd_sc_hd__inv_2_29/Y sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_593/B1 sky130_fd_sc_hd__xor2_1_387/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__buf_2_104 vccd1 vssd1 sky130_fd_sc_hd__buf_2_104/X sky130_fd_sc_hd__buf_2_104/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_115 vccd1 vssd1 sky130_fd_sc_hd__buf_2_115/X sky130_fd_sc_hd__buf_2_115/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_126 vccd1 vssd1 sky130_fd_sc_hd__buf_2_126/X sky130_fd_sc_hd__buf_2_126/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_19 sky130_fd_sc_hd__o22ai_1_44/B1 sky130_fd_sc_hd__o22ai_1_19/B1
+ sky130_fd_sc_hd__o22ai_1_19/Y sky130_fd_sc_hd__nor2_4_2/B sky130_fd_sc_hd__inv_4_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_137 vccd1 vssd1 sky130_fd_sc_hd__buf_2_137/X sky130_fd_sc_hd__buf_2_137/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_148 vccd1 vssd1 sky130_fd_sc_hd__buf_2_148/X sky130_fd_sc_hd__buf_2_148/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_159 vccd1 vssd1 sky130_fd_sc_hd__buf_2_159/X sky130_fd_sc_hd__buf_2_159/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__ha_2_4 vssd1 vccd1 sky130_fd_sc_hd__ha_2_4/A sky130_fd_sc_hd__ha_2_3/B
+ sky130_fd_sc_hd__ha_2_4/SUM sky130_fd_sc_hd__ha_2_4/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__a222oi_1_440 vccd1 vssd1 sky130_fd_sc_hd__and3_4_24/X sky130_fd_sc_hd__or2_0_71/B
+ sky130_fd_sc_hd__buf_2_29/X sky130_fd_sc_hd__nor2_1_183/Y sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__o21ai_1_717/B1 sky130_fd_sc_hd__nor2b_1_16/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_451 vccd1 vssd1 sky130_fd_sc_hd__and3_4_26/X sky130_fd_sc_hd__buf_2_27/X
+ sky130_fd_sc_hd__buf_2_15/X sky130_fd_sc_hd__nor2_2_31/Y sky130_fd_sc_hd__buf_2_4/A
+ sky130_fd_sc_hd__o21ai_1_731/B1 sky130_fd_sc_hd__nor2b_1_12/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_462 vccd1 vssd1 sky130_fd_sc_hd__and3_4_25/X sky130_fd_sc_hd__or2_0_71/B
+ sky130_fd_sc_hd__buf_2_29/X sky130_fd_sc_hd__nor2_1_186/Y sky130_fd_sc_hd__buf_2_30/X
+ sky130_fd_sc_hd__o21ai_1_745/B1 sky130_fd_sc_hd__nor2b_1_17/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_473 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__nor2_1_73/B sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__o21ai_1_760/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_15 vssd1 vccd1 sky130_fd_sc_hd__nand2_1_131/A sky130_fd_sc_hd__xor2_1_399/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_484 vccd1 vssd1 sky130_fd_sc_hd__and3_4_18/X sky130_fd_sc_hd__buf_2_26/X
+ sky130_fd_sc_hd__buf_2_24/X sky130_fd_sc_hd__nor2_2_32/Y sky130_fd_sc_hd__buf_2_27/X
+ sky130_fd_sc_hd__o21ai_1_773/B1 sky130_fd_sc_hd__nor2b_2_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_26 vssd1 vccd1 sky130_fd_sc_hd__and2_0_25/A sky130_fd_sc_hd__buf_4_1/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_495 vccd1 vssd1 sky130_fd_sc_hd__and3_4_21/X sky130_fd_sc_hd__buf_2_4/A
+ sky130_fd_sc_hd__buf_2_20/X sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__buf_2_21/X
+ sky130_fd_sc_hd__o21ai_1_788/B1 sky130_fd_sc_hd__and2b_4_12/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_37 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_37/X sky130_fd_sc_hd__buf_2_37/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_48 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_56/A sky130_fd_sc_hd__clkbuf_1_49/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_59 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_59/X sky130_fd_sc_hd__clkbuf_1_60/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__or2_0_17 sky130_fd_sc_hd__buf_4_5/X sky130_fd_sc_hd__or2_0_17/X
+ sky130_fd_sc_hd__buf_4_4/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_28 sky130_fd_sc_hd__or2_0_28/A sky130_fd_sc_hd__or2_0_28/X
+ sky130_fd_sc_hd__or2_0_28/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_39 sky130_fd_sc_hd__or2_0_58/A sky130_fd_sc_hd__or2_0_39/X
+ sky130_fd_sc_hd__or2_0_39/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__buf_12_4 sky130_fd_sc_hd__buf_12_4/A sky130_fd_sc_hd__buf_12_4/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_604 sky130_fd_sc_hd__buf_12_604/A sky130_fd_sc_hd__buf_12_604/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_615 sky130_fd_sc_hd__buf_12_615/A sky130_fd_sc_hd__buf_12_615/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_626 sky130_fd_sc_hd__buf_12_626/A sky130_fd_sc_hd__buf_12_626/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_637 sky130_fd_sc_hd__buf_12_637/A sky130_fd_sc_hd__buf_12_637/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_4_108 sky130_fd_sc_hd__clkinv_8_69/A sky130_fd_sc_hd__clkinv_4_109/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_12_648 sky130_fd_sc_hd__buf_12_648/A sky130_fd_sc_hd__buf_12_648/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_4_119 sky130_fd_sc_hd__clkinv_4_119/A sky130_fd_sc_hd__clkinv_8_75/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_12_659 sky130_fd_sc_hd__buf_12_659/A sky130_fd_sc_hd__buf_12_659/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__o22ai_1_130 sky130_fd_sc_hd__nor2b_1_20/A sky130_fd_sc_hd__xnor2_1_278/Y
+ sky130_fd_sc_hd__fa_2_456/CIN sky130_fd_sc_hd__xnor2_1_285/Y sky130_fd_sc_hd__o22ai_1_78/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_205 sky130_fd_sc_hd__nand2_1_205/Y sky130_fd_sc_hd__or2_0_60/A
+ sky130_fd_sc_hd__or2_0_60/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_804 sky130_fd_sc_hd__and2_0_303/A sky130_fd_sc_hd__clkinv_1_804/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_216 sky130_fd_sc_hd__nand2_1_216/Y sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__buf_4_5/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_815 sky130_fd_sc_hd__nand2_1_808/A sky130_fd_sc_hd__nor2_1_258/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_227 sky130_fd_sc_hd__xor2_1_117/B sky130_fd_sc_hd__o21ai_2_8/B1
+ sky130_fd_sc_hd__nand2_1_227/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_826 sky130_fd_sc_hd__clkinv_1_826/Y sky130_fd_sc_hd__nand2_1_831/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_2_30 sky130_fd_sc_hd__nor2_2_30/B sky130_fd_sc_hd__nor2_2_30/Y
+ sky130_fd_sc_hd__nor2_2_30/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__nand2_1_238 sky130_fd_sc_hd__xnor2_1_0/B sky130_fd_sc_hd__nand2_1_239/Y
+ sky130_fd_sc_hd__nand2_1_238/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_837 sky130_fd_sc_hd__clkinv_1_839/A sky130_fd_sc_hd__buf_8_75/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_249 sky130_fd_sc_hd__nand2_1_249/Y sky130_fd_sc_hd__nor2_1_43/A
+ sky130_fd_sc_hd__nor2_1_43/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_848 sky130_fd_sc_hd__clkinv_1_848/Y sky130_fd_sc_hd__clkinv_4_13/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_859 sky130_fd_sc_hd__clkinv_1_859/Y sky130_fd_sc_hd__inv_2_195/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__conb_1_15 sky130_fd_sc_hd__conb_1_15/LO sky130_fd_sc_hd__conb_1_15/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_26 sky130_fd_sc_hd__conb_1_26/LO sky130_fd_sc_hd__conb_1_26/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_37 sky130_fd_sc_hd__conb_1_37/LO sky130_fd_sc_hd__conb_1_37/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1309 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__conb_1_48 sky130_fd_sc_hd__conb_1_48/LO sky130_fd_sc_hd__conb_1_48/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_59 sky130_fd_sc_hd__conb_1_59/LO sky130_fd_sc_hd__conb_1_59/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__o21ai_1_390 vssd1 vccd1 sky130_fd_sc_hd__inv_2_26/Y sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__nand2_1_162/Y sky130_fd_sc_hd__xor2_1_205/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_800 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_811 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_822 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_833 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_844 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_855 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_866 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_750 sky130_fd_sc_hd__nand2_1_750/Y sky130_fd_sc_hd__or2_0_92/A
+ sky130_fd_sc_hd__or2_0_92/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_877 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_761 sky130_fd_sc_hd__xor2_1_663/B sky130_fd_sc_hd__nand2_1_777/Y
+ sky130_fd_sc_hd__or2_0_94/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_888 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_772 sky130_fd_sc_hd__nand2_1_772/Y sky130_fd_sc_hd__nor2_1_243/A
+ sky130_fd_sc_hd__nor2_1_243/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_899 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_783 sky130_fd_sc_hd__nand2_1_783/Y sky130_fd_sc_hd__or2_0_96/A
+ sky130_fd_sc_hd__or2_0_96/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_794 sky130_fd_sc_hd__xnor2_1_291/A sky130_fd_sc_hd__nand2_1_795/Y
+ sky130_fd_sc_hd__or2_0_100/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_1810 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1821 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1832 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1843 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1854 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1865 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_270 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__or2_0_60/A
+ sky130_fd_sc_hd__or2_0_61/A sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__or2_0_42/B
+ sky130_fd_sc_hd__o21ai_1_472/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_281 vccd1 vssd1 sky130_fd_sc_hd__and3_4_11/X sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__nor2_1_73/B sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__o21ai_1_488/B1 sky130_fd_sc_hd__and2b_4_8/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_292 vccd1 vssd1 sky130_fd_sc_hd__and3_4_17/X sky130_fd_sc_hd__buf_2_19/X
+ sky130_fd_sc_hd__buf_6_5/X sky130_fd_sc_hd__nor2_2_20/Y sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__o21ai_1_502/B1 sky130_fd_sc_hd__nor2b_2_4/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_440 sky130_fd_sc_hd__fa_2_435/CIN sky130_fd_sc_hd__fa_2_438/A
+ sky130_fd_sc_hd__fa_2_440/A sky130_fd_sc_hd__fa_2_440/B sky130_fd_sc_hd__o22ai_1_82/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_451 sky130_fd_sc_hd__fa_2_451/COUT sky130_fd_sc_hd__fa_2_451/SUM
+ sky130_fd_sc_hd__fa_2_451/A sky130_fd_sc_hd__fa_2_451/B sky130_fd_sc_hd__fa_2_453/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_462 sky130_fd_sc_hd__fa_2_460/CIN sky130_fd_sc_hd__fa_2_462/SUM
+ sky130_fd_sc_hd__fa_2_462/A sky130_fd_sc_hd__fa_2_462/B sky130_fd_sc_hd__fa_2_462/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_473 sky130_fd_sc_hd__or2_0_101/B sky130_fd_sc_hd__nor2_1_256/A
+ sky130_fd_sc_hd__fa_2_473/A sky130_fd_sc_hd__fa_2_473/B sky130_fd_sc_hd__nor2b_1_45/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_484 sky130_fd_sc_hd__nor2_1_261/B sky130_fd_sc_hd__or2_0_107/A
+ sky130_fd_sc_hd__fa_2_484/A sky130_fd_sc_hd__fa_2_484/B sky130_fd_sc_hd__nor2b_1_67/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__decap_8_12 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__nor2_1_205 sky130_fd_sc_hd__nor2_1_206/Y sky130_fd_sc_hd__nor2_1_205/Y
+ sky130_fd_sc_hd__nor2_1_209/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_216 sky130_fd_sc_hd__buf_2_26/X sky130_fd_sc_hd__nor2_1_216/Y
+ sky130_fd_sc_hd__buf_2_30/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_227 sky130_fd_sc_hd__mux2_2_38/X sky130_fd_sc_hd__nor2_1_227/Y
+ sky130_fd_sc_hd__mux2_2_24/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_238 sky130_fd_sc_hd__xor2_1_662/X sky130_fd_sc_hd__nor2_1_238/Y
+ sky130_fd_sc_hd__nor2_1_238/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_249 sky130_fd_sc_hd__nor2_1_249/B sky130_fd_sc_hd__nor2_1_249/Y
+ sky130_fd_sc_hd__nor2_1_249/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_401 sky130_fd_sc_hd__buf_12_401/A sky130_fd_sc_hd__buf_12_401/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_412 sky130_fd_sc_hd__buf_12_412/A sky130_fd_sc_hd__buf_12_598/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_423 sky130_fd_sc_hd__buf_12_423/A sky130_fd_sc_hd__buf_12_571/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_434 sky130_fd_sc_hd__buf_12_434/A sky130_fd_sc_hd__buf_12_642/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_445 sky130_fd_sc_hd__buf_12_445/A sky130_fd_sc_hd__buf_12_504/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_456 sky130_fd_sc_hd__buf_12_456/A sky130_fd_sc_hd__buf_12_607/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_467 sky130_fd_sc_hd__buf_12_467/A sky130_fd_sc_hd__buf_12_543/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_478 sky130_fd_sc_hd__buf_12_478/A sky130_fd_sc_hd__buf_12_590/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_107 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_489 sky130_fd_sc_hd__buf_12_489/A sky130_fd_sc_hd__buf_12_633/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_118 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_129 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_601 sky130_fd_sc_hd__nand2_1_638/A sky130_fd_sc_hd__nor2_1_214/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_612 sky130_fd_sc_hd__nand2_1_658/A sky130_fd_sc_hd__o21a_1_5/A2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_623 sky130_fd_sc_hd__buf_2_14/A sky130_fd_sc_hd__inv_6_0/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_634 sky130_fd_sc_hd__nand2_1_680/A sky130_fd_sc_hd__nor2_1_225/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_645 sky130_fd_sc_hd__clkinv_1_645/Y sky130_fd_sc_hd__nand2_1_703/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_208 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_208/B sky130_fd_sc_hd__a22o_1_14/B1
+ sky130_fd_sc_hd__xnor2_1_208/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_656 sky130_fd_sc_hd__o22ai_1_112/B1 sky130_fd_sc_hd__or2_0_78/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_219 vssd1 vccd1 sky130_fd_sc_hd__or2_0_84/A sky130_fd_sc_hd__xnor2_1_219/Y
+ sky130_fd_sc_hd__or2_0_79/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_667 sky130_fd_sc_hd__xor2_1_654/A sky130_fd_sc_hd__o21ai_1_878/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_678 sky130_fd_sc_hd__xnor2_1_212/A sky130_fd_sc_hd__and2_0_301/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_689 sky130_fd_sc_hd__nand2_1_764/A sky130_fd_sc_hd__nor2_1_252/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1106 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1117 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1128 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1139 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_10 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_351/Q sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__o211ai_1_26/Y sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__a222oi_1_10/Y sky130_fd_sc_hd__dfxtp_1_302/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_21 vccd1 vssd1 sky130_fd_sc_hd__xnor2_1_120/Y sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__xnor2_1_182/Y sky130_fd_sc_hd__xnor2_1_57/Y sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_21/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_32 vccd1 vssd1 sky130_fd_sc_hd__xor2_1_346/X sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__xor2_1_559/X sky130_fd_sc_hd__xor2_1_133/X sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_32/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_43 vccd1 vssd1 sky130_fd_sc_hd__xnor2_1_82/Y sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__inv_2_55/A sky130_fd_sc_hd__xnor2_1_19/Y sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_43/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_630 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_54 vccd1 vssd1 sky130_fd_sc_hd__and3_4_7/X sky130_fd_sc_hd__nor2_2_10/B
+ sky130_fd_sc_hd__buf_6_4/X sky130_fd_sc_hd__nor2_2_7/Y sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__a222oi_1_54/Y sky130_fd_sc_hd__nor2b_2_1/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_641 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_65 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__or2_0_58/A
+ sky130_fd_sc_hd__or2_0_9/B sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__or2_0_9/A
+ sky130_fd_sc_hd__a222oi_1_65/Y sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__xnor2_1_12 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_14/B sky130_fd_sc_hd__and3_1_0/A
+ sky130_fd_sc_hd__xor2_1_49/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_652 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_76 vccd1 vssd1 sky130_fd_sc_hd__and3_4_8/X sky130_fd_sc_hd__buf_6_4/X
+ sky130_fd_sc_hd__buf_6_0/X sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__a222oi_1_76/Y sky130_fd_sc_hd__nor2b_2_2/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_663 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_87 vccd1 vssd1 sky130_fd_sc_hd__and3_4_6/X sky130_fd_sc_hd__nor2_2_4/B
+ sky130_fd_sc_hd__buf_2_4/X sky130_fd_sc_hd__nor2_1_72/Y sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__a222oi_1_87/Y sky130_fd_sc_hd__nor2b_1_6/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__xnor2_1_23 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_23/B sky130_fd_sc_hd__xnor2_1_23/Y
+ sky130_fd_sc_hd__xnor2_1_23/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_674 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_98 vccd1 vssd1 sky130_fd_sc_hd__and3_4_6/X sky130_fd_sc_hd__nor2_2_5/A
+ sky130_fd_sc_hd__nor2_2_5/B sky130_fd_sc_hd__nor2_1_72/Y sky130_fd_sc_hd__nor2_2_4/B
+ sky130_fd_sc_hd__a222oi_1_98/Y sky130_fd_sc_hd__nor2b_1_6/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__xnor2_1_34 vssd1 vccd1 sky130_fd_sc_hd__fa_2_110/A sky130_fd_sc_hd__and3_4_6/C
+ sky130_fd_sc_hd__xnor2_1_34/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_685 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_45 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_45/B sky130_fd_sc_hd__inv_2_20/A
+ sky130_fd_sc_hd__xnor2_1_45/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_696 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_56 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_56/B sky130_fd_sc_hd__inv_2_16/A
+ sky130_fd_sc_hd__xnor2_1_56/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_580 sky130_fd_sc_hd__o21ai_2_15/B1 sky130_fd_sc_hd__nor2_2_27/A
+ sky130_fd_sc_hd__nor2_2_27/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_67 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_67/B sky130_fd_sc_hd__buf_2_7/A
+ sky130_fd_sc_hd__xnor2_1_67/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_408 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__xor2_1_408/X
+ sky130_fd_sc_hd__xor2_1_408/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_591 sky130_fd_sc_hd__xor2_1_572/B sky130_fd_sc_hd__nand2_1_592/Y
+ sky130_fd_sc_hd__or2_1_1/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_78 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_78/B sky130_fd_sc_hd__xnor2_1_78/Y
+ sky130_fd_sc_hd__xnor2_1_78/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_419 sky130_fd_sc_hd__o21a_1_3/X sky130_fd_sc_hd__xor2_1_419/X
+ sky130_fd_sc_hd__xor2_1_419/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xnor2_1_89 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_89/B sky130_fd_sc_hd__inv_2_41/A
+ sky130_fd_sc_hd__xnor2_1_89/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_2_1 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_1/Y sky130_fd_sc_hd__xnor2_2_1/A
+ sky130_fd_sc_hd__xnor2_2_1/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_2
Xsky130_fd_sc_hd__decap_12_1640 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1651 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1662 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1673 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1684 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1695 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__fa_2_270 sky130_fd_sc_hd__fa_2_267/CIN sky130_fd_sc_hd__fa_2_271/A
+ sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__fa_2_270/B sky130_fd_sc_hd__xor2_1_395/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_281 sky130_fd_sc_hd__fa_2_280/CIN sky130_fd_sc_hd__or2_0_48/A
+ sky130_fd_sc_hd__fa_2_281/A sky130_fd_sc_hd__fa_2_281/B sky130_fd_sc_hd__xor2_1_417/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_292 sky130_fd_sc_hd__fa_2_283/B sky130_fd_sc_hd__fa_2_298/CIN
+ sky130_fd_sc_hd__fa_2_292/A sky130_fd_sc_hd__fa_2_292/B sky130_fd_sc_hd__fa_2_292/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor4_1_4 wbs_adr_i[23] wbs_adr_i[22] sky130_fd_sc_hd__nor4_1_4/Y
+ wbs_adr_i[20] wbs_adr_i[21] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor4_1
Xsky130_fd_sc_hd__a22oi_1_3 sky130_fd_sc_hd__nor2_4_0/Y sky130_fd_sc_hd__nor2_2_0/Y
+ sky130_fd_sc_hd__a22oi_1_3/B2 sky130_fd_sc_hd__nor2_1_235/A sky130_fd_sc_hd__a22oi_1_3/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__decap_12_8 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_2_19 sky130_fd_sc_hd__clkinv_2_19/Y sky130_fd_sc_hd__inv_2_200/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__buf_12_220 sky130_fd_sc_hd__buf_6_78/X sky130_fd_sc_hd__buf_12_220/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_231 sky130_fd_sc_hd__buf_6_47/X sky130_fd_sc_hd__buf_12_429/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_242 sky130_fd_sc_hd__buf_6_49/X sky130_fd_sc_hd__buf_12_380/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_101 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_184/Q sky130_fd_sc_hd__dfxtp_1_152/Q sky130_fd_sc_hd__o21ai_1_7/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_253 sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__buf_12_253/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_112 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_174/Q sky130_fd_sc_hd__dfxtp_1_142/Q sky130_fd_sc_hd__o21ai_1_18/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_264 sky130_fd_sc_hd__buf_12_264/A sky130_fd_sc_hd__buf_12_398/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_123 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_163/Q sky130_fd_sc_hd__dfxtp_1_131/Q sky130_fd_sc_hd__o21ai_1_29/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_275 sky130_fd_sc_hd__buf_12_275/A sky130_fd_sc_hd__buf_12_667/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_134 sky130_fd_sc_hd__xnor2_1_73/Y sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xnor2_1_10/Y sky130_fd_sc_hd__o21ai_1_48/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_286 sky130_fd_sc_hd__buf_12_286/A sky130_fd_sc_hd__buf_12_568/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_145 sky130_fd_sc_hd__xor2_1_296/X sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xor2_1_83/X sky130_fd_sc_hd__o21ai_1_69/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_297 sky130_fd_sc_hd__buf_12_297/A sky130_fd_sc_hd__buf_12_487/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_156 sky130_fd_sc_hd__xor2_1_346/X sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xor2_1_133/X sky130_fd_sc_hd__o21ai_1_92/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_167 sky130_fd_sc_hd__nand2_1_123/A sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xnor2_1_44/Y sky130_fd_sc_hd__a22oi_1_167/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_178 sky130_fd_sc_hd__nand2_1_135/A sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xnor2_1_54/Y sky130_fd_sc_hd__a22oi_1_178/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_420 sky130_fd_sc_hd__nand2_1_341/A sky130_fd_sc_hd__nor2_1_112/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22oi_1_189 sky130_fd_sc_hd__xor2_1_421/X sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xor2_1_209/X sky130_fd_sc_hd__a22oi_1_189/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_431 sky130_fd_sc_hd__nor2_1_114/B sky130_fd_sc_hd__nand2_1_365/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_442 sky130_fd_sc_hd__a21oi_2_9/B1 sky130_fd_sc_hd__nand2_1_373/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_453 sky130_fd_sc_hd__nand2_1_388/A sky130_fd_sc_hd__nor2_1_124/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_464 sky130_fd_sc_hd__nand2_1_407/A sky130_fd_sc_hd__nor2_2_14/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_475 sky130_fd_sc_hd__nand2_1_428/A sky130_fd_sc_hd__nor2_1_140/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_486 sky130_fd_sc_hd__nand2_1_444/A sky130_fd_sc_hd__nor2_1_148/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_497 sky130_fd_sc_hd__a21oi_1_98/B1 sky130_fd_sc_hd__nand2_1_474/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_2_13 sky130_fd_sc_hd__nand2_2_13/Y sky130_fd_sc_hd__or2_0_72/X
+ sky130_fd_sc_hd__nand2_2_13/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__nor4b_2_0 sky130_fd_sc_hd__a21o_2_4/B1 sky130_fd_sc_hd__nor4b_2_0/Y
+ sky130_fd_sc_hd__nor4b_2_0/C wbs_adr_i[10] sky130_fd_sc_hd__nor4b_2_0/B vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__nor4b_2
Xsky130_fd_sc_hd__decap_12_460 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_471 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_482 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_493 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_205 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__xor2_1_205/X
+ sky130_fd_sc_hd__xor2_1_205/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_216 sky130_fd_sc_hd__fa_2_170/A sky130_fd_sc_hd__xor3_1_14/B
+ sky130_fd_sc_hd__xor2_1_216/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_227 sky130_fd_sc_hd__dfxtp_2_5/Q sky130_fd_sc_hd__fa_2_150/A
+ sky130_fd_sc_hd__xor2_1_227/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_238 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__fa_2_152/B
+ sky130_fd_sc_hd__xor2_1_238/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_249 sky130_fd_sc_hd__fa_2_217/A sky130_fd_sc_hd__xor2_1_249/X
+ sky130_fd_sc_hd__xor2_1_249/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1470 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_209 vssd1 vccd1 sky130_fd_sc_hd__buf_12_16/A sky130_fd_sc_hd__clkbuf_1_50/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o21ai_1_901 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_684/A sky130_fd_sc_hd__nor2_1_262/Y
+ sky130_fd_sc_hd__nand2_1_825/Y sky130_fd_sc_hd__xnor2_1_298/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1481 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_912 vssd1 vccd1 sky130_fd_sc_hd__a221oi_1_3/B2 sky130_fd_sc_hd__nand3_1_5/B
+ sky130_fd_sc_hd__o21ai_1_912/B1 sky130_fd_sc_hd__a31oi_1_1/A3 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1492 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_923 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_923/A2 la_data_out[54]
+ sky130_fd_sc_hd__xnor2_1_311/Y sky130_fd_sc_hd__o21ai_1_923/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_8_5 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__buf_2_10 vccd1 vssd1 sky130_fd_sc_hd__buf_2_10/X sky130_fd_sc_hd__buf_2_10/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_21 vccd1 vssd1 sky130_fd_sc_hd__buf_2_21/X sky130_fd_sc_hd__buf_6_1/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_32 vccd1 vssd1 sky130_fd_sc_hd__buf_2_32/X sky130_fd_sc_hd__inv_6_0/Y
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_43 vccd1 vssd1 sky130_fd_sc_hd__buf_2_43/X sky130_fd_sc_hd__buf_2_43/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_54 vccd1 vssd1 sky130_fd_sc_hd__buf_2_54/X sky130_fd_sc_hd__inv_12_0/Y
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_65 vccd1 vssd1 sky130_fd_sc_hd__buf_2_65/X sky130_fd_sc_hd__buf_6_7/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_76 vccd1 vssd1 sky130_fd_sc_hd__buf_2_76/X sky130_fd_sc_hd__buf_2_76/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_87 vccd1 vssd1 sky130_fd_sc_hd__buf_2_87/X sky130_fd_sc_hd__buf_2_87/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_98 vccd1 vssd1 sky130_fd_sc_hd__buf_2_98/X sky130_fd_sc_hd__buf_2_98/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__diode_2_5 sky130_fd_sc_hd__clkinv_4_23/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__and2_0_207 vccd1 vssd1 sky130_fd_sc_hd__and2_0_207/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_77/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_218 vccd1 vssd1 sky130_fd_sc_hd__and2_0_218/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_68/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_229 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_56/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_59/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__xor3_1_16 sky130_fd_sc_hd__xor3_1_16/X sky130_fd_sc_hd__xor3_1_17/X
+ sky130_fd_sc_hd__xor3_1_16/B sky130_fd_sc_hd__xor3_1_19/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__xor3_1_27 sky130_fd_sc_hd__xor3_1_27/X sky130_fd_sc_hd__xor3_1_28/X
+ sky130_fd_sc_hd__xor3_1_27/B sky130_fd_sc_hd__xor3_1_27/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__clkinv_1_250 sky130_fd_sc_hd__o21ai_1_89/A2 sky130_fd_sc_hd__xnor2_1_158/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_261 sky130_fd_sc_hd__o21ai_1_133/A2 sky130_fd_sc_hd__xor2_1_616/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_272 sky130_fd_sc_hd__and2_0_151/A sky130_fd_sc_hd__a222oi_1_16/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_283 sky130_fd_sc_hd__and2_0_216/A sky130_fd_sc_hd__a222oi_1_27/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_294 sky130_fd_sc_hd__and2_0_161/A sky130_fd_sc_hd__a222oi_1_38/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xor3_1_1 sky130_fd_sc_hd__xor3_1_1/X sky130_fd_sc_hd__xor3_1_1/C
+ sky130_fd_sc_hd__xor3_1_2/X sky130_fd_sc_hd__xor3_1_1/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__a21oi_1_2 sky130_fd_sc_hd__nor2_4_3/Y sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__a21oi_1_2/Y sky130_fd_sc_hd__nor3_2_0/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkbuf_4_15 sky130_fd_sc_hd__buf_2_136/A sky130_fd_sc_hd__buf_12_1/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_208 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_2/X sky130_fd_sc_hd__nand2_1_181/Y
+ sky130_fd_sc_hd__a21oi_1_41/Y sky130_fd_sc_hd__xnor2_1_11/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_26 sky130_fd_sc_hd__clkbuf_4_26/X sky130_fd_sc_hd__buf_12_67/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_219 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_219/A2 sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__a222oi_1_90/Y sky130_fd_sc_hd__xor2_1_45/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_37 sky130_fd_sc_hd__buf_8_14/A sky130_fd_sc_hd__buf_12_264/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_48 sky130_fd_sc_hd__buf_2_51/A sky130_fd_sc_hd__buf_4_40/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__a21oi_1_180 sky130_fd_sc_hd__xnor2_1_301/B sky130_fd_sc_hd__clkinv_1_828/Y
+ sky130_fd_sc_hd__xor2_1_686/A sky130_fd_sc_hd__or2_0_110/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_191 la_data_out[43] sky130_fd_sc_hd__xor2_1_694/X sky130_fd_sc_hd__a21oi_1_191/Y
+ sky130_fd_sc_hd__nand2_1_859/B vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_110 sky130_fd_sc_hd__buf_6_23/A sky130_fd_sc_hd__buf_6_81/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_121 sky130_fd_sc_hd__buf_6_21/X sky130_fd_sc_hd__buf_8_121/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_132 sky130_fd_sc_hd__buf_8_132/A sky130_fd_sc_hd__buf_8_132/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_143 sky130_fd_sc_hd__buf_4_26/A sky130_fd_sc_hd__buf_6_25/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nor2_4_5 sky130_fd_sc_hd__nor2_4_5/Y sky130_fd_sc_hd__ha_2_8/A sky130_fd_sc_hd__nor2_4_5/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__buf_8_154 sky130_fd_sc_hd__inv_2_71/Y sky130_fd_sc_hd__buf_8_154/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_165 sky130_fd_sc_hd__buf_8_165/A sky130_fd_sc_hd__buf_8_165/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__decap_12_290 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_408 sky130_fd_sc_hd__dfxtp_1_408/Q sky130_fd_sc_hd__dfxtp_1_410/CLK
+ sky130_fd_sc_hd__nor2b_1_107/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_419 sky130_fd_sc_hd__dfxtp_1_419/Q sky130_fd_sc_hd__dfxtp_1_427/CLK
+ sky130_fd_sc_hd__nor2b_1_96/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_720 vssd1 vccd1 sky130_fd_sc_hd__inv_2_44/Y sky130_fd_sc_hd__nand2b_1_15/Y
+ sky130_fd_sc_hd__o21ai_1_720/B1 sky130_fd_sc_hd__xor2_1_497/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_731 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_3/Y sky130_fd_sc_hd__nand2b_1_15/Y
+ sky130_fd_sc_hd__o21ai_1_731/B1 sky130_fd_sc_hd__xor2_1_508/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_742 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_742/A2 sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_742/B1 sky130_fd_sc_hd__xor2_1_518/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_753 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_772/B1 sky130_fd_sc_hd__nor2_1_182/A
+ sky130_fd_sc_hd__nor2_1_181/Y sky130_fd_sc_hd__o21ai_1_753/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_764 vssd1 vccd1 sky130_fd_sc_hd__xor2_2_2/X sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__o21ai_1_764/B1 sky130_fd_sc_hd__xor2_1_539/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_775 vssd1 vccd1 sky130_fd_sc_hd__nand2_2_13/Y sky130_fd_sc_hd__nand2b_1_21/Y
+ sky130_fd_sc_hd__a22oi_1_217/Y sky130_fd_sc_hd__xor2_1_549/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_786 vssd1 vccd1 sky130_fd_sc_hd__a21oi_1_127/Y sky130_fd_sc_hd__nor2_1_188/A
+ sky130_fd_sc_hd__a21oi_1_119/Y sky130_fd_sc_hd__o21ai_1_786/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_797 vssd1 vccd1 sky130_fd_sc_hd__inv_2_50/Y sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_797/B1 sky130_fd_sc_hd__xor2_1_571/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkinv_8_18 sky130_fd_sc_hd__clkinv_8_18/Y sky130_fd_sc_hd__clkinv_8_18/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_29 sky130_fd_sc_hd__clkinv_8_30/A sky130_fd_sc_hd__clkinv_8_88/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__xor2_1_60 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__fa_2_40/A
+ sky130_fd_sc_hd__xor2_1_60/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_16 sky130_fd_sc_hd__buf_12_16/A sky130_fd_sc_hd__buf_12_16/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_71 sky130_fd_sc_hd__xor2_1_6/B sky130_fd_sc_hd__xor2_1_71/X
+ sky130_fd_sc_hd__xor2_1_71/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_27 sky130_fd_sc_hd__buf_12_27/A sky130_fd_sc_hd__buf_12_27/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_82 sky130_fd_sc_hd__xor2_1_6/B sky130_fd_sc_hd__fa_2_53/A
+ sky130_fd_sc_hd__xor2_1_82/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_38 sky130_fd_sc_hd__inv_2_177/Y sky130_fd_sc_hd__buf_12_38/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_93 sky130_fd_sc_hd__xor2_1_6/B sky130_fd_sc_hd__xor2_1_93/X
+ sky130_fd_sc_hd__xor2_1_93/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_49 sky130_fd_sc_hd__buf_12_49/A sky130_fd_sc_hd__buf_12_49/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__o21ai_2_14 sky130_fd_sc_hd__o21ai_2_14/B1 sky130_fd_sc_hd__o21ai_2_14/Y
+ sky130_fd_sc_hd__xor2_1_543/A sky130_fd_sc_hd__nor2_2_25/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__o21ai_2
Xsky130_fd_sc_hd__xor2_1_580 sky130_fd_sc_hd__xor2_1_580/B sky130_fd_sc_hd__xor2_1_580/X
+ sky130_fd_sc_hd__xor2_1_580/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_591 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__xor2_1_591/X
+ sky130_fd_sc_hd__xor2_1_591/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a222oi_1_600 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_418/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_450/Q sky130_fd_sc_hd__nor2_4_19/B
+ sky130_fd_sc_hd__clkinv_1_797/A sky130_fd_sc_hd__dfxtp_1_386/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__maj3_1_1 sky130_fd_sc_hd__maj3_1_1/C sky130_fd_sc_hd__maj3_1_1/X
+ sky130_fd_sc_hd__maj3_1_1/B sky130_fd_sc_hd__maj3_1_1/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__and2_0_10 vccd1 vssd1 sky130_fd_sc_hd__and2_0_10/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_21 vccd1 vssd1 sky130_fd_sc_hd__and2_0_21/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__buf_2_30/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_32 vccd1 vssd1 sky130_fd_sc_hd__and2_0_32/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__or2_0_53/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_43 vccd1 vssd1 sky130_fd_sc_hd__and2_0_43/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__buf_2_20/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_54 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_2_3/D sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__nor2_2_4/B vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_65 vccd1 vssd1 sky130_fd_sc_hd__and2_0_65/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__or2_0_66/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_76 vccd1 vssd1 sky130_fd_sc_hd__and2_0_76/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__buf_4_5/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_409 sky130_fd_sc_hd__xnor2_2_0/B sky130_fd_sc_hd__nand2_1_410/Y
+ sky130_fd_sc_hd__nand2_1_409/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2_2_2 sky130_fd_sc_hd__nor2_2_2/B sky130_fd_sc_hd__nor2_2_2/Y
+ sky130_fd_sc_hd__nor2_2_2/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__and2_0_87 vccd1 vssd1 sky130_fd_sc_hd__and2_0_87/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__and2_0_87/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_98 vccd1 vssd1 sky130_fd_sc_hd__and2_0_98/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__or2_0_61/B vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_8_20 sky130_fd_sc_hd__buf_8_20/A sky130_fd_sc_hd__buf_8_20/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_31 sky130_fd_sc_hd__buf_8_31/A sky130_fd_sc_hd__buf_8_31/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_42 sky130_fd_sc_hd__buf_8_42/A sky130_fd_sc_hd__buf_8_42/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_53 sky130_fd_sc_hd__buf_8_53/A sky130_fd_sc_hd__buf_8_53/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_64 sky130_fd_sc_hd__buf_8_64/A sky130_fd_sc_hd__buf_8_64/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_75 sky130_fd_sc_hd__buf_8_75/A sky130_fd_sc_hd__buf_8_75/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_86 sky130_fd_sc_hd__buf_8_86/A sky130_fd_sc_hd__buf_8_86/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_205 sky130_fd_sc_hd__xor2_1_557/A sky130_fd_sc_hd__dfxtp_2_2/CLK
+ sky130_fd_sc_hd__and2_0_72/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_8_97 sky130_fd_sc_hd__buf_8_97/A sky130_fd_sc_hd__buf_8_97/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_216 sky130_fd_sc_hd__xnor2_1_134/A sky130_fd_sc_hd__dfxtp_1_217/CLK
+ sky130_fd_sc_hd__and2_0_100/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_227 sky130_fd_sc_hd__xnor2_1_109/A sky130_fd_sc_hd__dfxtp_1_230/CLK
+ sky130_fd_sc_hd__and2_0_38/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_238 sky130_fd_sc_hd__fa_2_217/A sky130_fd_sc_hd__dfxtp_2_5/CLK
+ sky130_fd_sc_hd__and2_0_63/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_249 sky130_fd_sc_hd__xnor2_1_61/A sky130_fd_sc_hd__clkinv_4_6/Y
+ sky130_fd_sc_hd__and2_0_27/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_550 vssd1 vccd1 sky130_fd_sc_hd__inv_2_34/Y sky130_fd_sc_hd__nand2b_2_3/Y
+ sky130_fd_sc_hd__o21ai_1_550/B1 sky130_fd_sc_hd__xor2_1_348/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_561 vssd1 vccd1 sky130_fd_sc_hd__inv_2_42/Y sky130_fd_sc_hd__nand2_1_416/Y
+ sky130_fd_sc_hd__a21oi_1_86/Y sky130_fd_sc_hd__xnor2_1_100/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_572 vssd1 vccd1 sky130_fd_sc_hd__inv_2_30/Y sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_572/B1 sky130_fd_sc_hd__xor2_1_369/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_583 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_384/A sky130_fd_sc_hd__nor2_1_147/Y
+ sky130_fd_sc_hd__nand2_1_442/Y sky130_fd_sc_hd__xnor2_1_107/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_594 vssd1 vccd1 sky130_fd_sc_hd__inv_2_34/Y sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_594/B1 sky130_fd_sc_hd__xor2_1_388/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__buf_2_105 vccd1 vssd1 sky130_fd_sc_hd__buf_2_105/X sky130_fd_sc_hd__buf_2_105/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_116 vccd1 vssd1 sky130_fd_sc_hd__buf_2_116/X sky130_fd_sc_hd__buf_2_116/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_127 vccd1 vssd1 sky130_fd_sc_hd__buf_2_127/X sky130_fd_sc_hd__buf_2_127/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_138 vccd1 vssd1 sky130_fd_sc_hd__buf_2_138/X sky130_fd_sc_hd__buf_2_138/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_149 vccd1 vssd1 sky130_fd_sc_hd__buf_2_149/X sky130_fd_sc_hd__buf_2_149/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__ha_2_5 vssd1 vccd1 sky130_fd_sc_hd__ha_2_5/A sky130_fd_sc_hd__ha_2_5/COUT
+ sky130_fd_sc_hd__ha_2_5/SUM sky130_fd_sc_hd__ha_2_5/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__nand2b_2_10 la_data_out[36] sky130_fd_sc_hd__nand2b_2_10/Y la_data_out[47]
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_2
Xsky130_fd_sc_hd__a222oi_1_430 vccd1 vssd1 sky130_fd_sc_hd__and3_4_26/X sky130_fd_sc_hd__buf_2_4/A
+ sky130_fd_sc_hd__buf_2_20/X sky130_fd_sc_hd__nor2_2_31/Y sky130_fd_sc_hd__buf_2_21/X
+ sky130_fd_sc_hd__o21ai_1_704/B1 sky130_fd_sc_hd__nor2b_1_12/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_441 vccd1 vssd1 sky130_fd_sc_hd__and3_4_18/X sky130_fd_sc_hd__buf_2_21/X
+ sky130_fd_sc_hd__nor2_1_87/A sky130_fd_sc_hd__nor2_2_32/Y sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__o21ai_1_719/B1 sky130_fd_sc_hd__nor2b_2_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_452 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__buf_4_2/X sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__o21ai_1_732/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_463 vccd1 vssd1 sky130_fd_sc_hd__and3_4_20/X sky130_fd_sc_hd__buf_2_21/X
+ sky130_fd_sc_hd__nor2_1_87/A sky130_fd_sc_hd__nor2_4_16/Y sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__o21ai_1_747/B1 sky130_fd_sc_hd__and2b_4_11/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_474 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__buf_6_4/X
+ sky130_fd_sc_hd__buf_6_0/X sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__o21ai_1_761/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_16 vssd1 vccd1 sky130_fd_sc_hd__nand2_1_129/A sky130_fd_sc_hd__xnor2_1_113/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_485 vccd1 vssd1 sky130_fd_sc_hd__and3_4_26/X sky130_fd_sc_hd__or2_0_71/B
+ sky130_fd_sc_hd__buf_2_29/X sky130_fd_sc_hd__nor2_2_31/Y sky130_fd_sc_hd__buf_2_30/X
+ sky130_fd_sc_hd__o21ai_1_774/B1 sky130_fd_sc_hd__nor2b_1_12/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_27 vssd1 vccd1 sky130_fd_sc_hd__and2_0_38/A sky130_fd_sc_hd__nor2_1_87/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_496 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__nor2_1_85/B sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__nor2_2_10/B
+ sky130_fd_sc_hd__o21ai_1_789/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_38 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_38/X sky130_fd_sc_hd__buf_2_38/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_49 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_49/X sky130_fd_sc_hd__clkbuf_1_49/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__or2_0_18 sky130_fd_sc_hd__buf_4_3/X sky130_fd_sc_hd__or2_0_18/X
+ sky130_fd_sc_hd__buf_4_2/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__or2_0_29 sky130_fd_sc_hd__or2_0_29/A sky130_fd_sc_hd__or2_0_29/X
+ sky130_fd_sc_hd__or2_0_29/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__and2_0_390 vccd1 vssd1 sky130_fd_sc_hd__and2_0_390/X sky130_fd_sc_hd__and2_0_401/B
+ sky130_fd_sc_hd__and2_0_390/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_12_5 sky130_fd_sc_hd__buf_12_5/A sky130_fd_sc_hd__buf_12_5/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_605 sky130_fd_sc_hd__buf_12_605/A sky130_fd_sc_hd__buf_12_605/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_616 sky130_fd_sc_hd__buf_12_616/A sky130_fd_sc_hd__buf_12_616/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_627 sky130_fd_sc_hd__buf_12_627/A sky130_fd_sc_hd__buf_12_627/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_638 sky130_fd_sc_hd__buf_12_638/A sky130_fd_sc_hd__buf_12_638/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__inv_2_190 sky130_fd_sc_hd__inv_2_190/A sky130_fd_sc_hd__inv_2_190/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__clkinv_4_109 sky130_fd_sc_hd__clkinv_4_109/A sky130_fd_sc_hd__clkinv_4_110/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_12_649 sky130_fd_sc_hd__buf_12_649/A sky130_fd_sc_hd__buf_12_649/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__o22ai_1_120 sky130_fd_sc_hd__nor2b_1_20/A sky130_fd_sc_hd__xnor2_1_267/Y
+ sky130_fd_sc_hd__fa_2_450/B sky130_fd_sc_hd__xnor2_1_270/Y sky130_fd_sc_hd__o22ai_1_78/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_131 sky130_fd_sc_hd__xnor2_2_6/Y sky130_fd_sc_hd__xnor2_1_279/Y
+ sky130_fd_sc_hd__fa_2_456/B sky130_fd_sc_hd__xnor2_1_282/Y sky130_fd_sc_hd__o22ai_1_98/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_206 sky130_fd_sc_hd__xor2_1_83/B sky130_fd_sc_hd__nand2_1_207/Y
+ sky130_fd_sc_hd__nand2_1_206/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_805 sky130_fd_sc_hd__fa_2_466/CIN sky130_fd_sc_hd__a21oi_1_169/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_217 sky130_fd_sc_hd__xor2_1_100/B sky130_fd_sc_hd__nand2_1_218/Y
+ sky130_fd_sc_hd__nand2_1_217/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_816 sky130_fd_sc_hd__clkinv_1_816/Y sky130_fd_sc_hd__nand2_1_811/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_2_20 sky130_fd_sc_hd__nor2_2_20/B sky130_fd_sc_hd__nor2_2_20/Y
+ sky130_fd_sc_hd__nor2_2_20/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__nand2_1_228 sky130_fd_sc_hd__o21ai_2_8/B1 sky130_fd_sc_hd__nor2_1_69/A
+ sky130_fd_sc_hd__nor2_1_69/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_827 sky130_fd_sc_hd__nand2_1_832/A sky130_fd_sc_hd__nor2_1_264/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_2_31 sky130_fd_sc_hd__nor2_2_31/B sky130_fd_sc_hd__nor2_2_31/Y
+ sky130_fd_sc_hd__nor2_2_31/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__nand2_1_239 sky130_fd_sc_hd__nand2_1_239/Y sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__nor2_1_73/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_838 sky130_fd_sc_hd__buf_8_87/A sky130_fd_sc_hd__clkinv_1_839/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_849 sky130_fd_sc_hd__clkinv_1_849/Y sky130_fd_sc_hd__clkinv_8_8/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__conb_1_16 sky130_fd_sc_hd__conb_1_16/LO sky130_fd_sc_hd__conb_1_16/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_27 sky130_fd_sc_hd__conb_1_27/LO sky130_fd_sc_hd__conb_1_27/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_38 sky130_fd_sc_hd__conb_1_38/LO sky130_fd_sc_hd__conb_1_38/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_49 sky130_fd_sc_hd__conb_1_49/LO sky130_fd_sc_hd__conb_1_49/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__o21ai_1_380 vssd1 vccd1 sky130_fd_sc_hd__buf_2_3/X sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__o21ai_1_380/B1 sky130_fd_sc_hd__xor2_1_195/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_391 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_103/Y sky130_fd_sc_hd__o21a_1_1/X
+ sky130_fd_sc_hd__nand2_1_314/Y sky130_fd_sc_hd__xnor2_1_60/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_801 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_812 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_823 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_834 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_845 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_856 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_740 sky130_fd_sc_hd__nand2_1_740/Y sky130_fd_sc_hd__or2_0_89/A
+ sky130_fd_sc_hd__or2_0_89/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_867 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_751 sky130_fd_sc_hd__xor2_1_658/A sky130_fd_sc_hd__nand2_1_752/Y
+ sky130_fd_sc_hd__nand2_1_751/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_878 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_762 sky130_fd_sc_hd__xnor2_1_215/A sky130_fd_sc_hd__nand2_1_778/Y
+ sky130_fd_sc_hd__or2_0_93/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_889 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_773 sky130_fd_sc_hd__nand2_1_773/Y sky130_fd_sc_hd__nor2_1_244/A
+ sky130_fd_sc_hd__nor2_1_244/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_784 sky130_fd_sc_hd__nand2_1_784/Y sky130_fd_sc_hd__o22ai_1_86/Y
+ sky130_fd_sc_hd__ha_2_14/SUM vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_795 sky130_fd_sc_hd__nand2_1_795/Y sky130_fd_sc_hd__or2_0_100/A
+ sky130_fd_sc_hd__or2_0_100/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_1800 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1811 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1822 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1833 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1844 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1855 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1866 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_260 vccd1 vssd1 sky130_fd_sc_hd__and3_4_14/X sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__buf_4_7/X sky130_fd_sc_hd__nor2_1_127/Y sky130_fd_sc_hd__buf_4_0/X
+ sky130_fd_sc_hd__o21ai_1_462/B1 sky130_fd_sc_hd__nor2b_1_10/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_271 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__buf_4_5/X sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__o21ai_1_475/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_282 vccd1 vssd1 sky130_fd_sc_hd__and3_4_14/X sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__inv_6_0/Y sky130_fd_sc_hd__nor2_1_127/Y sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__o21ai_1_489/B1 sky130_fd_sc_hd__nor2b_1_10/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_430 sky130_fd_sc_hd__nor2_1_244/A sky130_fd_sc_hd__nor2_1_246/B
+ sky130_fd_sc_hd__fa_2_430/A sky130_fd_sc_hd__fa_2_430/B sky130_fd_sc_hd__fa_2_430/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_293 vccd1 vssd1 sky130_fd_sc_hd__and3_4_14/X sky130_fd_sc_hd__or2_0_52/B
+ sky130_fd_sc_hd__or2_0_53/A sky130_fd_sc_hd__nor2_1_127/Y sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__o21ai_1_503/B1 sky130_fd_sc_hd__nor2b_1_10/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_441 sky130_fd_sc_hd__fa_2_437/B sky130_fd_sc_hd__fa_2_441/SUM
+ sky130_fd_sc_hd__fa_2_441/A sky130_fd_sc_hd__fa_2_441/B sky130_fd_sc_hd__ha_2_13/COUT
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_452 sky130_fd_sc_hd__fa_2_452/COUT sky130_fd_sc_hd__fa_2_451/B
+ sky130_fd_sc_hd__fa_2_452/A sky130_fd_sc_hd__fa_2_452/B sky130_fd_sc_hd__fa_2_452/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_463 sky130_fd_sc_hd__fa_2_460/B sky130_fd_sc_hd__fa_2_462/A
+ sky130_fd_sc_hd__fa_2_463/A sky130_fd_sc_hd__fa_2_463/B sky130_fd_sc_hd__nor2b_1_29/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_474 sky130_fd_sc_hd__nor2_1_256/B sky130_fd_sc_hd__or2_0_102/A
+ sky130_fd_sc_hd__fa_2_474/A sky130_fd_sc_hd__fa_2_474/B sky130_fd_sc_hd__nor2b_1_47/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_485 sky130_fd_sc_hd__or2_0_107/B sky130_fd_sc_hd__nor2_1_262/A
+ sky130_fd_sc_hd__fa_2_485/A sky130_fd_sc_hd__fa_2_485/B sky130_fd_sc_hd__nor2b_1_69/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__decap_8_13 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__nor2_1_206 sky130_fd_sc_hd__nor2_1_206/B sky130_fd_sc_hd__nor2_1_206/Y
+ sky130_fd_sc_hd__nor2_1_206/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_217 sky130_fd_sc_hd__buf_2_29/X sky130_fd_sc_hd__nor2_1_217/Y
+ sky130_fd_sc_hd__buf_2_30/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_228 sky130_fd_sc_hd__mux2_2_46/X sky130_fd_sc_hd__nor2_1_228/Y
+ sky130_fd_sc_hd__mux2_2_31/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_239 sky130_fd_sc_hd__xor2_1_664/X sky130_fd_sc_hd__nor2_1_239/Y
+ sky130_fd_sc_hd__nor2_1_239/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_402 sky130_fd_sc_hd__buf_12_402/A sky130_fd_sc_hd__buf_12_570/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_413 sky130_fd_sc_hd__buf_12_413/A sky130_fd_sc_hd__buf_12_488/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_424 sky130_fd_sc_hd__buf_12_424/A sky130_fd_sc_hd__buf_12_481/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_435 sky130_fd_sc_hd__buf_12_75/X sky130_fd_sc_hd__buf_12_480/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_446 sky130_fd_sc_hd__buf_12_446/A sky130_fd_sc_hd__buf_12_634/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_457 sky130_fd_sc_hd__buf_12_457/A sky130_fd_sc_hd__buf_12_640/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_468 sky130_fd_sc_hd__buf_12_468/A sky130_fd_sc_hd__buf_12_650/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_479 sky130_fd_sc_hd__buf_12_479/A sky130_fd_sc_hd__buf_12_524/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_108 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_119 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_602 sky130_fd_sc_hd__clkinv_1_602/Y sky130_fd_sc_hd__nand2_1_645/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_613 sky130_fd_sc_hd__and3_4_19/A sky130_fd_sc_hd__xor2_1_637/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_624 sky130_fd_sc_hd__fa_2_419/CIN sky130_fd_sc_hd__a21oi_1_138/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_635 sky130_fd_sc_hd__clkinv_1_635/Y sky130_fd_sc_hd__nand2_1_683/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_646 sky130_fd_sc_hd__nand2_1_704/A sky130_fd_sc_hd__nor2_1_231/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_209 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_209/B sky130_fd_sc_hd__a22o_1_13/B1
+ sky130_fd_sc_hd__xnor2_1_209/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_657 sky130_fd_sc_hd__o22ai_1_103/B1 sky130_fd_sc_hd__or2_0_79/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_668 sky130_fd_sc_hd__clkinv_1_668/Y sky130_fd_sc_hd__nand2_1_738/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_679 sky130_fd_sc_hd__xor2_1_659/A sky130_fd_sc_hd__o21ai_1_884/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1107 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1118 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1129 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_11 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_352/Q sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__o211ai_1_27/Y sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__a222oi_1_11/Y sky130_fd_sc_hd__dfxtp_1_303/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_22 vccd1 vssd1 sky130_fd_sc_hd__xnor2_1_123/Y sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__xnor2_1_185/Y sky130_fd_sc_hd__xnor2_1_60/Y sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_22/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_33 vccd1 vssd1 sky130_fd_sc_hd__xor2_1_367/X sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__xor2_1_580/X sky130_fd_sc_hd__xor2_1_154/X sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_33/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_620 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_44 vccd1 vssd1 sky130_fd_sc_hd__xor2_1_296/X sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__inv_2_56/A sky130_fd_sc_hd__xor2_1_83/X sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_44/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_631 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_55 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__or2_0_42/B
+ sky130_fd_sc_hd__or2_0_39/B sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__or2_0_58/A
+ sky130_fd_sc_hd__a222oi_1_55/Y sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_642 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_66 vccd1 vssd1 sky130_fd_sc_hd__and3_4_1/X sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__buf_4_4/X sky130_fd_sc_hd__nor2_2_9/Y sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__a222oi_1_66/Y sky130_fd_sc_hd__and2b_4_3/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_653 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_13 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_13/B sky130_fd_sc_hd__xnor2_1_13/Y
+ sky130_fd_sc_hd__xnor2_1_13/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__a222oi_1_77 vccd1 vssd1 sky130_fd_sc_hd__and3_4_5/X sky130_fd_sc_hd__nor2_2_5/A
+ sky130_fd_sc_hd__nor2_2_5/B sky130_fd_sc_hd__nor2_1_68/Y sky130_fd_sc_hd__nor2_2_4/B
+ sky130_fd_sc_hd__a222oi_1_77/Y sky130_fd_sc_hd__nor2b_1_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_664 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_24 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_24/B sky130_fd_sc_hd__inv_2_14/A
+ sky130_fd_sc_hd__xnor2_1_24/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__a222oi_1_88 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__or2_0_60/B sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__or2_0_60/A
+ sky130_fd_sc_hd__a222oi_1_88/Y sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_675 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_99 vccd1 vssd1 sky130_fd_sc_hd__and3_4_8/X sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__nor2_1_85/B sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__nor2_2_10/B
+ sky130_fd_sc_hd__a222oi_1_99/Y sky130_fd_sc_hd__nor2b_2_2/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__xnor2_1_35 vssd1 vccd1 sky130_fd_sc_hd__o21ai_2_7/Y sky130_fd_sc_hd__xnor2_1_35/Y
+ sky130_fd_sc_hd__xnor2_1_35/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_46 vssd1 vccd1 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__nor2_2_8/A
+ sky130_fd_sc_hd__xnor2_1_46/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_686 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_570 sky130_fd_sc_hd__xor2_1_543/B sky130_fd_sc_hd__o21ai_2_14/B1
+ sky130_fd_sc_hd__nand2_1_570/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_697 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_57 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_57/B sky130_fd_sc_hd__xnor2_1_57/Y
+ sky130_fd_sc_hd__xnor2_1_57/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_581 sky130_fd_sc_hd__xnor2_1_126/B sky130_fd_sc_hd__nand2_1_582/Y
+ sky130_fd_sc_hd__nand2_1_581/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_68 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_71/A sky130_fd_sc_hd__nor2b_1_7/A
+ sky130_fd_sc_hd__xnor2_1_68/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xor2_1_409 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__nor2_4_13/B
+ sky130_fd_sc_hd__xor2_1_409/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_592 sky130_fd_sc_hd__nand2_1_592/Y sky130_fd_sc_hd__or2_1_1/A
+ sky130_fd_sc_hd__or2_1_1/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_79 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_79/B sky130_fd_sc_hd__xnor2_1_79/Y
+ sky130_fd_sc_hd__xnor2_1_79/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_1150 sky130_fd_sc_hd__buf_2_47/A sky130_fd_sc_hd__clkinv_4_89/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_2_2 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_2/Y sky130_fd_sc_hd__xnor2_2_2/A
+ sky130_fd_sc_hd__xnor2_2_2/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_2
Xsky130_fd_sc_hd__decap_12_1630 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1641 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1652 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1663 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1674 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1685 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1696 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__fa_2_260 sky130_fd_sc_hd__fa_2_257/A sky130_fd_sc_hd__fa_2_263/A
+ sky130_fd_sc_hd__fa_2_260/A sky130_fd_sc_hd__fa_2_260/B sky130_fd_sc_hd__fa_2_260/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_271 sky130_fd_sc_hd__fa_2_269/A sky130_fd_sc_hd__fa_2_272/CIN
+ sky130_fd_sc_hd__fa_2_271/A sky130_fd_sc_hd__fa_2_271/B sky130_fd_sc_hd__fa_2_271/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_282 sky130_fd_sc_hd__xor2_1_426/B sky130_fd_sc_hd__or2_1_9/B
+ sky130_fd_sc_hd__fa_2_282/A sky130_fd_sc_hd__fa_2_282/B sky130_fd_sc_hd__fa_2_287/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor4_1_5 wbs_adr_i[27] wbs_adr_i[25] sky130_fd_sc_hd__nor4_1_5/Y
+ wbs_adr_i[26] wbs_adr_i[24] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor4_1
Xsky130_fd_sc_hd__fa_2_293 sky130_fd_sc_hd__fa_2_283/A sky130_fd_sc_hd__fa_2_296/CIN
+ sky130_fd_sc_hd__fa_2_293/A sky130_fd_sc_hd__fa_2_293/B sky130_fd_sc_hd__xor2_1_453/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22oi_1_4 sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__a22oi_1_4/B2 sky130_fd_sc_hd__a22oi_1_4/A2 sky130_fd_sc_hd__nand2_2_1/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__decap_12_9 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_210 sky130_fd_sc_hd__buf_6_51/X sky130_fd_sc_hd__buf_12_412/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_221 sky130_fd_sc_hd__buf_6_80/X sky130_fd_sc_hd__buf_12_399/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_232 sky130_fd_sc_hd__bufinv_8_1/Y sky130_fd_sc_hd__buf_12_313/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_243 sky130_fd_sc_hd__buf_6_39/X sky130_fd_sc_hd__buf_12_373/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_90 sky130_fd_sc_hd__xnor2_1_104/B sky130_fd_sc_hd__a21oi_1_90/B1
+ sky130_fd_sc_hd__xor2_1_367/A sky130_fd_sc_hd__nand2_1_430/A vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_1_102 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_183/Q sky130_fd_sc_hd__dfxtp_1_151/Q sky130_fd_sc_hd__o21ai_1_8/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_254 sky130_fd_sc_hd__buf_6_24/X sky130_fd_sc_hd__buf_12_290/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_113 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_173/Q sky130_fd_sc_hd__dfxtp_1_141/Q sky130_fd_sc_hd__o21ai_1_19/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_265 sky130_fd_sc_hd__buf_6_50/X sky130_fd_sc_hd__buf_12_426/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_124 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_162/Q sky130_fd_sc_hd__dfxtp_1_130/Q sky130_fd_sc_hd__o21ai_1_30/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_276 sky130_fd_sc_hd__buf_12_276/A sky130_fd_sc_hd__buf_12_605/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_135 sky130_fd_sc_hd__xnor2_1_73/Y sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xnor2_1_10/Y sky130_fd_sc_hd__o21ai_1_49/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_287 sky130_fd_sc_hd__buf_12_287/A sky130_fd_sc_hd__buf_12_287/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_146 sky130_fd_sc_hd__xnor2_1_86/Y sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xnor2_1_23/Y sky130_fd_sc_hd__o21ai_1_72/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_298 sky130_fd_sc_hd__buf_12_298/A sky130_fd_sc_hd__buf_8_165/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_157 sky130_fd_sc_hd__xor2_1_346/X sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xor2_1_133/X sky130_fd_sc_hd__o21ai_1_93/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_168 sky130_fd_sc_hd__xor2_1_384/X sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xor2_1_171/X sky130_fd_sc_hd__a22oi_1_168/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_410 sky130_fd_sc_hd__nand2_1_458/A sky130_fd_sc_hd__nor2_2_16/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22oi_1_179 sky130_fd_sc_hd__nand2_1_135/A sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xnor2_1_54/Y sky130_fd_sc_hd__a22oi_1_179/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_421 sky130_fd_sc_hd__nand2_1_344/A sky130_fd_sc_hd__nor2_1_110/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_432 sky130_fd_sc_hd__nor2_1_114/A sky130_fd_sc_hd__nand2_1_371/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_443 sky130_fd_sc_hd__o21ai_1_486/A2 sky130_fd_sc_hd__xnor2_1_83/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_454 sky130_fd_sc_hd__o21ai_1_515/B1 sky130_fd_sc_hd__o21ai_1_516/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_465 sky130_fd_sc_hd__nand2_1_409/A sky130_fd_sc_hd__nor2_1_131/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_476 sky130_fd_sc_hd__a21oi_1_90/B1 sky130_fd_sc_hd__nand2_1_431/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_487 sky130_fd_sc_hd__xor2_1_384/A sky130_fd_sc_hd__o21ai_1_595/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_498 sky130_fd_sc_hd__a21oi_1_99/B1 sky130_fd_sc_hd__nand2_1_471/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_2_14 sky130_fd_sc_hd__buf_4_8/A sky130_fd_sc_hd__nand2_2_14/A
+ sky130_fd_sc_hd__dfxtp_1_0/Q vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__decap_12_450 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_461 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_472 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_483 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_494 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_206 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__and3_4_3/A
+ sky130_fd_sc_hd__xor2_1_206/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_217 sky130_fd_sc_hd__fa_2_239/A sky130_fd_sc_hd__xor3_1_13/A
+ sky130_fd_sc_hd__xor2_1_217/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_228 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__xor2_1_228/X
+ sky130_fd_sc_hd__xor2_1_228/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_239 sky130_fd_sc_hd__dfxtp_2_5/Q sky130_fd_sc_hd__fa_2_152/A
+ sky130_fd_sc_hd__xor2_1_239/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1460 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1471 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_902 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_685/A sky130_fd_sc_hd__nor2_1_263/Y
+ sky130_fd_sc_hd__nand2_1_829/Y sky130_fd_sc_hd__xnor2_1_299/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1482 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_913 vssd1 vccd1 sky130_fd_sc_hd__nor2_2_1/B sky130_fd_sc_hd__o21ai_1_913/A1
+ sky130_fd_sc_hd__a31oi_1_2/Y sky130_fd_sc_hd__o21ai_1_913/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1493 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_924 vssd1 vccd1 sky130_fd_sc_hd__nand2_1_865/B sky130_fd_sc_hd__a21o_2_3/B1
+ sky130_fd_sc_hd__a21o_2_4/A2 sky130_fd_sc_hd__inv_2_114/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_8_6 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__buf_2_11 vccd1 vssd1 sky130_fd_sc_hd__buf_2_11/X sky130_fd_sc_hd__buf_2_11/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_22 vccd1 vssd1 sky130_fd_sc_hd__buf_2_22/X sky130_fd_sc_hd__buf_2_22/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_33 vccd1 vssd1 sky130_fd_sc_hd__buf_8_90/A sky130_fd_sc_hd__buf_8_88/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_44 vccd1 vssd1 sky130_fd_sc_hd__buf_2_44/X sky130_fd_sc_hd__buf_2_44/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_55 vccd1 vssd1 sky130_fd_sc_hd__buf_8_91/A sky130_fd_sc_hd__inv_12_0/Y
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_66 vccd1 vssd1 sky130_fd_sc_hd__buf_6_8/A sky130_fd_sc_hd__buf_2_66/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_77 vccd1 vssd1 sky130_fd_sc_hd__buf_2_77/X sky130_fd_sc_hd__buf_2_77/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_88 vccd1 vssd1 sky130_fd_sc_hd__buf_2_88/X sky130_fd_sc_hd__buf_2_88/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_99 vccd1 vssd1 sky130_fd_sc_hd__buf_2_99/X sky130_fd_sc_hd__buf_2_99/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o211ai_1_60 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o22ai_1_3/B1
+ sky130_fd_sc_hd__fa_2_414/B sky130_fd_sc_hd__nand2_1_80/Y sky130_fd_sc_hd__a21oi_1_31/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__diode_2_6 sky130_fd_sc_hd__inv_12_0/Y vssd1 vccd1 vccd1 vssd1 sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__and2_0_208 vccd1 vssd1 sky130_fd_sc_hd__and2_0_208/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_76/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_219 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_54/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_67/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__xor3_1_17 sky130_fd_sc_hd__xor3_1_17/X sky130_fd_sc_hd__xor3_1_18/X
+ sky130_fd_sc_hd__xor3_1_17/B sky130_fd_sc_hd__xor3_1_17/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__xor3_1_28 sky130_fd_sc_hd__xor3_1_28/X sky130_fd_sc_hd__xor3_1_28/C
+ sky130_fd_sc_hd__xor3_1_28/B sky130_fd_sc_hd__xor3_1_28/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__clkinv_1_240 sky130_fd_sc_hd__o22ai_1_0/B1 sky130_fd_sc_hd__dfxtp_1_95/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_251 sky130_fd_sc_hd__o21ai_1_93/A2 sky130_fd_sc_hd__xor2_1_559/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_262 sky130_fd_sc_hd__o21ai_1_137/A2 sky130_fd_sc_hd__xnor2_1_179/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_273 sky130_fd_sc_hd__and2_0_148/A sky130_fd_sc_hd__a222oi_1_17/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_284 sky130_fd_sc_hd__and2_0_211/A sky130_fd_sc_hd__a222oi_1_28/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_295 sky130_fd_sc_hd__and2_0_156/A sky130_fd_sc_hd__a222oi_1_39/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xor3_1_2 sky130_fd_sc_hd__xor3_1_2/X sky130_fd_sc_hd__xor3_1_2/C
+ sky130_fd_sc_hd__xor3_1_3/X sky130_fd_sc_hd__xor3_1_2/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__a21oi_1_3 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_32/Y
+ sky130_fd_sc_hd__a21oi_1_3/Y sky130_fd_sc_hd__dfxtp_1_92/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkbuf_4_16 sky130_fd_sc_hd__buf_6_11/A sky130_fd_sc_hd__clkbuf_4_16/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and3_4_20 sky130_fd_sc_hd__nor2_4_16/B sky130_fd_sc_hd__nor2_4_16/A
+ sky130_fd_sc_hd__and3_4_20/C sky130_fd_sc_hd__and3_4_20/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__o21ai_1_209 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_209/A2 sky130_fd_sc_hd__nor2_1_55/Y
+ sky130_fd_sc_hd__nand2_1_189/Y sky130_fd_sc_hd__o21ai_1_209/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_27 sky130_fd_sc_hd__clkbuf_4_27/X sky130_fd_sc_hd__buf_8_15/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_38 la_data_out[63] sky130_fd_sc_hd__dfxtp_1_478/Q vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_49 la_data_out[85] sky130_fd_sc_hd__or2_0_80/A vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__a21oi_1_170 sky130_fd_sc_hd__xnor2_1_291/B sky130_fd_sc_hd__clkinv_1_808/Y
+ sky130_fd_sc_hd__xor2_1_676/A sky130_fd_sc_hd__or2_0_100/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_181 sky130_fd_sc_hd__xnor2_1_302/A sky130_fd_sc_hd__clkinv_1_830/Y
+ sky130_fd_sc_hd__xor2_1_687/A sky130_fd_sc_hd__or2_0_111/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_192 sky130_fd_sc_hd__ha_2_32/A la_data_out[39] sky130_fd_sc_hd__a21oi_1_192/Y
+ sky130_fd_sc_hd__ha_2_48/B vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_100 sky130_fd_sc_hd__buf_8_100/A sky130_fd_sc_hd__buf_8_100/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_111 sky130_fd_sc_hd__buf_8_111/A sky130_fd_sc_hd__buf_8_111/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_122 sky130_fd_sc_hd__inv_2_164/Y sky130_fd_sc_hd__buf_8_122/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_133 sky130_fd_sc_hd__buf_8_133/A sky130_fd_sc_hd__buf_8_133/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_144 sky130_fd_sc_hd__buf_8_144/A sky130_fd_sc_hd__buf_8_144/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nor2_4_6 sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__nor2_4_6/A
+ sky130_fd_sc_hd__nor2_4_7/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__buf_8_155 sky130_fd_sc_hd__buf_8_155/A sky130_fd_sc_hd__buf_6_82/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__decap_12_280 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_291 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_409 sky130_fd_sc_hd__dfxtp_1_409/Q sky130_fd_sc_hd__dfxtp_1_410/CLK
+ sky130_fd_sc_hd__nor2b_1_106/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_710 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_10/X sky130_fd_sc_hd__nand2_1_535/Y
+ sky130_fd_sc_hd__a21oi_1_113/Y sky130_fd_sc_hd__xnor2_1_142/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1290 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_721 vssd1 vccd1 sky130_fd_sc_hd__inv_2_50/Y sky130_fd_sc_hd__nand2b_2_6/Y
+ sky130_fd_sc_hd__o21ai_1_721/B1 sky130_fd_sc_hd__xor2_1_498/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_732 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_767/A2 sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_732/B1 sky130_fd_sc_hd__xor2_1_510/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_743 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_10/X sky130_fd_sc_hd__nand2_1_557/Y
+ sky130_fd_sc_hd__a21oi_1_117/Y sky130_fd_sc_hd__xnor2_1_150/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_754 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_2/Y sky130_fd_sc_hd__nand2b_1_21/Y
+ sky130_fd_sc_hd__o21ai_1_754/B1 sky130_fd_sc_hd__xor2_1_528/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_765 vssd1 vccd1 sky130_fd_sc_hd__buf_2_13/X sky130_fd_sc_hd__nand2b_1_21/Y
+ sky130_fd_sc_hd__o21ai_1_765/B1 sky130_fd_sc_hd__xor2_1_540/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_776 vssd1 vccd1 sky130_fd_sc_hd__inv_2_44/Y sky130_fd_sc_hd__nand2b_2_6/Y
+ sky130_fd_sc_hd__o21ai_1_776/B1 sky130_fd_sc_hd__xor2_1_550/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_787 vssd1 vccd1 sky130_fd_sc_hd__inv_2_49/Y sky130_fd_sc_hd__nand2b_2_6/Y
+ sky130_fd_sc_hd__o21ai_1_787/B1 sky130_fd_sc_hd__xor2_1_561/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_798 vssd1 vccd1 sky130_fd_sc_hd__inv_2_52/Y sky130_fd_sc_hd__nand2_1_588/Y
+ sky130_fd_sc_hd__a21oi_1_121/Y sky130_fd_sc_hd__xnor2_1_163/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkinv_8_19 sky130_fd_sc_hd__clkinv_8_20/A sky130_fd_sc_hd__clkinv_8_19/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__xor2_1_50 sky130_fd_sc_hd__xor2_1_6/B sky130_fd_sc_hd__fa_2_29/A
+ sky130_fd_sc_hd__xor2_1_50/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_61 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__xor2_1_61/X
+ sky130_fd_sc_hd__xor2_1_61/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_17 sky130_fd_sc_hd__inv_2_75/Y sky130_fd_sc_hd__buf_12_17/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_72 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__fa_2_50/B
+ sky130_fd_sc_hd__xor2_1_72/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_28 sky130_fd_sc_hd__inv_2_135/Y sky130_fd_sc_hd__buf_12_28/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_83 sky130_fd_sc_hd__xor2_1_83/B sky130_fd_sc_hd__xor2_1_83/X
+ sky130_fd_sc_hd__xor2_1_83/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_39 sky130_fd_sc_hd__buf_12_39/A sky130_fd_sc_hd__buf_12_39/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_94 sky130_fd_sc_hd__fa_2_97/A sky130_fd_sc_hd__fa_2_69/B
+ sky130_fd_sc_hd__xor2_1_94/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2b_1_0 sky130_fd_sc_hd__o21ai_2_4/A2 sky130_fd_sc_hd__nand2_1_8/B
+ sky130_fd_sc_hd__nor2_1_0/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__o21ai_2_15 sky130_fd_sc_hd__o21ai_2_15/B1 sky130_fd_sc_hd__o21ai_2_15/Y
+ sky130_fd_sc_hd__xor2_1_559/A sky130_fd_sc_hd__nor2_2_27/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__o21ai_2
Xsky130_fd_sc_hd__xor2_1_570 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__xor2_1_570/X
+ sky130_fd_sc_hd__xor2_1_570/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_581 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__fa_2_394/B
+ sky130_fd_sc_hd__xor2_1_581/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_592 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__fa_2_399/B
+ sky130_fd_sc_hd__xor2_1_592/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a222oi_1_601 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_419/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_451/Q sky130_fd_sc_hd__nor2_4_19/B
+ sky130_fd_sc_hd__clkinv_1_798/A sky130_fd_sc_hd__dfxtp_1_387/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__maj3_1_2 sky130_fd_sc_hd__maj3_1_2/C sky130_fd_sc_hd__maj3_1_2/X
+ sky130_fd_sc_hd__maj3_1_2/B la_data_out[55] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__and2_0_11 vccd1 vssd1 sky130_fd_sc_hd__and2_0_11/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_22 vccd1 vssd1 sky130_fd_sc_hd__and2_0_22/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__buf_6_2/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_33 vccd1 vssd1 sky130_fd_sc_hd__and2_0_33/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__or2_0_72/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_44 vccd1 vssd1 sky130_fd_sc_hd__and2_0_44/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__nor2_1_73/B vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_55 vccd1 vssd1 sky130_fd_sc_hd__and2_0_55/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__buf_2_4/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_66 vccd1 vssd1 sky130_fd_sc_hd__and2_0_66/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__or2_0_61/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_77 vccd1 vssd1 sky130_fd_sc_hd__and2_0_77/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__buf_4_4/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nor2_2_3 sky130_fd_sc_hd__nor2_2_3/B sky130_fd_sc_hd__nor2_2_3/Y
+ sky130_fd_sc_hd__nor2_2_3/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__and2_0_88 vccd1 vssd1 sky130_fd_sc_hd__and2_0_88/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__buf_6_4/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_99 vccd1 vssd1 sky130_fd_sc_hd__and2_0_99/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__or2_0_9/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_8_10 sky130_fd_sc_hd__buf_8_10/A sky130_fd_sc_hd__buf_8_10/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_21 sky130_fd_sc_hd__buf_8_9/X sky130_fd_sc_hd__buf_8_21/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_32 sky130_fd_sc_hd__buf_8_32/A sky130_fd_sc_hd__buf_8_32/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_43 sky130_fd_sc_hd__buf_8_43/A sky130_fd_sc_hd__buf_8_43/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_54 sky130_fd_sc_hd__buf_8_54/A sky130_fd_sc_hd__buf_8_54/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_65 sky130_fd_sc_hd__inv_4_14/Y sky130_fd_sc_hd__buf_8_65/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_76 sky130_fd_sc_hd__buf_8_76/A sky130_fd_sc_hd__buf_8_76/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_87 sky130_fd_sc_hd__buf_8_87/A sky130_fd_sc_hd__buf_8_87/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_206 sky130_fd_sc_hd__fa_2_379/A sky130_fd_sc_hd__dfxtp_2_0/CLK
+ sky130_fd_sc_hd__and2_0_77/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_8_98 sky130_fd_sc_hd__buf_8_98/A sky130_fd_sc_hd__buf_8_98/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_217 sky130_fd_sc_hd__nor2_1_167/A sky130_fd_sc_hd__dfxtp_1_217/CLK
+ sky130_fd_sc_hd__and2_0_59/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_228 sky130_fd_sc_hd__xor2_1_383/A sky130_fd_sc_hd__dfxtp_1_230/CLK
+ sky130_fd_sc_hd__and2_0_49/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_239 sky130_fd_sc_hd__xnor2_1_84/A sky130_fd_sc_hd__clkinv_4_4/Y
+ sky130_fd_sc_hd__and2_0_64/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_540 vssd1 vccd1 sky130_fd_sc_hd__inv_2_32/Y sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_540/B1 sky130_fd_sc_hd__xor2_1_338/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_551 vssd1 vccd1 sky130_fd_sc_hd__inv_2_30/Y sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_551/B1 sky130_fd_sc_hd__xor2_1_349/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_562 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_562/A2 sky130_fd_sc_hd__nor2_1_137/Y
+ sky130_fd_sc_hd__nand2_1_424/Y sky130_fd_sc_hd__o21ai_1_562/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_573 vssd1 vccd1 sky130_fd_sc_hd__inv_2_42/Y sky130_fd_sc_hd__nand2_1_427/Y
+ sky130_fd_sc_hd__a21oi_1_89/Y sky130_fd_sc_hd__xnor2_1_103/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_584 vssd1 vccd1 sky130_fd_sc_hd__inv_2_32/Y sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_584/B1 sky130_fd_sc_hd__xor2_1_378/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_595 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_389/A sky130_fd_sc_hd__nor2_1_149/Y
+ sky130_fd_sc_hd__nand2_1_447/Y sky130_fd_sc_hd__o21ai_1_595/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__buf_2_106 vccd1 vssd1 sky130_fd_sc_hd__buf_2_106/X sky130_fd_sc_hd__buf_2_106/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_117 vccd1 vssd1 sky130_fd_sc_hd__buf_2_117/X sky130_fd_sc_hd__buf_2_117/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_128 vccd1 vssd1 sky130_fd_sc_hd__buf_2_128/X sky130_fd_sc_hd__buf_2_128/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_139 vccd1 vssd1 sky130_fd_sc_hd__buf_2_139/X sky130_fd_sc_hd__buf_2_65/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__ha_2_6 vssd1 vccd1 sky130_fd_sc_hd__ha_2_6/A sky130_fd_sc_hd__ha_2_4/B
+ sky130_fd_sc_hd__nor3_1_0/C sky130_fd_sc_hd__ha_2_6/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__a222oi_1_420 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__or2_0_61/A
+ sky130_fd_sc_hd__or2_0_61/B sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__or2_0_58/B
+ sky130_fd_sc_hd__o21ai_1_691/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_360 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1_1/D sky130_fd_sc_hd__dfxtp_1_2/Q
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_431 vccd1 vssd1 sky130_fd_sc_hd__and3_4_23/X sky130_fd_sc_hd__or2_0_52/B
+ sky130_fd_sc_hd__buf_2_25/A sky130_fd_sc_hd__nor2_1_178/Y sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__o21ai_1_705/B1 sky130_fd_sc_hd__nor2b_1_15/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_442 vccd1 vssd1 sky130_fd_sc_hd__and3_4_26/X sky130_fd_sc_hd__buf_2_15/X
+ sky130_fd_sc_hd__buf_2_4/A sky130_fd_sc_hd__nor2_2_31/Y sky130_fd_sc_hd__buf_2_20/X
+ sky130_fd_sc_hd__o21ai_1_720/B1 sky130_fd_sc_hd__nor2b_1_12/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_453 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__or2_0_66/A sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__or2_0_60/B
+ sky130_fd_sc_hd__o21ai_1_733/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_464 vccd1 vssd1 sky130_fd_sc_hd__and3_4_18/X sky130_fd_sc_hd__buf_2_15/X
+ sky130_fd_sc_hd__buf_2_4/A sky130_fd_sc_hd__nor2_2_32/Y sky130_fd_sc_hd__buf_2_20/X
+ sky130_fd_sc_hd__o21ai_1_748/B1 sky130_fd_sc_hd__nor2b_2_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_475 vccd1 vssd1 sky130_fd_sc_hd__and3_4_18/X sky130_fd_sc_hd__buf_2_24/X
+ sky130_fd_sc_hd__buf_2_27/X sky130_fd_sc_hd__nor2_2_32/Y sky130_fd_sc_hd__buf_2_15/X
+ sky130_fd_sc_hd__o21ai_1_762/B1 sky130_fd_sc_hd__nor2b_2_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_17 vssd1 vccd1 sky130_fd_sc_hd__nand2_1_127/A sky130_fd_sc_hd__xor2_1_389/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_486 vccd1 vssd1 sky130_fd_sc_hd__and3_4_20/X sky130_fd_sc_hd__buf_2_15/X
+ sky130_fd_sc_hd__buf_2_4/A sky130_fd_sc_hd__nor2_4_16/Y sky130_fd_sc_hd__buf_2_20/X
+ sky130_fd_sc_hd__o21ai_1_776/B1 sky130_fd_sc_hd__and2b_4_11/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_28 vssd1 vccd1 sky130_fd_sc_hd__and2_0_49/A sky130_fd_sc_hd__nor2_1_85/B
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_497 vccd1 vssd1 sky130_fd_sc_hd__and3_4_26/X sky130_fd_sc_hd__or2_0_72/B
+ sky130_fd_sc_hd__or2_0_72/A sky130_fd_sc_hd__nor2_2_31/Y sky130_fd_sc_hd__or2_0_71/B
+ sky130_fd_sc_hd__o21ai_1_790/B1 sky130_fd_sc_hd__nor2b_1_12/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_39 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_39/X sky130_fd_sc_hd__a22o_1_79/A2
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__or2_0_19 sky130_fd_sc_hd__buf_4_2/X sky130_fd_sc_hd__or2_0_19/X
+ sky130_fd_sc_hd__buf_4_4/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__and2_0_380 vccd1 vssd1 sky130_fd_sc_hd__and2_0_380/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_54/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_391 vccd1 vssd1 sky130_fd_sc_hd__and2_0_391/X sky130_fd_sc_hd__and2_0_401/B
+ sky130_fd_sc_hd__and2_0_391/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__conb_1_0 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__conb_1_0/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__buf_12_6 sky130_fd_sc_hd__buf_12_6/A sky130_fd_sc_hd__buf_12_6/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_606 sky130_fd_sc_hd__buf_12_606/A sky130_fd_sc_hd__buf_12_606/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_617 sky130_fd_sc_hd__buf_12_617/A sky130_fd_sc_hd__buf_12_617/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_628 sky130_fd_sc_hd__buf_12_628/A sky130_fd_sc_hd__buf_12_628/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__inv_2_180 sky130_fd_sc_hd__inv_2_180/A sky130_fd_sc_hd__inv_2_180/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_12_639 sky130_fd_sc_hd__buf_12_639/A sky130_fd_sc_hd__buf_12_639/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__inv_2_191 sky130_fd_sc_hd__buf_6_88/A sky130_fd_sc_hd__inv_2_191/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__o22ai_1_110 sky130_fd_sc_hd__xnor2_1_260/Y sky130_fd_sc_hd__xnor2_1_259/Y
+ sky130_fd_sc_hd__fa_2_448/B sky130_fd_sc_hd__inv_2_65/Y sky130_fd_sc_hd__o22ai_1_99/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_121 sky130_fd_sc_hd__xnor2_1_271/Y sky130_fd_sc_hd__xnor2_1_268/Y
+ sky130_fd_sc_hd__fa_2_450/A sky130_fd_sc_hd__nor2b_1_24/A sky130_fd_sc_hd__nand2_1_722/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_132 sky130_fd_sc_hd__xnor2_1_283/Y sky130_fd_sc_hd__xnor2_1_280/Y
+ sky130_fd_sc_hd__fa_2_456/A sky130_fd_sc_hd__nor2b_1_19/A sky130_fd_sc_hd__o22ai_1_66/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_207 sky130_fd_sc_hd__nand2_1_207/Y sky130_fd_sc_hd__nor2_1_62/A
+ sky130_fd_sc_hd__nor2_1_62/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_806 sky130_fd_sc_hd__clkinv_1_806/Y sky130_fd_sc_hd__nand2_1_791/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_2_10 sky130_fd_sc_hd__nor2_2_10/B sky130_fd_sc_hd__nor2_2_10/Y
+ sky130_fd_sc_hd__buf_6_4/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__nand2_1_218 sky130_fd_sc_hd__nand2_1_218/Y sky130_fd_sc_hd__nor2_1_65/A
+ sky130_fd_sc_hd__nor2_1_65/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_817 sky130_fd_sc_hd__nand2_1_812/A sky130_fd_sc_hd__nor2_1_259/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_2_21 sky130_fd_sc_hd__nor2_2_21/B sky130_fd_sc_hd__nor2_2_21/Y
+ sky130_fd_sc_hd__nor2_2_21/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__nand2_1_229 sky130_fd_sc_hd__nand2_1_229/Y sky130_fd_sc_hd__nand2_1_239/Y
+ sky130_fd_sc_hd__nand2_1_235/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_828 sky130_fd_sc_hd__clkinv_1_828/Y sky130_fd_sc_hd__nand2_1_835/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_2_32 sky130_fd_sc_hd__nor2_2_32/B sky130_fd_sc_hd__nor2_2_32/Y
+ sky130_fd_sc_hd__nor2_2_32/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__clkinv_1_839 sky130_fd_sc_hd__buf_8_88/A sky130_fd_sc_hd__clkinv_1_839/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o211ai_1_0 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_0/A2
+ sky130_fd_sc_hd__o211ai_1_0/Y sky130_fd_sc_hd__a22oi_1_32/Y sky130_fd_sc_hd__a22oi_1_33/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__conb_1_17 sky130_fd_sc_hd__conb_1_17/LO sky130_fd_sc_hd__conb_1_17/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_28 sky130_fd_sc_hd__conb_1_28/LO sky130_fd_sc_hd__conb_1_28/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_39 sky130_fd_sc_hd__conb_1_39/LO sky130_fd_sc_hd__conb_1_39/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__o21ai_1_370 vssd1 vccd1 sky130_fd_sc_hd__buf_2_1/X sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__o21ai_1_370/B1 sky130_fd_sc_hd__xor2_1_184/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_381 vssd1 vccd1 sky130_fd_sc_hd__inv_2_26/Y sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__nand2_1_160/Y sky130_fd_sc_hd__xor2_1_196/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_392 vssd1 vccd1 sky130_fd_sc_hd__buf_2_2/X sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__o21ai_1_392/B1 sky130_fd_sc_hd__xor2_1_208/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_802 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_813 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_824 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_835 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_846 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_730 sky130_fd_sc_hd__xnor2_1_206/A sky130_fd_sc_hd__nand2_1_731/Y
+ sky130_fd_sc_hd__or2_0_86/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_857 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_741 sky130_fd_sc_hd__xnor2_1_209/A sky130_fd_sc_hd__nand2_1_742/Y
+ sky130_fd_sc_hd__or2_0_88/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_868 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_752 sky130_fd_sc_hd__nand2_1_752/Y sky130_fd_sc_hd__nor2_1_241/A
+ sky130_fd_sc_hd__a22o_1_8/A2 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_879 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__mux2_2_50 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_50/A1 sky130_fd_sc_hd__buf_4_13/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__xnor2_2_4/A vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_763 sky130_fd_sc_hd__xnor2_1_216/A sky130_fd_sc_hd__nand2_1_780/Y
+ sky130_fd_sc_hd__nand2_1_763/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_774 sky130_fd_sc_hd__nand2_1_774/Y sky130_fd_sc_hd__or2_1_12/X
+ sky130_fd_sc_hd__nor2_1_242/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_785 sky130_fd_sc_hd__nand2_1_785/Y sky130_fd_sc_hd__or2_0_97/A
+ sky130_fd_sc_hd__or2_0_97/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_796 sky130_fd_sc_hd__xor2_1_677/B sky130_fd_sc_hd__nand2_1_797/Y
+ sky130_fd_sc_hd__nand2_1_796/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_1801 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1812 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1823 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1834 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1845 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1856 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1867 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__or2b_2_0 sky130_fd_sc_hd__or2b_2_0/A sky130_fd_sc_hd__nor2_4_8/B
+ sky130_fd_sc_hd__or2b_2_0/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__or2b_2
Xsky130_fd_sc_hd__a222oi_1_250 vccd1 vssd1 sky130_fd_sc_hd__and3_4_17/X sky130_fd_sc_hd__and2_0_45/A
+ sky130_fd_sc_hd__and2_0_87/A sky130_fd_sc_hd__nor2_2_20/Y sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__o21ai_1_449/B1 sky130_fd_sc_hd__nor2b_2_4/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_190 vssd1 vccd1 sky130_fd_sc_hd__buf_12_34/A sky130_fd_sc_hd__clkbuf_1_60/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_261 vccd1 vssd1 sky130_fd_sc_hd__and3_4_15/X sky130_fd_sc_hd__buf_2_23/X
+ sky130_fd_sc_hd__buf_2_31/X sky130_fd_sc_hd__nor2_1_130/Y sky130_fd_sc_hd__buf_2_19/X
+ sky130_fd_sc_hd__o21ai_1_463/B1 sky130_fd_sc_hd__nor2b_1_11/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_272 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__or2_0_60/B
+ sky130_fd_sc_hd__or2_0_60/A sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__or2_0_61/A
+ sky130_fd_sc_hd__o21ai_1_476/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_420 sky130_fd_sc_hd__or2_1_12/A sky130_fd_sc_hd__nor2_1_243/B
+ sky130_fd_sc_hd__fa_2_420/A sky130_fd_sc_hd__fa_2_420/B sky130_fd_sc_hd__fa_2_421/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_283 vccd1 vssd1 sky130_fd_sc_hd__and3_4_17/X sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__buf_6_1/X sky130_fd_sc_hd__nor2_2_20/Y sky130_fd_sc_hd__and2_0_38/A
+ sky130_fd_sc_hd__o21ai_1_491/B1 sky130_fd_sc_hd__nor2b_2_4/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_431 sky130_fd_sc_hd__fa_2_428/CIN sky130_fd_sc_hd__fa_2_433/CIN
+ sky130_fd_sc_hd__fa_2_431/A sky130_fd_sc_hd__fa_2_431/B sky130_fd_sc_hd__o22ai_1_69/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_294 vccd1 vssd1 sky130_fd_sc_hd__and3_4_15/X sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__buf_6_2/X sky130_fd_sc_hd__nor2_1_130/Y sky130_fd_sc_hd__buf_4_7/X
+ sky130_fd_sc_hd__o21ai_1_504/B1 sky130_fd_sc_hd__nor2b_1_11/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_442 sky130_fd_sc_hd__fa_2_438/B sky130_fd_sc_hd__fa_2_442/SUM
+ sky130_fd_sc_hd__fa_2_442/A sky130_fd_sc_hd__fa_2_442/B sky130_fd_sc_hd__o22ai_1_91/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_453 sky130_fd_sc_hd__fa_2_453/COUT sky130_fd_sc_hd__fa_2_453/SUM
+ sky130_fd_sc_hd__fa_2_453/A sky130_fd_sc_hd__fa_2_453/B sky130_fd_sc_hd__fa_2_453/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_464 sky130_fd_sc_hd__fa_2_462/CIN sky130_fd_sc_hd__fa_2_464/SUM
+ sky130_fd_sc_hd__fa_2_464/A sky130_fd_sc_hd__fa_2_464/B sky130_fd_sc_hd__fa_2_464/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_475 sky130_fd_sc_hd__or2_0_102/B sky130_fd_sc_hd__nor2_1_257/A
+ sky130_fd_sc_hd__fa_2_475/A sky130_fd_sc_hd__fa_2_475/B sky130_fd_sc_hd__nor2b_1_49/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_486 sky130_fd_sc_hd__nor2_1_262/B sky130_fd_sc_hd__or2_0_108/A
+ sky130_fd_sc_hd__fa_2_486/A sky130_fd_sc_hd__fa_2_486/B sky130_fd_sc_hd__nor2b_1_71/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__decap_8_14 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__nor2_1_207 sky130_fd_sc_hd__buf_2_15/X sky130_fd_sc_hd__nor2_1_207/Y
+ sky130_fd_sc_hd__buf_2_4/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_218 sky130_fd_sc_hd__or2_0_71/B sky130_fd_sc_hd__nor2_1_218/Y
+ sky130_fd_sc_hd__buf_2_29/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_229 sky130_fd_sc_hd__mux2_2_48/X sky130_fd_sc_hd__nor2_1_229/Y
+ sky130_fd_sc_hd__mux2_4_2/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_403 sky130_fd_sc_hd__buf_12_76/X sky130_fd_sc_hd__buf_12_636/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_414 sky130_fd_sc_hd__buf_12_89/X sky130_fd_sc_hd__buf_12_496/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_425 sky130_fd_sc_hd__buf_12_425/A sky130_fd_sc_hd__buf_12_651/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_436 sky130_fd_sc_hd__buf_12_436/A sky130_fd_sc_hd__buf_12_574/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_447 sky130_fd_sc_hd__buf_12_447/A sky130_fd_sc_hd__buf_12_661/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_458 sky130_fd_sc_hd__buf_12_458/A sky130_fd_sc_hd__buf_12_625/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_469 sky130_fd_sc_hd__buf_12_469/A sky130_fd_sc_hd__buf_12_518/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_109 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_603 sky130_fd_sc_hd__clkinv_1_603/Y sky130_fd_sc_hd__nand2_1_642/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_614 sky130_fd_sc_hd__or2b_2_2/A sky130_fd_sc_hd__dfxtp_1_191/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_625 sky130_fd_sc_hd__clkinv_1_625/Y sky130_fd_sc_hd__nand2_1_663/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_636 sky130_fd_sc_hd__nand2_1_684/A sky130_fd_sc_hd__nor2_1_226/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_647 sky130_fd_sc_hd__clkinv_1_647/Y sky130_fd_sc_hd__nand2_1_707/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_658 sky130_fd_sc_hd__o22ai_1_133/B1 sky130_fd_sc_hd__or2_0_77/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_669 sky130_fd_sc_hd__clkinv_1_669/Y sky130_fd_sc_hd__nand2_1_740/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1108 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1119 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_12 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_353/Q sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__o211ai_1_28/Y sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__a222oi_1_12/Y sky130_fd_sc_hd__dfxtp_1_304/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_23 vccd1 vssd1 sky130_fd_sc_hd__xor2_1_419/X sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__xor2_1_632/X sky130_fd_sc_hd__xor2_1_207/X sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_23/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_610 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_34 vccd1 vssd1 sky130_fd_sc_hd__xor2_1_359/X sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__xor2_1_572/X sky130_fd_sc_hd__xor2_1_146/X sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_34/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_621 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_45 vccd1 vssd1 sky130_fd_sc_hd__xor2_1_234/X sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__inv_2_58/A sky130_fd_sc_hd__xor2_1_21/X sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_45/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_632 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_56 vccd1 vssd1 sky130_fd_sc_hd__and3_4_2/X sky130_fd_sc_hd__or2_0_60/B
+ sky130_fd_sc_hd__or2_0_60/A sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__or2_0_61/A
+ sky130_fd_sc_hd__a222oi_1_56/Y sky130_fd_sc_hd__and2b_4_4/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_643 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_67 vccd1 vssd1 sky130_fd_sc_hd__and3_1_0/X sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__buf_2_32/X sky130_fd_sc_hd__nor2_1_56/Y sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__a222oi_1_67/Y sky130_fd_sc_hd__nor2b_1_3/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_654 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_78 vccd1 vssd1 sky130_fd_sc_hd__and3_4_7/X sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__nor2_1_85/B sky130_fd_sc_hd__nor2_2_7/Y sky130_fd_sc_hd__nor2_2_10/B
+ sky130_fd_sc_hd__a222oi_1_78/Y sky130_fd_sc_hd__nor2b_2_1/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__xnor2_1_14 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_14/B sky130_fd_sc_hd__and3_1_0/C
+ sky130_fd_sc_hd__fa_2_56/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_25 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_104/A sky130_fd_sc_hd__and3_4_5/B
+ sky130_fd_sc_hd__xnor2_1_27/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_665 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_89 vccd1 vssd1 sky130_fd_sc_hd__and3_4_2/X sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__buf_4_4/X sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__a222oi_1_89/Y sky130_fd_sc_hd__and2b_4_4/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_676 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_36 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_149/A sky130_fd_sc_hd__and3_4_7/B
+ sky130_fd_sc_hd__xnor2_1_38/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_560 sky130_fd_sc_hd__xor2_1_526/B sky130_fd_sc_hd__nand2_1_561/Y
+ sky130_fd_sc_hd__nand2_1_560/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_687 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_47 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_47/B sky130_fd_sc_hd__inv_2_9/A
+ sky130_fd_sc_hd__xnor2_1_47/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_571 sky130_fd_sc_hd__o21ai_2_14/B1 sky130_fd_sc_hd__nor2_2_25/A
+ sky130_fd_sc_hd__nor2_2_25/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_698 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_58 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_58/B sky130_fd_sc_hd__inv_2_15/A
+ sky130_fd_sc_hd__xnor2_1_58/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_582 sky130_fd_sc_hd__nand2_1_582/Y sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__nor2_1_73/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_69 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_69/B sky130_fd_sc_hd__xnor2_1_69/Y
+ sky130_fd_sc_hd__xnor2_1_69/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_593 sky130_fd_sc_hd__nand2_1_593/Y sky130_fd_sc_hd__nand2_1_606/Y
+ sky130_fd_sc_hd__nand2_1_601/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_1140 sky130_fd_sc_hd__buf_4_39/A sky130_fd_sc_hd__buf_4_42/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1151 sky130_fd_sc_hd__buf_2_48/A sky130_fd_sc_hd__inv_4_21/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_2_3 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_3/Y sky130_fd_sc_hd__inv_2_52/Y
+ sky130_fd_sc_hd__xnor2_2_3/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_2
Xsky130_fd_sc_hd__decap_12_1620 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1631 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1642 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1653 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1664 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1675 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1686 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1697 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__or4_1_0 sky130_fd_sc_hd__ha_2_7/A sky130_fd_sc_hd__ha_2_4/A sky130_fd_sc_hd__or4_1_0/X
+ sky130_fd_sc_hd__or4_1_1/C sky130_fd_sc_hd__ha_2_5/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__or4_1
Xsky130_fd_sc_hd__fa_2_250 sky130_fd_sc_hd__fa_2_246/CIN sky130_fd_sc_hd__fa_2_252/A
+ sky130_fd_sc_hd__fa_2_250/A sky130_fd_sc_hd__fa_2_250/B sky130_fd_sc_hd__xor2_1_361/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_261 sky130_fd_sc_hd__fa_2_259/B sky130_fd_sc_hd__fa_2_263/CIN
+ sky130_fd_sc_hd__fa_2_261/A sky130_fd_sc_hd__fa_2_261/B sky130_fd_sc_hd__xor2_1_378/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_272 sky130_fd_sc_hd__nor2_1_149/A sky130_fd_sc_hd__nor2_1_152/B
+ sky130_fd_sc_hd__fa_2_272/A sky130_fd_sc_hd__fa_2_272/B sky130_fd_sc_hd__fa_2_272/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_283 sky130_fd_sc_hd__xor3_1_21/C sky130_fd_sc_hd__fa_2_287/CIN
+ sky130_fd_sc_hd__fa_2_283/A sky130_fd_sc_hd__fa_2_283/B sky130_fd_sc_hd__fa_2_290/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_294 sky130_fd_sc_hd__fa_2_288/CIN sky130_fd_sc_hd__fa_2_291/B
+ sky130_fd_sc_hd__fa_2_294/A sky130_fd_sc_hd__fa_2_294/B sky130_fd_sc_hd__xor2_1_449/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22oi_1_5 sky130_fd_sc_hd__nor2_4_0/Y sky130_fd_sc_hd__nor2_2_0/Y
+ sky130_fd_sc_hd__a22oi_1_5/B2 sky130_fd_sc_hd__or2_0_87/A sky130_fd_sc_hd__nand2_2_1/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_200 sky130_fd_sc_hd__buf_6_61/X sky130_fd_sc_hd__buf_12_200/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_211 sky130_fd_sc_hd__buf_6_32/X sky130_fd_sc_hd__buf_12_387/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_222 sky130_fd_sc_hd__buf_6_75/X sky130_fd_sc_hd__buf_12_430/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_233 sky130_fd_sc_hd__buf_6_41/X sky130_fd_sc_hd__buf_12_404/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_80 sky130_fd_sc_hd__a21oi_1_80/A1 sky130_fd_sc_hd__nor2_1_119/A
+ sky130_fd_sc_hd__a21oi_1_80/Y sky130_fd_sc_hd__or2_0_41/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_244 sky130_fd_sc_hd__buf_6_79/X sky130_fd_sc_hd__buf_12_441/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_91 sky130_fd_sc_hd__o21ai_1_595/Y sky130_fd_sc_hd__o21ai_1_576/Y
+ sky130_fd_sc_hd__a21oi_1_91/Y sky130_fd_sc_hd__nor2_1_141/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_1_103 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_190/Q sky130_fd_sc_hd__dfxtp_1_158/Q sky130_fd_sc_hd__o21ai_1_9/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_255 sky130_fd_sc_hd__buf_12_74/X sky130_fd_sc_hd__buf_12_392/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_114 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_172/Q sky130_fd_sc_hd__dfxtp_1_140/Q sky130_fd_sc_hd__o21ai_1_20/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_266 sky130_fd_sc_hd__buf_6_73/X sky130_fd_sc_hd__buf_12_266/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_125 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_159/Q sky130_fd_sc_hd__dfxtp_1_127/Q sky130_fd_sc_hd__o21ai_1_31/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_277 sky130_fd_sc_hd__buf_12_3/X sky130_fd_sc_hd__buf_12_624/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_136 sky130_fd_sc_hd__xor2_1_255/X sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xor2_1_42/X sky130_fd_sc_hd__o21ai_1_52/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_288 sky130_fd_sc_hd__buf_12_4/X sky130_fd_sc_hd__buf_12_672/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_147 sky130_fd_sc_hd__xnor2_1_86/Y sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xnor2_1_23/Y sky130_fd_sc_hd__o21ai_1_73/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_299 sky130_fd_sc_hd__buf_12_64/X sky130_fd_sc_hd__buf_12_555/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_158 sky130_fd_sc_hd__xor2_1_359/X sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xor2_1_146/X sky130_fd_sc_hd__o21ai_1_98/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_400 sky130_fd_sc_hd__nand2_1_306/A sky130_fd_sc_hd__nor2_1_102/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22oi_1_169 sky130_fd_sc_hd__xor2_1_384/X sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xor2_1_171/X sky130_fd_sc_hd__a22oi_1_169/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_411 sky130_fd_sc_hd__nand2_1_462/A sky130_fd_sc_hd__nor2_2_17/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_422 sky130_fd_sc_hd__o21ai_1_434/A2 sky130_fd_sc_hd__xnor2_1_72/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_433 sky130_fd_sc_hd__nand2_1_359/A sky130_fd_sc_hd__nor2_1_116/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_444 sky130_fd_sc_hd__nor2_1_119/A sky130_fd_sc_hd__nand2_1_382/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_455 sky130_fd_sc_hd__nor2_1_125/B sky130_fd_sc_hd__nand2_1_397/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_466 sky130_fd_sc_hd__a21oi_2_12/B1 sky130_fd_sc_hd__nand2_1_415/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_477 sky130_fd_sc_hd__xnor2_1_104/B sky130_fd_sc_hd__a21oi_1_91/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_488 sky130_fd_sc_hd__nand2_1_446/A sky130_fd_sc_hd__nor2_1_149/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_499 sky130_fd_sc_hd__xnor2_1_119/B sky130_fd_sc_hd__a21oi_1_100/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a222oi_1_0 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_341/Q sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__o211ai_1_16/Y sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__a222oi_1_0/Y sky130_fd_sc_hd__dfxtp_1_292/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_440 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_451 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_462 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_473 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_484 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_495 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_207 sky130_fd_sc_hd__o21a_1_1/X sky130_fd_sc_hd__xor2_1_207/X
+ sky130_fd_sc_hd__xor2_1_207/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_390 sky130_fd_sc_hd__nor2_1_126/A sky130_fd_sc_hd__or2_0_44/X
+ sky130_fd_sc_hd__or2_0_45/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_218 sky130_fd_sc_hd__fa_2_217/A sky130_fd_sc_hd__xor3_1_18/C
+ sky130_fd_sc_hd__xor2_1_218/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_229 sky130_fd_sc_hd__xor2_1_383/B sky130_fd_sc_hd__fa_2_144/B
+ sky130_fd_sc_hd__xor2_1_229/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1450 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1461 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1472 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_903 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_686/A sky130_fd_sc_hd__nor2_1_264/Y
+ sky130_fd_sc_hd__nand2_1_833/Y sky130_fd_sc_hd__xnor2_1_300/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1483 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_914 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_914/A2 sky130_fd_sc_hd__nor2_1_274/Y
+ sky130_fd_sc_hd__nor3_1_2/Y sky130_fd_sc_hd__nor2_1_268/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1494 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_925 vssd1 vccd1 sky130_fd_sc_hd__nand2_1_866/B sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a21o_2_3/A2 sky130_fd_sc_hd__o21ai_1_925/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_8_7 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__buf_2_12 vccd1 vssd1 sky130_fd_sc_hd__buf_2_12/X sky130_fd_sc_hd__buf_2_12/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_23 vccd1 vssd1 sky130_fd_sc_hd__buf_2_23/X sky130_fd_sc_hd__buf_2_27/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_34 vccd1 vssd1 sky130_fd_sc_hd__buf_8_89/A la_data_out[42]
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_45 vccd1 vssd1 sky130_fd_sc_hd__buf_2_45/X sky130_fd_sc_hd__buf_2_45/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_56 vccd1 vssd1 sky130_fd_sc_hd__buf_8_92/A sky130_fd_sc_hd__buf_8_7/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_67 vccd1 vssd1 sky130_fd_sc_hd__buf_2_68/A sky130_fd_sc_hd__buf_2_67/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_78 vccd1 vssd1 sky130_fd_sc_hd__buf_2_78/X sky130_fd_sc_hd__buf_2_78/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_89 vccd1 vssd1 sky130_fd_sc_hd__buf_2_89/X sky130_fd_sc_hd__buf_2_89/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o211ai_1_50 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o22ai_1_13/B1
+ sky130_fd_sc_hd__fah_1_13/A sky130_fd_sc_hd__nand2_1_70/Y sky130_fd_sc_hd__a21oi_1_21/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_61 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o22ai_1_0/B1
+ sky130_fd_sc_hd__or2_0_70/B sky130_fd_sc_hd__nand2_1_81/Y sky130_fd_sc_hd__a21oi_1_32/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__diode_2_7 sky130_fd_sc_hd__conb_1_147/HI vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__and2_0_209 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_52/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_75/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__xor3_1_18 sky130_fd_sc_hd__xor3_1_18/X sky130_fd_sc_hd__xor3_1_18/C
+ sky130_fd_sc_hd__xor3_1_18/B sky130_fd_sc_hd__xor3_1_18/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__xor3_1_29 sky130_fd_sc_hd__xor3_1_29/X sky130_fd_sc_hd__xor3_1_29/C
+ sky130_fd_sc_hd__xor3_1_29/B sky130_fd_sc_hd__xor3_1_29/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__clkinv_1_230 sky130_fd_sc_hd__nor2_1_9/A sky130_fd_sc_hd__dfxtp_1_132/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_241 sky130_fd_sc_hd__o22ai_1_1/A2 sky130_fd_sc_hd__dfxtp_1_160/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_252 sky130_fd_sc_hd__o21ai_1_98/A2 sky130_fd_sc_hd__xor2_1_572/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_263 sky130_fd_sc_hd__o21ai_1_141/A2 sky130_fd_sc_hd__xor2_1_624/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_274 sky130_fd_sc_hd__and2_0_141/A sky130_fd_sc_hd__a222oi_1_18/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_285 sky130_fd_sc_hd__and2_0_206/A sky130_fd_sc_hd__a222oi_1_29/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_296 sky130_fd_sc_hd__and2_0_241/A sky130_fd_sc_hd__a222oi_1_40/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xor3_1_3 sky130_fd_sc_hd__xor3_1_3/X sky130_fd_sc_hd__xor3_1_3/C
+ sky130_fd_sc_hd__xor3_1_4/X sky130_fd_sc_hd__xor3_1_3/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__a21oi_1_4 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_33/Y
+ sky130_fd_sc_hd__a21oi_1_4/Y sky130_fd_sc_hd__dfxtp_1_91/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__and3_4_10 sky130_fd_sc_hd__nor2_4_12/B sky130_fd_sc_hd__nor2_4_12/A
+ sky130_fd_sc_hd__and3_4_10/C sky130_fd_sc_hd__and3_4_10/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__clkbuf_4_17 sky130_fd_sc_hd__a22o_1_48/A2 sky130_fd_sc_hd__clkbuf_4_17/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and3_4_21 sky130_fd_sc_hd__nor2_4_17/B sky130_fd_sc_hd__nor2_4_17/A
+ sky130_fd_sc_hd__and3_4_21/C sky130_fd_sc_hd__and3_4_21/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__clkbuf_4_28 sky130_fd_sc_hd__buf_4_29/A sky130_fd_sc_hd__clkbuf_4_28/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_39 la_data_out[62] sky130_fd_sc_hd__dfxtp_1_477/Q vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__a21oi_1_160 sky130_fd_sc_hd__xnor2_1_213/B sky130_fd_sc_hd__o21ai_1_885/Y
+ sky130_fd_sc_hd__xor2_1_660/A sky130_fd_sc_hd__nor2_1_242/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_171 sky130_fd_sc_hd__xnor2_1_292/B sky130_fd_sc_hd__clkinv_1_810/Y
+ sky130_fd_sc_hd__xor2_1_677/A sky130_fd_sc_hd__or2_0_101/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_182 sky130_fd_sc_hd__or2_0_112/X sky130_fd_sc_hd__clkinv_1_831/Y
+ sky130_fd_sc_hd__xor2_1_688/B sky130_fd_sc_hd__nor2b_1_85/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_193 la_data_out[45] sky130_fd_sc_hd__o21ai_1_918/Y sky130_fd_sc_hd__a21o_2_0/A2
+ sky130_fd_sc_hd__o21ai_1_918/A2 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_101 sky130_fd_sc_hd__buf_8_101/A sky130_fd_sc_hd__buf_6_83/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_112 sky130_fd_sc_hd__buf_8_112/A sky130_fd_sc_hd__buf_6_55/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_123 sky130_fd_sc_hd__buf_8_123/A sky130_fd_sc_hd__buf_6_68/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_134 sky130_fd_sc_hd__buf_8_134/A sky130_fd_sc_hd__buf_8_134/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_145 sky130_fd_sc_hd__buf_8_145/A sky130_fd_sc_hd__buf_8_145/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nor2_4_7 sky130_fd_sc_hd__nor2_4_7/Y sky130_fd_sc_hd__nor2_4_7/A
+ sky130_fd_sc_hd__nor2_4_7/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__buf_8_156 sky130_fd_sc_hd__buf_8_156/A sky130_fd_sc_hd__buf_8_156/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__decap_12_270 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_281 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_292 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_700 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_3/Y sky130_fd_sc_hd__nand2b_1_21/Y
+ sky130_fd_sc_hd__o21ai_1_700/B1 sky130_fd_sc_hd__xor2_1_479/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1280 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_711 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_176/Y sky130_fd_sc_hd__nor2_1_177/Y
+ sky130_fd_sc_hd__nand2_1_543/Y sky130_fd_sc_hd__o21ai_1_711/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1291 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_722 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_751/A2 sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_722/B1 sky130_fd_sc_hd__xor2_1_499/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_733 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_733/A2 sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_733/B1 sky130_fd_sc_hd__xor2_1_511/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_744 vssd1 vccd1 sky130_fd_sc_hd__buf_2_12/X sky130_fd_sc_hd__nand2b_1_15/Y
+ sky130_fd_sc_hd__o21ai_1_744/B1 sky130_fd_sc_hd__xor2_1_519/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_755 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_861/A2 sky130_fd_sc_hd__nand2b_1_20/Y
+ sky130_fd_sc_hd__nand2_1_495/Y sky130_fd_sc_hd__xor2_1_529/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_766 vssd1 vccd1 sky130_fd_sc_hd__inv_2_48/Y sky130_fd_sc_hd__nand2b_1_15/Y
+ sky130_fd_sc_hd__o21ai_1_766/B1 sky130_fd_sc_hd__xor2_1_541/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_777 vssd1 vccd1 sky130_fd_sc_hd__inv_2_45/Y sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__o21ai_1_777/B1 sky130_fd_sc_hd__xor2_1_551/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_788 vssd1 vccd1 sky130_fd_sc_hd__inv_2_43/Y sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__o21ai_1_788/B1 sky130_fd_sc_hd__xor2_1_562/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_799 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_799/A2 sky130_fd_sc_hd__nor2_1_193/Y
+ sky130_fd_sc_hd__nand2_1_596/Y sky130_fd_sc_hd__o21ai_1_799/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_40 sky130_fd_sc_hd__xor2_1_6/B sky130_fd_sc_hd__xor2_1_40/X
+ sky130_fd_sc_hd__xor2_1_40/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_51 sky130_fd_sc_hd__xor2_1_9/B sky130_fd_sc_hd__xor2_1_51/X
+ sky130_fd_sc_hd__xor2_1_51/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_62 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__fa_2_36/B
+ sky130_fd_sc_hd__xor2_1_62/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_18 sky130_fd_sc_hd__inv_2_77/Y sky130_fd_sc_hd__buf_12_18/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_73 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__fa_2_54/B
+ sky130_fd_sc_hd__xor2_1_73/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_29 sky130_fd_sc_hd__buf_12_29/A sky130_fd_sc_hd__buf_12_29/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_84 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__xor2_1_84/X
+ sky130_fd_sc_hd__xor2_1_84/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_95 sky130_fd_sc_hd__fa_2_75/A sky130_fd_sc_hd__fa_2_72/B
+ sky130_fd_sc_hd__xor2_1_95/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2b_1_1 sky130_fd_sc_hd__nand2b_1_1/Y sky130_fd_sc_hd__nor2_2_8/A
+ sky130_fd_sc_hd__nor2_2_8/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__o21ai_2_16 sky130_fd_sc_hd__o21ai_2_16/B1 sky130_fd_sc_hd__o21ai_2_16/Y
+ sky130_fd_sc_hd__o21ai_2_16/A2 sky130_fd_sc_hd__o21ai_2_16/A1 vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__o21ai_2
Xsky130_fd_sc_hd__xor2_1_560 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__xor2_1_560/X
+ sky130_fd_sc_hd__xor2_1_560/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_571 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__fa_2_386/B
+ sky130_fd_sc_hd__xor2_1_571/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_582 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__fa_2_394/A
+ sky130_fd_sc_hd__xor2_1_582/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_593 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__fa_2_399/A
+ sky130_fd_sc_hd__xor2_1_593/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a222oi_1_602 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_420/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_452/Q sky130_fd_sc_hd__nor2_4_19/B
+ sky130_fd_sc_hd__clkinv_1_799/A sky130_fd_sc_hd__dfxtp_1_388/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__maj3_1_3 sky130_fd_sc_hd__maj3_1_3/C sky130_fd_sc_hd__maj3_1_3/X
+ sky130_fd_sc_hd__maj3_1_3/B sky130_fd_sc_hd__maj3_1_3/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__and2_0_12 vccd1 vssd1 sky130_fd_sc_hd__and2_0_12/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_12/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_23 vccd1 vssd1 sky130_fd_sc_hd__and2_0_23/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__nor2_2_5/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_34 vccd1 vssd1 sky130_fd_sc_hd__and2_0_34/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__or2_0_53/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_45 vccd1 vssd1 sky130_fd_sc_hd__and2_0_45/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__and2_0_45/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_56 vccd1 vssd1 sky130_fd_sc_hd__and2_0_56/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__buf_2_19/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_67 vccd1 vssd1 sky130_fd_sc_hd__and2_0_67/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__or2_0_60/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_78 vccd1 vssd1 sky130_fd_sc_hd__and2_0_78/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__buf_6_0/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nor2_2_4 sky130_fd_sc_hd__nor2_2_4/B sky130_fd_sc_hd__nor2_2_4/Y
+ sky130_fd_sc_hd__nor2_2_5/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__and2_0_89 vccd1 vssd1 sky130_fd_sc_hd__and2_0_89/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__or2_0_9/B vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_8_11 sky130_fd_sc_hd__inv_2_74/Y sky130_fd_sc_hd__buf_8_11/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_22 sky130_fd_sc_hd__buf_8_22/A sky130_fd_sc_hd__buf_8_22/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_33 sky130_fd_sc_hd__buf_8_33/A sky130_fd_sc_hd__buf_8_33/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_44 sky130_fd_sc_hd__buf_8_44/A sky130_fd_sc_hd__buf_8_44/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_55 sky130_fd_sc_hd__buf_8_55/A sky130_fd_sc_hd__buf_8_55/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_66 sky130_fd_sc_hd__buf_8_66/A sky130_fd_sc_hd__buf_8_66/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_77 la_data_out[41] sky130_fd_sc_hd__buf_8_77/X vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xnor2_1_190 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_190/B sky130_fd_sc_hd__and2_0_273/A
+ sky130_fd_sc_hd__xnor2_1_190/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__buf_8_88 sky130_fd_sc_hd__buf_8_88/A sky130_fd_sc_hd__buf_8_88/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_207 sky130_fd_sc_hd__xnor2_1_153/A sky130_fd_sc_hd__dfxtp_2_0/CLK
+ sky130_fd_sc_hd__and2_0_80/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_8_99 sky130_fd_sc_hd__buf_8_99/A sky130_fd_sc_hd__buf_8_99/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_218 sky130_fd_sc_hd__dfxtp_1_218/Q sky130_fd_sc_hd__dfxtp_2_5/CLK
+ sky130_fd_sc_hd__and2_0_11/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_229 sky130_fd_sc_hd__xor2_1_383/B sky130_fd_sc_hd__dfxtp_1_230/CLK
+ sky130_fd_sc_hd__and2_0_45/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_530 vssd1 vccd1 sky130_fd_sc_hd__inv_2_37/Y sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_530/B1 sky130_fd_sc_hd__xor2_1_329/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_541 vssd1 vccd1 sky130_fd_sc_hd__buf_2_11/X sky130_fd_sc_hd__nand2b_1_9/Y
+ sky130_fd_sc_hd__o21ai_1_541/B1 sky130_fd_sc_hd__xor2_1_339/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_552 vssd1 vccd1 sky130_fd_sc_hd__inv_2_38/Y sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_552/B1 sky130_fd_sc_hd__xor2_1_350/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_563 vssd1 vccd1 sky130_fd_sc_hd__buf_2_10/X sky130_fd_sc_hd__nand2b_1_9/Y
+ sky130_fd_sc_hd__o21ai_1_563/B1 sky130_fd_sc_hd__xor2_1_360/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_574 vssd1 vccd1 sky130_fd_sc_hd__buf_2_7/X sky130_fd_sc_hd__nand2b_1_9/Y
+ sky130_fd_sc_hd__o21ai_1_574/B1 sky130_fd_sc_hd__xor2_1_371/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_585 vssd1 vccd1 sky130_fd_sc_hd__inv_2_42/Y sky130_fd_sc_hd__nand2_1_438/Y
+ sky130_fd_sc_hd__a21oi_1_93/Y sky130_fd_sc_hd__xnor2_1_108/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_596 vssd1 vccd1 sky130_fd_sc_hd__buf_2_8/X sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_596/B1 sky130_fd_sc_hd__xor2_1_390/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__buf_2_107 vccd1 vssd1 sky130_fd_sc_hd__buf_2_107/X sky130_fd_sc_hd__buf_2_107/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_118 vccd1 vssd1 sky130_fd_sc_hd__buf_2_118/X sky130_fd_sc_hd__buf_2_118/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_129 vccd1 vssd1 sky130_fd_sc_hd__buf_2_129/X sky130_fd_sc_hd__buf_2_129/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__xor2_1_390 sky130_fd_sc_hd__fa_2_281/A sky130_fd_sc_hd__xor2_1_390/X
+ sky130_fd_sc_hd__xor2_1_390/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__ha_2_7 vssd1 vccd1 sky130_fd_sc_hd__ha_2_7/A sky130_fd_sc_hd__ha_2_6/B
+ sky130_fd_sc_hd__nor3_1_0/A sky130_fd_sc_hd__ha_2_7/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__a222oi_1_410 vccd1 vssd1 sky130_fd_sc_hd__and3_4_21/X sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__buf_4_5/X sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__o21ai_1_678/B1 sky130_fd_sc_hd__and2b_4_12/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_350 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2_2/A sky130_fd_sc_hd__a222oi_1_6/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_421 vccd1 vssd1 sky130_fd_sc_hd__and3_4_20/X sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__nor2_1_73/B sky130_fd_sc_hd__nor2_4_16/Y sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__o21ai_1_694/B1 sky130_fd_sc_hd__and2b_4_11/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_432 vccd1 vssd1 sky130_fd_sc_hd__and3_4_24/X sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__buf_6_2/X sky130_fd_sc_hd__nor2_1_183/Y sky130_fd_sc_hd__buf_4_7/X
+ sky130_fd_sc_hd__o21ai_1_706/B1 sky130_fd_sc_hd__nor2b_1_16/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_443 vccd1 vssd1 sky130_fd_sc_hd__and3_4_20/X sky130_fd_sc_hd__nor2_2_10/B
+ sky130_fd_sc_hd__buf_6_4/X sky130_fd_sc_hd__nor2_4_16/Y sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__o21ai_1_721/B1 sky130_fd_sc_hd__and2b_4_11/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_454 vccd1 vssd1 sky130_fd_sc_hd__and3_4_21/X sky130_fd_sc_hd__buf_6_4/X
+ sky130_fd_sc_hd__buf_6_0/X sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__o21ai_1_736/B1 sky130_fd_sc_hd__and2b_4_12/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_465 vccd1 vssd1 sky130_fd_sc_hd__and3_4_21/X sky130_fd_sc_hd__nor2_2_10/B
+ sky130_fd_sc_hd__buf_6_4/X sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__o21ai_1_749/B1 sky130_fd_sc_hd__and2b_4_12/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_476 vccd1 vssd1 sky130_fd_sc_hd__and3_4_20/X sky130_fd_sc_hd__buf_2_4/A
+ sky130_fd_sc_hd__buf_2_20/X sky130_fd_sc_hd__nor2_4_16/Y sky130_fd_sc_hd__buf_2_21/X
+ sky130_fd_sc_hd__o21ai_1_763/B1 sky130_fd_sc_hd__and2b_4_11/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_18 vssd1 vccd1 sky130_fd_sc_hd__nand2_1_123/A sky130_fd_sc_hd__xnor2_1_107/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_487 vccd1 vssd1 sky130_fd_sc_hd__and3_4_21/X sky130_fd_sc_hd__buf_2_20/X
+ sky130_fd_sc_hd__buf_2_21/X sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__o21ai_1_777/B1 sky130_fd_sc_hd__and2b_4_12/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_29 vssd1 vccd1 sky130_fd_sc_hd__and2_0_45/A sky130_fd_sc_hd__nor2_2_10/B
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_498 vccd1 vssd1 sky130_fd_sc_hd__and3_4_18/X sky130_fd_sc_hd__buf_2_29/X
+ sky130_fd_sc_hd__buf_2_30/X sky130_fd_sc_hd__nor2_2_32/Y sky130_fd_sc_hd__buf_2_26/X
+ sky130_fd_sc_hd__o21ai_1_791/B1 sky130_fd_sc_hd__nor2b_2_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__and2_0_370 vccd1 vssd1 sky130_fd_sc_hd__and2_0_370/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_63/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_381 vccd1 vssd1 sky130_fd_sc_hd__and2_0_381/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_79/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_392 vccd1 vssd1 sky130_fd_sc_hd__and2_0_392/X sky130_fd_sc_hd__and2_0_401/B
+ sky130_fd_sc_hd__and2_0_392/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__conb_1_1 sky130_fd_sc_hd__conb_1_1/LO sky130_fd_sc_hd__conb_1_1/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__buf_12_7 sky130_fd_sc_hd__buf_12_7/A sky130_fd_sc_hd__buf_12_7/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_607 sky130_fd_sc_hd__buf_12_607/A sky130_fd_sc_hd__buf_12_607/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_618 sky130_fd_sc_hd__buf_12_618/A sky130_fd_sc_hd__buf_12_618/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__inv_2_170 sky130_fd_sc_hd__inv_2_170/A sky130_fd_sc_hd__inv_2_170/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_12_629 sky130_fd_sc_hd__buf_12_629/A sky130_fd_sc_hd__buf_12_629/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__inv_2_181 sky130_fd_sc_hd__inv_2_181/A sky130_fd_sc_hd__inv_2_181/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_192 la_data_out[36] sky130_fd_sc_hd__nor2_2_1/B vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__o22ai_1_100 sky130_fd_sc_hd__xnor2_2_6/Y sky130_fd_sc_hd__xnor2_1_249/Y
+ sky130_fd_sc_hd__ha_2_15/A sky130_fd_sc_hd__xnor2_1_250/Y sky130_fd_sc_hd__o22ai_1_98/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_111 sky130_fd_sc_hd__xnor2_1_286/Y sky130_fd_sc_hd__xnor2_1_272/Y
+ sky130_fd_sc_hd__fa_2_452/A sky130_fd_sc_hd__nor2b_1_24/A sky130_fd_sc_hd__nand2_1_722/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_122 sky130_fd_sc_hd__xnor2_2_6/Y sky130_fd_sc_hd__xnor2_1_269/Y
+ sky130_fd_sc_hd__fa_2_455/CIN sky130_fd_sc_hd__xnor2_1_279/Y sky130_fd_sc_hd__o22ai_1_98/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_133 sky130_fd_sc_hd__nor2b_1_25/A sky130_fd_sc_hd__o22ai_1_133/B1
+ sky130_fd_sc_hd__ha_2_17/B sky130_fd_sc_hd__nand2b_1_29/Y sky130_fd_sc_hd__nand2_1_717/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_208 sky130_fd_sc_hd__or2_0_5/B sky130_fd_sc_hd__nor2_1_64/Y
+ sky130_fd_sc_hd__nor2_1_70/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_807 sky130_fd_sc_hd__nand2_1_792/A sky130_fd_sc_hd__nor2_1_254/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_2_11 sky130_fd_sc_hd__nor2_2_11/B sky130_fd_sc_hd__nor2_2_11/Y
+ sky130_fd_sc_hd__nor2_2_11/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__nand2_1_219 sky130_fd_sc_hd__nor2_1_67/A sky130_fd_sc_hd__or2_0_18/X
+ sky130_fd_sc_hd__or2_0_19/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_818 sky130_fd_sc_hd__clkinv_1_818/Y sky130_fd_sc_hd__nand2_1_815/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_2_22 sky130_fd_sc_hd__nor2_2_22/B sky130_fd_sc_hd__nor2_2_22/Y
+ sky130_fd_sc_hd__nor2_2_22/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__clkinv_1_829 sky130_fd_sc_hd__nand2_1_836/A sky130_fd_sc_hd__nor2_1_265/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o211ai_1_1 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_1/A2
+ sky130_fd_sc_hd__o211ai_1_1/Y sky130_fd_sc_hd__a22oi_1_34/Y sky130_fd_sc_hd__a22oi_1_35/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__conb_1_18 sky130_fd_sc_hd__conb_1_18/LO sky130_fd_sc_hd__conb_1_18/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_29 sky130_fd_sc_hd__conb_1_29/LO sky130_fd_sc_hd__conb_1_29/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__o21ai_1_360 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_176/A sky130_fd_sc_hd__nor2_1_91/Y
+ sky130_fd_sc_hd__nand2_1_276/Y sky130_fd_sc_hd__o21ai_1_360/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_371 vssd1 vccd1 sky130_fd_sc_hd__inv_2_19/Y sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__o21ai_1_371/B1 sky130_fd_sc_hd__xor2_1_185/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_382 vssd1 vccd1 sky130_fd_sc_hd__buf_2_1/X sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__o21ai_1_382/B1 sky130_fd_sc_hd__xor2_1_198/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_393 vssd1 vccd1 sky130_fd_sc_hd__nand2_4_4/Y sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__a22oi_1_200/Y sky130_fd_sc_hd__xor2_1_210/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_803 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_814 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_825 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_836 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_720 sky130_fd_sc_hd__o22ai_1_66/B2 sky130_fd_sc_hd__nor2b_1_19/A
+ sky130_fd_sc_hd__xor2_1_671/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_847 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_731 sky130_fd_sc_hd__nand2_1_731/Y sky130_fd_sc_hd__or2_0_86/A
+ sky130_fd_sc_hd__or2_0_86/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_858 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_742 sky130_fd_sc_hd__nand2_1_742/Y sky130_fd_sc_hd__or2_0_88/A
+ sky130_fd_sc_hd__or2_0_88/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_869 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__mux2_2_40 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_40/A1 sky130_fd_sc_hd__buf_2_87/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__fa_2_419/B vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_753 sky130_fd_sc_hd__xnor2_1_212/B sky130_fd_sc_hd__nand2_1_754/Y
+ sky130_fd_sc_hd__or2_0_95/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_51 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_51/A1 sky130_fd_sc_hd__buf_4_19/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__or2_0_80/A vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_764 sky130_fd_sc_hd__xor2_1_664/B sky130_fd_sc_hd__nand2_1_781/Y
+ sky130_fd_sc_hd__nand2_1_764/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_775 sky130_fd_sc_hd__nand2_1_775/Y sky130_fd_sc_hd__nor2_1_246/A
+ sky130_fd_sc_hd__nor2_1_246/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_786 sky130_fd_sc_hd__and2_0_302/B sky130_fd_sc_hd__or2_0_98/A
+ sky130_fd_sc_hd__or2_0_98/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_797 sky130_fd_sc_hd__nand2_1_797/Y sky130_fd_sc_hd__nor2_1_255/A
+ sky130_fd_sc_hd__nor2_1_255/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_1802 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1813 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1824 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1835 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1846 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1857 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1868 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__or2b_2_1 sky130_fd_sc_hd__or2b_2_1/A sky130_fd_sc_hd__and3_4_9/B
+ sky130_fd_sc_hd__or2b_2_1/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__or2b_2
Xsky130_fd_sc_hd__a222oi_1_240 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__or2_0_39/B
+ sky130_fd_sc_hd__or2_0_58/A sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__or2_0_9/B
+ sky130_fd_sc_hd__o21ai_1_434/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_180 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_46/A sky130_fd_sc_hd__xor2_1_697/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_251 vccd1 vssd1 sky130_fd_sc_hd__and3_4_16/X sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__and2_0_38/A sky130_fd_sc_hd__nor2_2_19/Y sky130_fd_sc_hd__and2_0_49/A
+ sky130_fd_sc_hd__o21ai_1_450/B1 sky130_fd_sc_hd__nor2b_2_3/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_191 vssd1 vccd1 sky130_fd_sc_hd__buf_8_32/A sky130_fd_sc_hd__buf_8_34/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_262 vccd1 vssd1 sky130_fd_sc_hd__and3_4_10/X sky130_fd_sc_hd__and2_0_87/A
+ sky130_fd_sc_hd__buf_6_0/X sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__o21ai_1_464/B1 sky130_fd_sc_hd__and2b_4_7/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_410 sky130_fd_sc_hd__fa_2_408/CIN sky130_fd_sc_hd__fa_2_411/A
+ sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__fa_2_410/B sky130_fd_sc_hd__xor2_1_621/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_273 vccd1 vssd1 sky130_fd_sc_hd__and3_4_11/X sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__buf_4_3/X sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__o21ai_1_478/B1 sky130_fd_sc_hd__and2b_4_8/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_421 sky130_fd_sc_hd__fah_1_17/B sky130_fd_sc_hd__fa_2_421/SUM
+ sky130_fd_sc_hd__fa_2_421/A sky130_fd_sc_hd__fa_2_421/B sky130_fd_sc_hd__fa_2_421/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_284 vccd1 vssd1 sky130_fd_sc_hd__and3_4_10/X sky130_fd_sc_hd__and2_0_49/A
+ sky130_fd_sc_hd__and2_0_45/A sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__and2_0_87/A
+ sky130_fd_sc_hd__o21ai_1_492/B1 sky130_fd_sc_hd__and2b_4_7/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_432 sky130_fd_sc_hd__fa_2_428/A sky130_fd_sc_hd__fa_2_433/B
+ sky130_fd_sc_hd__fa_2_432/A sky130_fd_sc_hd__fa_2_432/B sky130_fd_sc_hd__o22ai_1_72/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_295 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__buf_4_5/X sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__o21ai_1_505/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_443 sky130_fd_sc_hd__nor2_1_249/A sky130_fd_sc_hd__or2_0_96/B
+ sky130_fd_sc_hd__fa_2_443/A sky130_fd_sc_hd__fa_2_443/B sky130_fd_sc_hd__o22ai_1_89/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_454 sky130_fd_sc_hd__fa_2_453/CIN sky130_fd_sc_hd__fah_1_18/B
+ sky130_fd_sc_hd__fa_2_454/A sky130_fd_sc_hd__fa_2_454/B sky130_fd_sc_hd__ha_2_16/COUT
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_465 sky130_fd_sc_hd__fa_2_462/B sky130_fd_sc_hd__fa_2_464/A
+ sky130_fd_sc_hd__fa_2_465/A sky130_fd_sc_hd__fa_2_465/B sky130_fd_sc_hd__nor2b_1_31/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_476 sky130_fd_sc_hd__nor2_1_257/B sky130_fd_sc_hd__or2_0_103/A
+ sky130_fd_sc_hd__fa_2_476/A sky130_fd_sc_hd__fa_2_476/B sky130_fd_sc_hd__nor2b_1_51/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_487 sky130_fd_sc_hd__or2_0_108/B sky130_fd_sc_hd__nor2_1_263/A
+ sky130_fd_sc_hd__fa_2_487/A sky130_fd_sc_hd__fa_2_487/B sky130_fd_sc_hd__nor2b_1_73/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor2_1_208 sky130_fd_sc_hd__nor2_1_210/Y sky130_fd_sc_hd__nor2_1_208/Y
+ sky130_fd_sc_hd__nor2_1_212/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_219 sky130_fd_sc_hd__xor2_1_633/X sky130_fd_sc_hd__nor2_1_219/Y
+ sky130_fd_sc_hd__nor2_1_219/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_404 sky130_fd_sc_hd__buf_12_404/A sky130_fd_sc_hd__buf_12_527/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_415 sky130_fd_sc_hd__buf_12_68/X sky130_fd_sc_hd__buf_12_628/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_426 sky130_fd_sc_hd__buf_12_426/A sky130_fd_sc_hd__buf_12_485/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_437 sky130_fd_sc_hd__buf_12_437/A sky130_fd_sc_hd__buf_12_583/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_448 sky130_fd_sc_hd__buf_12_448/A sky130_fd_sc_hd__buf_12_599/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_459 sky130_fd_sc_hd__buf_12_459/A sky130_fd_sc_hd__buf_12_612/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_604 sky130_fd_sc_hd__xnor2_1_181/B sky130_fd_sc_hd__o21ai_2_17/A2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_615 sky130_fd_sc_hd__clkinv_1_615/Y sky130_fd_sc_hd__inv_2_52/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_626 sky130_fd_sc_hd__nand2_1_664/A sky130_fd_sc_hd__nor2_1_221/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_637 sky130_fd_sc_hd__clkinv_1_637/Y sky130_fd_sc_hd__nand2_1_687/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_648 sky130_fd_sc_hd__nand2_1_708/A sky130_fd_sc_hd__nor2_1_232/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_659 sky130_fd_sc_hd__nand2_1_723/A sky130_fd_sc_hd__nor2_1_234/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1109 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_190 vssd1 vccd1 sky130_fd_sc_hd__buf_2_3/X sky130_fd_sc_hd__nand2b_1_3/Y
+ sky130_fd_sc_hd__a222oi_1_67/Y sky130_fd_sc_hd__xor2_1_19/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_13 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_354/Q sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__o211ai_1_29/Y sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__a222oi_1_13/Y sky130_fd_sc_hd__dfxtp_1_305/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_600 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_24 vccd1 vssd1 sky130_fd_sc_hd__xor2_1_421/X sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__xor2_1_634/X sky130_fd_sc_hd__xor2_1_209/X sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_24/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_35 vccd1 vssd1 sky130_fd_sc_hd__xnor2_1_98/Y sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__xnor2_1_161/Y sky130_fd_sc_hd__xnor2_1_35/Y sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_35/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_611 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_622 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_46 vccd1 vssd1 sky130_fd_sc_hd__xnor2_1_73/Y sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__inv_2_63/A sky130_fd_sc_hd__xnor2_1_10/Y sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_46/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_633 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_57 vccd1 vssd1 sky130_fd_sc_hd__and3_4_8/X sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__buf_4_3/X sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__a222oi_1_57/Y sky130_fd_sc_hd__nor2b_2_2/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_644 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_68 vccd1 vssd1 sky130_fd_sc_hd__and3_4_6/X sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__buf_6_1/X sky130_fd_sc_hd__nor2_1_72/Y sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__a222oi_1_68/Y sky130_fd_sc_hd__nor2b_1_6/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_655 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_79 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__or2_0_60/B
+ sky130_fd_sc_hd__or2_0_60/A sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__or2_0_61/A
+ sky130_fd_sc_hd__a222oi_1_79/Y sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__xnor2_1_15 vssd1 vccd1 sky130_fd_sc_hd__o21ai_2_6/Y sky130_fd_sc_hd__xnor2_1_15/Y
+ sky130_fd_sc_hd__xnor2_1_15/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_666 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_26 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_26/B sky130_fd_sc_hd__inv_2_10/A
+ sky130_fd_sc_hd__xnor2_1_26/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_550 sky130_fd_sc_hd__nand2_1_550/Y sky130_fd_sc_hd__nor2_2_23/A
+ sky130_fd_sc_hd__nor2_2_23/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_677 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_37 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_37/B sky130_fd_sc_hd__inv_2_22/A
+ sky130_fd_sc_hd__xnor2_1_37/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_561 sky130_fd_sc_hd__nand2_1_561/Y sky130_fd_sc_hd__nor2_2_26/A
+ sky130_fd_sc_hd__nor2_2_26/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_688 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_48 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_183/A sky130_fd_sc_hd__and3_4_1/C
+ sky130_fd_sc_hd__xnor2_1_51/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_572 sky130_fd_sc_hd__nand2_1_572/Y sky130_fd_sc_hd__nand2_1_582/Y
+ sky130_fd_sc_hd__nand2_1_578/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_59 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_61/A sky130_fd_sc_hd__and3_4_3/C
+ sky130_fd_sc_hd__xor2_1_206/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_699 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_583 sky130_fd_sc_hd__nand2_1_583/Y sky130_fd_sc_hd__nand2_1_596/Y
+ sky130_fd_sc_hd__nand2_1_590/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_594 sky130_fd_sc_hd__nand2_1_594/Y sky130_fd_sc_hd__nor2_1_192/Y
+ sky130_fd_sc_hd__nand2_1_599/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_1130 sky130_fd_sc_hd__clkinv_4_73/A sky130_fd_sc_hd__a22o_1_50/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1141 sky130_fd_sc_hd__buf_2_184/A sky130_fd_sc_hd__inv_4_15/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1610 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_2_4 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_4/Y sky130_fd_sc_hd__xnor2_2_4/A
+ sky130_fd_sc_hd__xnor2_2_4/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_2
Xsky130_fd_sc_hd__decap_12_1621 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1632 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1643 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1654 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1665 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1676 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1687 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_390 sky130_fd_sc_hd__dfxtp_1_390/Q sky130_fd_sc_hd__dfxtp_1_392/CLK
+ sky130_fd_sc_hd__nor2b_1_93/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1698 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__or4_1_1 sky130_fd_sc_hd__or4_1_1/C sky130_fd_sc_hd__ha_2_7/A sky130_fd_sc_hd__or4_1_1/X
+ sky130_fd_sc_hd__or4_1_1/B sky130_fd_sc_hd__or4_1_2/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__or4_1
Xsky130_fd_sc_hd__fa_2_240 sky130_fd_sc_hd__nor2_2_15/A sky130_fd_sc_hd__or2_0_35/B
+ sky130_fd_sc_hd__fa_2_240/A sky130_fd_sc_hd__fa_2_240/B sky130_fd_sc_hd__fa_2_240/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_251 sky130_fd_sc_hd__fah_1_3/B sky130_fd_sc_hd__fah_1_2/CI
+ sky130_fd_sc_hd__fa_2_251/A sky130_fd_sc_hd__fa_2_251/B sky130_fd_sc_hd__fah_1_5/COUT
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_262 sky130_fd_sc_hd__fa_2_258/CIN sky130_fd_sc_hd__fa_2_260/A
+ sky130_fd_sc_hd__fa_2_262/A sky130_fd_sc_hd__fa_2_262/B sky130_fd_sc_hd__xor2_1_382/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_273 sky130_fd_sc_hd__fa_2_271/CIN sky130_fd_sc_hd__fa_2_274/B
+ sky130_fd_sc_hd__fa_2_273/A sky130_fd_sc_hd__fa_2_273/B sky130_fd_sc_hd__xor2_1_401/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_284 sky130_fd_sc_hd__xor3_1_22/C sky130_fd_sc_hd__fa_2_286/CIN
+ sky130_fd_sc_hd__fa_2_284/A sky130_fd_sc_hd__fa_2_284/B sky130_fd_sc_hd__xor2_1_441/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_0 vccd1 vssd1 sky130_fd_sc_hd__and2_0_0/X la_data_out[36]
+ sky130_fd_sc_hd__nor2_4_0/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__fa_2_295 sky130_fd_sc_hd__fa_2_286/A sky130_fd_sc_hd__fa_2_296/A
+ sky130_fd_sc_hd__fa_2_295/A sky130_fd_sc_hd__fa_2_295/B sky130_fd_sc_hd__xor2_1_455/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22oi_1_6 sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__a22oi_1_6/B2 sky130_fd_sc_hd__a22oi_1_6/A2 sky130_fd_sc_hd__nand2_2_2/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_201 sky130_fd_sc_hd__buf_6_60/X sky130_fd_sc_hd__buf_12_369/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_212 sky130_fd_sc_hd__buf_6_83/X sky130_fd_sc_hd__buf_12_212/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_223 sky130_fd_sc_hd__buf_6_56/X sky130_fd_sc_hd__buf_12_455/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_70 sky130_fd_sc_hd__xnor2_1_91/B sky130_fd_sc_hd__a21oi_1_70/B1
+ sky130_fd_sc_hd__xor2_1_313/A sky130_fd_sc_hd__or2_0_34/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_234 sky130_fd_sc_hd__buf_6_72/X sky130_fd_sc_hd__buf_12_393/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_81 sky130_fd_sc_hd__nand2_1_400/Y sky130_fd_sc_hd__o21ai_1_498/Y
+ sky130_fd_sc_hd__o21a_1_2/A2 sky130_fd_sc_hd__nor2_1_123/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_245 sky130_fd_sc_hd__buf_6_42/X sky130_fd_sc_hd__buf_12_338/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_92 sky130_fd_sc_hd__nor2_1_143/Y sky130_fd_sc_hd__nand2_1_432/Y
+ sky130_fd_sc_hd__a21oi_1_92/Y sky130_fd_sc_hd__nand2_1_443/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_1_104 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_182/Q sky130_fd_sc_hd__dfxtp_1_150/Q sky130_fd_sc_hd__o21ai_1_10/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_256 sky130_fd_sc_hd__buf_12_256/A sky130_fd_sc_hd__buf_12_389/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_115 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_171/Q sky130_fd_sc_hd__dfxtp_1_139/Q sky130_fd_sc_hd__o21ai_1_21/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_267 sky130_fd_sc_hd__buf_6_46/X sky130_fd_sc_hd__buf_12_267/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_126 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_160/Q sky130_fd_sc_hd__dfxtp_1_128/Q sky130_fd_sc_hd__o21ai_1_32/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_278 sky130_fd_sc_hd__buf_12_278/A sky130_fd_sc_hd__buf_12_604/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_137 sky130_fd_sc_hd__xor2_1_255/X sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xor2_1_42/X sky130_fd_sc_hd__o21ai_1_53/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_289 sky130_fd_sc_hd__buf_12_63/X sky130_fd_sc_hd__buf_12_515/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_148 sky130_fd_sc_hd__xor2_1_313/X sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xor2_1_100/X sky130_fd_sc_hd__o21ai_1_76/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_159 sky130_fd_sc_hd__xor2_1_367/X sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xor2_1_154/X sky130_fd_sc_hd__o21ai_1_99/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_401 sky130_fd_sc_hd__nand2_1_310/A sky130_fd_sc_hd__nor2_2_6/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_412 sky130_fd_sc_hd__xor2_2_1/B sky130_fd_sc_hd__a21oi_1_69/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_423 sky130_fd_sc_hd__nor2_1_111/B sky130_fd_sc_hd__nand2_1_354/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_434 sky130_fd_sc_hd__a21oi_2_8/B1 sky130_fd_sc_hd__nand2_1_362/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_445 sky130_fd_sc_hd__a21oi_1_80/A1 sky130_fd_sc_hd__o21a_1_2/A2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_456 sky130_fd_sc_hd__o21ai_1_515/A1 sky130_fd_sc_hd__nor2_1_126/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_467 sky130_fd_sc_hd__o21ai_1_562/A2 sky130_fd_sc_hd__nand2_1_421/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_478 sky130_fd_sc_hd__nand2_1_430/A sky130_fd_sc_hd__nor2_1_142/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_489 sky130_fd_sc_hd__nand2_1_448/A sky130_fd_sc_hd__nor2_1_150/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a222oi_1_1 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_342/Q sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__o211ai_1_17/Y sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__a222oi_1_1/Y sky130_fd_sc_hd__dfxtp_1_293/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_430 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_441 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_452 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_463 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_474 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_485 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_496 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_380 sky130_fd_sc_hd__nor2_1_123/A sky130_fd_sc_hd__or2_0_46/X
+ sky130_fd_sc_hd__or2_0_47/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_208 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__xor2_1_208/X
+ sky130_fd_sc_hd__xor2_1_208/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_391 sky130_fd_sc_hd__xnor2_1_89/A sky130_fd_sc_hd__nand2_1_392/Y
+ sky130_fd_sc_hd__or2_0_47/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_990 sky130_fd_sc_hd__clkinv_1_990/Y sky130_fd_sc_hd__clkinv_2_35/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xor2_1_219 sky130_fd_sc_hd__xor2_1_362/B sky130_fd_sc_hd__xor3_1_18/B
+ sky130_fd_sc_hd__xor2_1_219/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1440 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1451 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1462 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1473 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_904 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_687/A sky130_fd_sc_hd__nor2_1_265/Y
+ sky130_fd_sc_hd__nand2_1_837/Y sky130_fd_sc_hd__xnor2_1_301/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1484 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_915 vssd1 vccd1 sky130_fd_sc_hd__ha_2_53/SUM sky130_fd_sc_hd__o21ai_1_915/A1
+ sky130_fd_sc_hd__a21oi_1_189/Y sky130_fd_sc_hd__o21ai_1_915/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1495 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_926 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_926/A2 sky130_fd_sc_hd__a21o_2_1/B1
+ sky130_fd_sc_hd__or3_1_0/X sky130_fd_sc_hd__o21ai_1_926/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_8_8 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__buf_2_13 vccd1 vssd1 sky130_fd_sc_hd__buf_2_13/X sky130_fd_sc_hd__buf_2_13/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_24 vccd1 vssd1 sky130_fd_sc_hd__buf_2_24/X sky130_fd_sc_hd__buf_4_0/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_35 vccd1 vssd1 sky130_fd_sc_hd__buf_8_82/A sky130_fd_sc_hd__ha_2_30/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_46 vccd1 vssd1 sky130_fd_sc_hd__buf_2_46/X sky130_fd_sc_hd__buf_2_46/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_57 vccd1 vssd1 sky130_fd_sc_hd__buf_8_3/A sky130_fd_sc_hd__buf_8_5/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_68 vccd1 vssd1 sky130_fd_sc_hd__buf_6_9/A sky130_fd_sc_hd__buf_2_68/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_79 vccd1 vssd1 sky130_fd_sc_hd__buf_2_79/X sky130_fd_sc_hd__buf_2_79/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o211ai_1_40 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o22ai_1_23/B1
+ sky130_fd_sc_hd__fa_2_346/A sky130_fd_sc_hd__nand2_1_60/Y sky130_fd_sc_hd__a21oi_1_11/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_51 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o22ai_1_12/B1
+ sky130_fd_sc_hd__fah_1_14/B sky130_fd_sc_hd__nand2_1_71/Y sky130_fd_sc_hd__a21oi_1_22/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_62 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o22ai_1_1/B1
+ sky130_fd_sc_hd__nor2_1_220/A sky130_fd_sc_hd__nand2_1_82/Y sky130_fd_sc_hd__a21oi_1_33/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__diode_2_8 sky130_fd_sc_hd__conb_1_147/HI vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__xor3_1_19 sky130_fd_sc_hd__xor3_1_19/X sky130_fd_sc_hd__xor3_1_19/C
+ sky130_fd_sc_hd__xor3_1_19/B sky130_fd_sc_hd__xor3_1_19/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__clkinv_1_220 sky130_fd_sc_hd__o22ai_1_8/A2 sky130_fd_sc_hd__dfxtp_1_167/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_231 sky130_fd_sc_hd__o22ai_1_5/B1 sky130_fd_sc_hd__dfxtp_1_100/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_242 sky130_fd_sc_hd__nor2_1_5/A sky130_fd_sc_hd__dfxtp_1_128/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_253 sky130_fd_sc_hd__o21ai_1_99/A2 sky130_fd_sc_hd__xor2_1_580/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_264 sky130_fd_sc_hd__o21ai_1_145/A2 sky130_fd_sc_hd__xnor2_1_182/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_275 sky130_fd_sc_hd__and2_0_136/A sky130_fd_sc_hd__a222oi_1_19/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_286 sky130_fd_sc_hd__and2_0_201/A sky130_fd_sc_hd__a222oi_1_30/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_297 sky130_fd_sc_hd__and2_0_236/A sky130_fd_sc_hd__a222oi_1_41/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xor3_1_4 sky130_fd_sc_hd__xor3_1_4/X sky130_fd_sc_hd__xor3_1_4/C
+ sky130_fd_sc_hd__xor3_1_4/B sky130_fd_sc_hd__xor3_1_5/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__a21oi_1_5 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_34/Y
+ sky130_fd_sc_hd__a21oi_1_5/Y sky130_fd_sc_hd__dfxtp_1_90/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__and3_4_11 sky130_fd_sc_hd__nor2_4_13/B sky130_fd_sc_hd__nor2_4_13/A
+ sky130_fd_sc_hd__and3_4_11/C sky130_fd_sc_hd__and3_4_11/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__clkbuf_4_18 sky130_fd_sc_hd__clkbuf_4_18/X sky130_fd_sc_hd__buf_6_8/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and3_4_22 sky130_fd_sc_hd__nor2_4_18/B sky130_fd_sc_hd__nor2_4_18/A
+ sky130_fd_sc_hd__and3_4_22/C sky130_fd_sc_hd__and3_4_22/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__clkbuf_4_29 sky130_fd_sc_hd__clkbuf_4_29/X sky130_fd_sc_hd__buf_8_159/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__a21oi_1_150 sky130_fd_sc_hd__or2_0_83/X sky130_fd_sc_hd__clkinv_1_649/Y
+ sky130_fd_sc_hd__xor2_1_651/A sky130_fd_sc_hd__xnor2_1_200/A vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_161 sky130_fd_sc_hd__xnor2_1_213/B sky130_fd_sc_hd__clkinv_1_681/Y
+ sky130_fd_sc_hd__xor2_1_661/A sky130_fd_sc_hd__nand2_1_758/A vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_172 sky130_fd_sc_hd__xnor2_1_293/B sky130_fd_sc_hd__clkinv_1_812/Y
+ sky130_fd_sc_hd__xor2_1_678/A sky130_fd_sc_hd__or2_0_102/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_183 sky130_fd_sc_hd__nand3_1_5/C sky130_fd_sc_hd__a21oi_1_184/Y
+ sky130_fd_sc_hd__nand2_1_848/A sky130_fd_sc_hd__o21ai_1_907/Y vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_194 sky130_fd_sc_hd__ha_2_53/SUM sky130_fd_sc_hd__ha_2_53/COUT
+ sky130_fd_sc_hd__nand2_1_858/A sky130_fd_sc_hd__o21ai_1_915/A1 vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_102 sky130_fd_sc_hd__inv_2_173/A sky130_fd_sc_hd__buf_8_102/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_113 sky130_fd_sc_hd__buf_8_113/A sky130_fd_sc_hd__buf_6_31/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_124 sky130_fd_sc_hd__buf_8_124/A sky130_fd_sc_hd__buf_8_124/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_135 sky130_fd_sc_hd__inv_2_185/Y sky130_fd_sc_hd__buf_8_135/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_146 sky130_fd_sc_hd__buf_8_146/A sky130_fd_sc_hd__buf_8_146/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nor2_4_8 sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__or2b_2_0/A
+ sky130_fd_sc_hd__nor2_4_8/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__buf_8_157 sky130_fd_sc_hd__buf_8_157/A sky130_fd_sc_hd__buf_8_157/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__decap_12_260 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_271 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_282 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_293 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1270 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_701 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_126/Y sky130_fd_sc_hd__nand2b_2_6/Y
+ sky130_fd_sc_hd__o21ai_1_701/B1 sky130_fd_sc_hd__xor2_1_480/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1281 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_712 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_742/A2 sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_712/B1 sky130_fd_sc_hd__xor2_1_490/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1292 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_723 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_723/A2 sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_723/B1 sky130_fd_sc_hd__xor2_1_500/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_734 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_10/X sky130_fd_sc_hd__or2_0_55/B
+ sky130_fd_sc_hd__o21a_1_4/A2 sky130_fd_sc_hd__xnor2_1_148/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_745 vssd1 vccd1 sky130_fd_sc_hd__inv_2_46/Y sky130_fd_sc_hd__nand2b_1_21/Y
+ sky130_fd_sc_hd__o21ai_1_745/B1 sky130_fd_sc_hd__xor2_1_520/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_756 vssd1 vccd1 sky130_fd_sc_hd__inv_2_45/Y sky130_fd_sc_hd__nand2b_2_6/Y
+ sky130_fd_sc_hd__o21ai_1_756/B1 sky130_fd_sc_hd__xor2_1_531/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_767 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_767/A2 sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_767/B1 sky130_fd_sc_hd__xor2_1_542/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_778 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_9/X sky130_fd_sc_hd__nand2b_1_16/Y
+ sky130_fd_sc_hd__o21ai_1_778/B1 sky130_fd_sc_hd__xor2_1_552/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_789 vssd1 vccd1 sky130_fd_sc_hd__xor2_2_2/X sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_789/B1 sky130_fd_sc_hd__xor2_1_563/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_30 sky130_fd_sc_hd__fa_2_75/A sky130_fd_sc_hd__fa_2_13/B
+ sky130_fd_sc_hd__xor2_1_30/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_41 sky130_fd_sc_hd__fa_2_97/A sky130_fd_sc_hd__fa_2_23/B
+ sky130_fd_sc_hd__xor2_1_41/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_52 sky130_fd_sc_hd__fa_2_75/A sky130_fd_sc_hd__fa_2_31/B
+ sky130_fd_sc_hd__xor2_1_52/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_63 sky130_fd_sc_hd__xor2_1_63/B sky130_fd_sc_hd__xor2_1_63/X
+ sky130_fd_sc_hd__xor2_1_63/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_19 sky130_fd_sc_hd__buf_12_19/A sky130_fd_sc_hd__buf_12_19/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_74 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__fa_2_54/A
+ sky130_fd_sc_hd__xor2_1_74/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_85 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__fa_2_62/B
+ sky130_fd_sc_hd__xor2_1_85/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_96 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__fa_2_68/A
+ sky130_fd_sc_hd__xor2_1_96/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2b_1_2 sky130_fd_sc_hd__nand2b_1_2/Y sky130_fd_sc_hd__xnor2_1_8/Y
+ sky130_fd_sc_hd__xnor2_1_5/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__o21ai_2_17 sky130_fd_sc_hd__o21ai_2_17/B1 sky130_fd_sc_hd__inv_2_52/A
+ sky130_fd_sc_hd__o21ai_2_17/A2 sky130_fd_sc_hd__o21ai_2_17/A1 vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__o21ai_2
Xsky130_fd_sc_hd__xor2_1_550 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__fa_2_369/A
+ sky130_fd_sc_hd__xor2_1_550/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_561 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__fa_2_380/B
+ sky130_fd_sc_hd__xor2_1_561/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_572 sky130_fd_sc_hd__xor2_1_572/B sky130_fd_sc_hd__xor2_1_572/X
+ sky130_fd_sc_hd__xor2_1_572/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_583 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__xor2_1_583/X
+ sky130_fd_sc_hd__xor2_1_583/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_594 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__fa_2_398/B
+ sky130_fd_sc_hd__xor2_1_594/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a221oi_1_0 sky130_fd_sc_hd__nand4_1_1/C sky130_fd_sc_hd__o22ai_1_136/Y
+ sky130_fd_sc_hd__a221oi_1_0/A1 sky130_fd_sc_hd__dfxtp_1_360/Q sky130_fd_sc_hd__nand4_1_0/D
+ sky130_fd_sc_hd__dfxtp_1_359/Q vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__a221oi_1
Xsky130_fd_sc_hd__a222oi_1_603 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_421/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_453/Q sky130_fd_sc_hd__nor2_4_19/B
+ sky130_fd_sc_hd__clkinv_1_800/A sky130_fd_sc_hd__dfxtp_1_389/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a32oi_1_0 sky130_fd_sc_hd__o21ai_2_0/B1 sky130_fd_sc_hd__a32oi_1_0/Y
+ sky130_fd_sc_hd__inv_2_5/A sky130_fd_sc_hd__o21ai_2_0/B1 sky130_fd_sc_hd__o21ai_2_1/A2
+ sky130_fd_sc_hd__inv_2_7/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__a32oi_1
Xsky130_fd_sc_hd__and2_0_13 vccd1 vssd1 sky130_fd_sc_hd__and2_0_13/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_13/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_24 vccd1 vssd1 sky130_fd_sc_hd__and2_0_24/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__buf_2_24/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_35 vccd1 vssd1 sky130_fd_sc_hd__and2_0_35/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__buf_2_29/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_46 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_2_2/D sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__nor2_2_10/B vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_57 vccd1 vssd1 sky130_fd_sc_hd__and2_0_57/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__or2_0_4/B vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_68 vccd1 vssd1 sky130_fd_sc_hd__and2_0_68/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__or2_0_61/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_79 vccd1 vssd1 sky130_fd_sc_hd__and2_0_79/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__buf_6_4/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nor2_2_5 sky130_fd_sc_hd__nor2_2_5/B sky130_fd_sc_hd__nor2_2_5/Y
+ sky130_fd_sc_hd__nor2_2_5/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__buf_8_12 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__buf_8_12/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_23 sky130_fd_sc_hd__buf_8_23/A sky130_fd_sc_hd__buf_8_23/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_34 sky130_fd_sc_hd__buf_8_34/A sky130_fd_sc_hd__buf_8_34/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_45 sky130_fd_sc_hd__inv_2_78/Y sky130_fd_sc_hd__buf_8_45/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_56 sky130_fd_sc_hd__buf_8_70/A sky130_fd_sc_hd__buf_8_56/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_67 sky130_fd_sc_hd__buf_8_67/A sky130_fd_sc_hd__buf_8_67/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xnor2_1_180 vssd1 vccd1 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__nor2_4_17/A
+ sky130_fd_sc_hd__xnor2_1_180/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__buf_8_78 sky130_fd_sc_hd__buf_8_78/A sky130_fd_sc_hd__buf_8_78/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xnor2_1_191 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_191/B sky130_fd_sc_hd__and2_0_271/A
+ sky130_fd_sc_hd__xnor2_1_191/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__buf_8_89 sky130_fd_sc_hd__buf_8_89/A sky130_fd_sc_hd__buf_8_89/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_208 sky130_fd_sc_hd__xor2_1_530/A sky130_fd_sc_hd__dfxtp_2_0/CLK
+ sky130_fd_sc_hd__and2_0_65/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_219 sky130_fd_sc_hd__xor2_1_424/A sky130_fd_sc_hd__dfxtp_2_5/CLK
+ sky130_fd_sc_hd__and2_0_32/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_520 vssd1 vccd1 sky130_fd_sc_hd__inv_2_35/Y sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_520/B1 sky130_fd_sc_hd__xor2_1_319/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_531 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_7/X sky130_fd_sc_hd__nand2_1_395/Y
+ sky130_fd_sc_hd__a21oi_1_83/Y sky130_fd_sc_hd__xnor2_1_92/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_542 vssd1 vccd1 sky130_fd_sc_hd__buf_2_9/X sky130_fd_sc_hd__nand2b_2_3/Y
+ sky130_fd_sc_hd__o21ai_1_542/B1 sky130_fd_sc_hd__xor2_1_340/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_553 vssd1 vccd1 sky130_fd_sc_hd__buf_2_7/X sky130_fd_sc_hd__nand2b_1_8/Y
+ sky130_fd_sc_hd__o21ai_1_553/B1 sky130_fd_sc_hd__xor2_1_351/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_564 vssd1 vccd1 sky130_fd_sc_hd__inv_2_27/Y sky130_fd_sc_hd__nand2b_1_8/Y
+ sky130_fd_sc_hd__nand2_1_327/Y sky130_fd_sc_hd__xor2_1_361/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_575 vssd1 vccd1 sky130_fd_sc_hd__inv_2_29/Y sky130_fd_sc_hd__nand2b_2_3/Y
+ sky130_fd_sc_hd__o21ai_1_575/B1 sky130_fd_sc_hd__xor2_1_372/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_586 vssd1 vccd1 sky130_fd_sc_hd__buf_2_11/X sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_586/B1 sky130_fd_sc_hd__xor2_1_379/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_597 vssd1 vccd1 sky130_fd_sc_hd__inv_2_28/Y sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_597/B1 sky130_fd_sc_hd__xor2_1_391/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__buf_2_108 vccd1 vssd1 sky130_fd_sc_hd__buf_2_108/X sky130_fd_sc_hd__buf_2_108/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_119 vccd1 vssd1 sky130_fd_sc_hd__buf_2_119/X sky130_fd_sc_hd__buf_2_119/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__xor2_1_380 sky130_fd_sc_hd__fa_2_281/A sky130_fd_sc_hd__fa_2_261/A
+ sky130_fd_sc_hd__xor2_1_380/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_391 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__fa_2_268/B
+ sky130_fd_sc_hd__xor2_1_391/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__ha_2_8 vssd1 vccd1 sky130_fd_sc_hd__ha_2_8/A sky130_fd_sc_hd__ha_2_7/B
+ sky130_fd_sc_hd__nor3_1_0/B sky130_fd_sc_hd__ha_2_8/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__a222oi_1_400 vccd1 vssd1 sky130_fd_sc_hd__and3_1_2/X sky130_fd_sc_hd__or2_0_52/B
+ sky130_fd_sc_hd__buf_2_25/A sky130_fd_sc_hd__nor2_1_174/Y sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__o21ai_1_666/B1 sky130_fd_sc_hd__nor2b_1_14/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_340 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1_11/D sky130_fd_sc_hd__dfxtp_1_12/Q
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_411 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__or2_0_61/B
+ sky130_fd_sc_hd__or2_0_58/B sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__or2_0_58/A
+ sky130_fd_sc_hd__o21ai_1_679/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_351 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2_1/A sky130_fd_sc_hd__a222oi_1_5/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_422 vccd1 vssd1 sky130_fd_sc_hd__and3_4_23/X sky130_fd_sc_hd__buf_2_25/A
+ sky130_fd_sc_hd__inv_6_0/Y sky130_fd_sc_hd__nor2_1_178/Y sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__o21ai_1_695/B1 sky130_fd_sc_hd__nor2b_1_15/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_433 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__or2_0_66/A sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__or2_0_60/B
+ sky130_fd_sc_hd__o21ai_1_707/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_444 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__buf_4_4/X sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__o21ai_1_722/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_455 vccd1 vssd1 sky130_fd_sc_hd__and3_4_26/X sky130_fd_sc_hd__buf_2_24/X
+ sky130_fd_sc_hd__buf_2_27/X sky130_fd_sc_hd__nor2_2_31/Y sky130_fd_sc_hd__buf_2_15/X
+ sky130_fd_sc_hd__o21ai_1_737/B1 sky130_fd_sc_hd__nor2b_1_12/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_466 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__buf_4_3/X sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__o21ai_1_750/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_477 vccd1 vssd1 sky130_fd_sc_hd__and3_4_21/X sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__nor2_1_85/B sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__nor2_2_10/B
+ sky130_fd_sc_hd__o21ai_1_764/B1 sky130_fd_sc_hd__and2b_4_12/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_19 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_9/B2 sky130_fd_sc_hd__inv_4_7/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_488 vccd1 vssd1 sky130_fd_sc_hd__and3_4_18/X sky130_fd_sc_hd__buf_2_30/X
+ sky130_fd_sc_hd__buf_2_26/X sky130_fd_sc_hd__nor2_2_32/Y sky130_fd_sc_hd__buf_2_24/X
+ sky130_fd_sc_hd__o21ai_1_778/B1 sky130_fd_sc_hd__nor2b_2_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_499 vccd1 vssd1 sky130_fd_sc_hd__and3_4_20/X sky130_fd_sc_hd__buf_2_26/X
+ sky130_fd_sc_hd__buf_2_24/X sky130_fd_sc_hd__nor2_4_16/Y sky130_fd_sc_hd__buf_2_27/X
+ sky130_fd_sc_hd__o21ai_1_792/B1 sky130_fd_sc_hd__and2b_4_11/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__and2_0_360 vccd1 vssd1 sky130_fd_sc_hd__and2_0_360/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__buf_2_49/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_371 vccd1 vssd1 sky130_fd_sc_hd__and2_0_371/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_64/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_382 vccd1 vssd1 sky130_fd_sc_hd__and2_0_382/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_78/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_393 vccd1 vssd1 sky130_fd_sc_hd__and2_0_393/X sky130_fd_sc_hd__and2_0_401/B
+ sky130_fd_sc_hd__and2_0_393/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__conb_1_2 sky130_fd_sc_hd__conb_1_2/LO sky130_fd_sc_hd__conb_1_2/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__buf_12_8 sky130_fd_sc_hd__buf_12_8/A sky130_fd_sc_hd__buf_12_8/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_608 sky130_fd_sc_hd__buf_12_608/A sky130_fd_sc_hd__buf_12_608/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__inv_2_160 sky130_fd_sc_hd__inv_2_160/A sky130_fd_sc_hd__inv_4_10/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_12_619 sky130_fd_sc_hd__buf_12_619/A sky130_fd_sc_hd__buf_12_619/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__inv_2_171 sky130_fd_sc_hd__inv_2_171/A sky130_fd_sc_hd__inv_2_171/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_182 sky130_fd_sc_hd__inv_2_182/A sky130_fd_sc_hd__inv_2_182/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_193 sky130_fd_sc_hd__inv_2_71/A sky130_fd_sc_hd__ha_2_34/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__o22ai_1_101 sky130_fd_sc_hd__xnor2_2_4/Y sky130_fd_sc_hd__o22ai_1_101/B1
+ sky130_fd_sc_hd__fa_2_444/B sky130_fd_sc_hd__nand2b_1_26/Y sky130_fd_sc_hd__o22ai_1_96/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_112 sky130_fd_sc_hd__nor2b_1_24/A sky130_fd_sc_hd__o22ai_1_112/B1
+ sky130_fd_sc_hd__ha_2_16/B sky130_fd_sc_hd__nand2b_1_28/Y sky130_fd_sc_hd__nand2_1_722/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_123 sky130_fd_sc_hd__nor2b_1_20/A sky130_fd_sc_hd__xnor2_1_270/Y
+ sky130_fd_sc_hd__fa_2_455/B sky130_fd_sc_hd__xnor2_1_278/Y sky130_fd_sc_hd__o22ai_1_78/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_134 sky130_fd_sc_hd__xnor2_1_289/Y sky130_fd_sc_hd__xnor2_1_288/Y
+ sky130_fd_sc_hd__ha_2_17/A sky130_fd_sc_hd__inv_2_65/Y sky130_fd_sc_hd__o22ai_1_99/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_209 sky130_fd_sc_hd__nor2_1_64/A sky130_fd_sc_hd__or2_0_20/X
+ sky130_fd_sc_hd__or2_0_17/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_808 sky130_fd_sc_hd__clkinv_1_808/Y sky130_fd_sc_hd__nand2_1_795/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_2_12 sky130_fd_sc_hd__nor2_2_12/B sky130_fd_sc_hd__nor2_2_12/Y
+ sky130_fd_sc_hd__nor2_2_12/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__clkinv_1_819 sky130_fd_sc_hd__nand2_1_816/A sky130_fd_sc_hd__nor2_1_260/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_2_23 sky130_fd_sc_hd__nor2_2_23/B sky130_fd_sc_hd__nor2_2_23/Y
+ sky130_fd_sc_hd__nor2_2_23/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__o211ai_1_2 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_2/A2
+ sky130_fd_sc_hd__o211ai_1_2/Y sky130_fd_sc_hd__a22oi_1_36/Y sky130_fd_sc_hd__a22oi_1_37/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__conb_1_19 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__conb_1_19/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__o21ai_1_350 vssd1 vccd1 sky130_fd_sc_hd__inv_2_11/Y sky130_fd_sc_hd__nand2_1_267/Y
+ sky130_fd_sc_hd__a21oi_1_58/Y sky130_fd_sc_hd__xnor2_1_45/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_361 vssd1 vccd1 sky130_fd_sc_hd__buf_2_5/X sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__o21ai_1_361/B1 sky130_fd_sc_hd__xor2_1_177/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_372 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_191/B sky130_fd_sc_hd__nor2_1_98/Y
+ sky130_fd_sc_hd__nand2_1_290/Y sky130_fd_sc_hd__o21ai_1_372/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_383 vssd1 vccd1 sky130_fd_sc_hd__nand2_1_298/Y sky130_fd_sc_hd__a21oi_1_67/Y
+ sky130_fd_sc_hd__a21oi_1_64/Y sky130_fd_sc_hd__xnor2_1_54/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_394 vssd1 vccd1 sky130_fd_sc_hd__inv_2_26/Y sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__nand2_1_161/Y sky130_fd_sc_hd__xor2_1_211/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_804 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_815 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_826 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_710 sky130_fd_sc_hd__xnor2_1_200/B sky130_fd_sc_hd__nand2_1_711/Y
+ sky130_fd_sc_hd__or2_0_83/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_837 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_721 sky130_fd_sc_hd__o22ai_1_99/B2 sky130_fd_sc_hd__inv_2_65/Y
+ la_data_out[77] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_848 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_732 sky130_fd_sc_hd__xnor2_1_207/A sky130_fd_sc_hd__nand2_1_733/Y
+ sky130_fd_sc_hd__nand2_1_732/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_859 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__mux2_2_30 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_30/A1 sky130_fd_sc_hd__buf_2_72/X
+ sky130_fd_sc_hd__mux2_8_0/S sky130_fd_sc_hd__fa_2_417/A vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_743 sky130_fd_sc_hd__xor2_1_656/B sky130_fd_sc_hd__nand2_1_744/Y
+ sky130_fd_sc_hd__nand2_1_743/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_41 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_41/A1 sky130_fd_sc_hd__buf_2_145/X
+ sky130_fd_sc_hd__mux2_8_0/S sky130_fd_sc_hd__or2_0_77/B vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_754 sky130_fd_sc_hd__nand2_1_754/Y sky130_fd_sc_hd__or2_0_95/A
+ sky130_fd_sc_hd__or2_0_95/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_52 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_52/A1 sky130_fd_sc_hd__buf_2_147/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__or2_0_81/A vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_765 sky130_fd_sc_hd__xor2_1_665/A sky130_fd_sc_hd__nand2_1_782/Y
+ sky130_fd_sc_hd__nand2_1_765/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_776 sky130_fd_sc_hd__nand2_1_776/Y sky130_fd_sc_hd__nor2_1_247/A
+ sky130_fd_sc_hd__nor2_1_247/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_787 sky130_fd_sc_hd__or2_0_98/B sky130_fd_sc_hd__nand2b_1_24/Y
+ sky130_fd_sc_hd__o22ai_1_99/B2 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_798 sky130_fd_sc_hd__xnor2_1_292/A sky130_fd_sc_hd__nand2_1_799/Y
+ sky130_fd_sc_hd__or2_0_101/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_1803 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1814 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1825 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1836 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1847 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_550 wbs_dat_o[29] sky130_fd_sc_hd__dfxtp_1_552/CLK sky130_fd_sc_hd__nor2b_1_128/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1858 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1869 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__or2b_2_2 sky130_fd_sc_hd__or2b_2_2/A sky130_fd_sc_hd__nor2_4_15/B
+ sky130_fd_sc_hd__or2b_2_2/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__or2b_2
Xsky130_sram_1kbyte_1rw1r_32x256_8_10 sky130_fd_sc_hd__buf_4_8/X sky130_fd_sc_hd__buf_4_8/X
+ sky130_fd_sc_hd__buf_12_655/X sky130_fd_sc_hd__buf_12_325/X sky130_fd_sc_hd__buf_12_662/X
+ sky130_fd_sc_hd__buf_12_631/X sky130_fd_sc_hd__buf_12_641/X sky130_fd_sc_hd__buf_12_574/X
+ sky130_fd_sc_hd__buf_12_639/X sky130_fd_sc_hd__clkinv_1_955/Y sky130_fd_sc_hd__buf_12_618/X
+ sky130_fd_sc_hd__buf_12_392/X sky130_fd_sc_hd__buf_12_592/X vccd1 sky130_fd_sc_hd__clkinv_8_17/Y
+ sky130_fd_sc_hd__clkbuf_1_145/A sky130_fd_sc_hd__clkbuf_1_144/A sky130_fd_sc_hd__clkbuf_1_80/A
+ sky130_fd_sc_hd__clkbuf_1_79/A sky130_fd_sc_hd__clkbuf_1_78/A sky130_fd_sc_hd__clkbuf_1_77/A
+ sky130_fd_sc_hd__clkbuf_1_314/A sky130_fd_sc_hd__clkbuf_1_75/A sky130_fd_sc_hd__clkbuf_1_274/A
+ sky130_fd_sc_hd__clkbuf_1_74/A sky130_fd_sc_hd__clkbuf_1_73/A sky130_fd_sc_hd__clkbuf_1_72/A
+ sky130_fd_sc_hd__clkbuf_1_71/A sky130_fd_sc_hd__clkbuf_1_70/A sky130_fd_sc_hd__clkbuf_1_69/A
+ sky130_fd_sc_hd__clkbuf_1_68/A sky130_fd_sc_hd__buf_12_585/X sky130_fd_sc_hd__buf_2_155/A
+ sky130_fd_sc_hd__clkbuf_1_304/A sky130_fd_sc_hd__clkbuf_1_87/A sky130_fd_sc_hd__clkbuf_1_86/A
+ sky130_fd_sc_hd__clkbuf_1_85/A sky130_fd_sc_hd__clkbuf_1_84/A sky130_fd_sc_hd__clkbuf_1_83/A
+ sky130_fd_sc_hd__clkbuf_1_82/A sky130_fd_sc_hd__clkbuf_1_81/A sky130_fd_sc_hd__clkbuf_1_159/A
+ sky130_fd_sc_hd__clkbuf_1_158/A sky130_fd_sc_hd__clkbuf_1_156/A sky130_fd_sc_hd__clkbuf_1_153/A
+ sky130_fd_sc_hd__clkbuf_1_146/A sky130_fd_sc_hd__clkbuf_1_148/A sky130_fd_sc_hd__clkbuf_1_157/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[10] sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[11]
+ sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[12] sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[13]
+ sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[14] sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[15]
+ sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[16] sky130_fd_sc_hd__buf_12_663/X sky130_fd_sc_hd__buf_12_259/X
+ sky130_fd_sc_hd__buf_12_29/X sky130_fd_sc_hd__buf_12_258/X sky130_fd_sc_hd__buf_12_19/X
+ sky130_fd_sc_hd__clkinv_8_22/Y sky130_fd_sc_hd__buf_2_51/X sky130_fd_sc_hd__buf_2_50/X
+ sky130_fd_sc_hd__buf_6_6/X sky130_fd_sc_hd__inv_2_107/Y sky130_fd_sc_hd__inv_2_105/Y
+ sky130_fd_sc_hd__buf_2_49/X sky130_fd_sc_hd__buf_2_48/X sky130_fd_sc_hd__clkbuf_1_322/X
+ sky130_fd_sc_hd__buf_2_47/X sky130_fd_sc_hd__buf_2_46/X sky130_fd_sc_hd__buf_2_45/X
+ sky130_fd_sc_hd__clkinv_2_17/Y sky130_fd_sc_hd__buf_2_44/X sky130_fd_sc_hd__buf_2_42/X
+ sky130_fd_sc_hd__clkbuf_1_41/X sky130_fd_sc_hd__clkbuf_4_9/X sky130_fd_sc_hd__clkbuf_1_138/X
+ sky130_fd_sc_hd__clkbuf_1_139/X sky130_fd_sc_hd__buf_2_39/X sky130_fd_sc_hd__clkbuf_1_40/X
+ sky130_fd_sc_hd__clkbuf_1_312/X sky130_fd_sc_hd__clkbuf_1_236/X sky130_fd_sc_hd__clkbuf_1_323/X
+ sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[0] sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[1]
+ sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[2] sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[3]
+ sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[4] sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[5]
+ sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[6] sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[7]
+ sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[8] sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[9]
+ sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[25] sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[26]
+ sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[27] sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[28]
+ sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[29] sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[30]
+ sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[31] sky130_fd_sc_hd__clkinv_1_847/Y sky130_fd_sc_hd__clkinv_1_871/Y
+ sky130_fd_sc_hd__inv_2_95/Y sky130_fd_sc_hd__clkinv_1_866/Y sky130_fd_sc_hd__inv_2_94/Y
+ sky130_fd_sc_hd__clkinv_1_861/Y sky130_fd_sc_hd__clkbuf_1_319/X sky130_fd_sc_hd__clkinv_1_855/Y
+ sky130_fd_sc_hd__clkinv_1_851/Y sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[17] sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[18]
+ sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[19] sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[20]
+ sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[21] sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[22]
+ sky130_fd_sc_hd__buf_12_517/X sky130_fd_sc_hd__buf_12_620/X sky130_fd_sc_hd__buf_12_466/X
+ sky130_fd_sc_hd__buf_12_573/X sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[23] sky130_sram_1kbyte_1rw1r_32x256_8_10/dout0[24]
+ sky130_sram_1kbyte_1rw1r_32x256_8_10/sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/gnd_uq26
+ vssd1 sky130_sram_1kbyte_1rw1r_32x256_8
Xsky130_fd_sc_hd__a222oi_1_230 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__or2_0_58/A
+ sky130_fd_sc_hd__or2_0_9/B sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__or2_0_9/A
+ sky130_fd_sc_hd__o21ai_1_421/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_170 vssd1 vccd1 sky130_fd_sc_hd__a22o_1_33/B2 sky130_fd_sc_hd__clkbuf_1_170/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_241 vccd1 vssd1 sky130_fd_sc_hd__and3_4_17/X sky130_fd_sc_hd__and2_0_87/A
+ sky130_fd_sc_hd__buf_6_0/X sky130_fd_sc_hd__nor2_2_20/Y sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__o21ai_1_437/B1 sky130_fd_sc_hd__nor2b_2_4/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_181 vssd1 vccd1 sky130_fd_sc_hd__a22o_1_23/B2 sky130_fd_sc_hd__clkbuf_1_181/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_252 vccd1 vssd1 sky130_fd_sc_hd__and3_4_15/X sky130_fd_sc_hd__buf_2_31/X
+ sky130_fd_sc_hd__buf_2_19/X sky130_fd_sc_hd__nor2_1_130/Y sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__o21ai_1_451/B1 sky130_fd_sc_hd__nor2b_1_11/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_192 vssd1 vccd1 sky130_fd_sc_hd__buf_12_49/A sky130_fd_sc_hd__buf_8_42/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_400 sky130_fd_sc_hd__fah_1_8/B sky130_fd_sc_hd__fah_1_10/CI
+ sky130_fd_sc_hd__fa_2_400/A sky130_fd_sc_hd__fa_2_400/B sky130_fd_sc_hd__xor2_1_598/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_263 vccd1 vssd1 sky130_fd_sc_hd__and3_4_15/X sky130_fd_sc_hd__buf_4_0/X
+ sky130_fd_sc_hd__buf_2_23/X sky130_fd_sc_hd__nor2_1_130/Y sky130_fd_sc_hd__buf_2_31/X
+ sky130_fd_sc_hd__o21ai_1_465/B1 sky130_fd_sc_hd__nor2b_1_11/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_411 sky130_fd_sc_hd__nor2_1_211/A sky130_fd_sc_hd__or2_0_62/B
+ sky130_fd_sc_hd__fa_2_411/A sky130_fd_sc_hd__fa_2_411/B sky130_fd_sc_hd__fa_2_411/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_274 vccd1 vssd1 sky130_fd_sc_hd__and3_4_15/X sky130_fd_sc_hd__buf_4_7/X
+ sky130_fd_sc_hd__buf_4_0/X sky130_fd_sc_hd__nor2_1_130/Y sky130_fd_sc_hd__buf_2_23/X
+ sky130_fd_sc_hd__o21ai_1_479/B1 sky130_fd_sc_hd__nor2b_1_11/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_422 sky130_fd_sc_hd__fa_2_420/B sky130_fd_sc_hd__fa_2_424/CIN
+ sky130_fd_sc_hd__fa_2_422/A sky130_fd_sc_hd__fa_2_422/B sky130_fd_sc_hd__fa_2_422/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_285 vccd1 vssd1 sky130_fd_sc_hd__and3_4_15/X sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__buf_4_7/X sky130_fd_sc_hd__nor2_1_130/Y sky130_fd_sc_hd__buf_4_0/X
+ sky130_fd_sc_hd__o21ai_1_493/B1 sky130_fd_sc_hd__nor2b_1_11/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_433 sky130_fd_sc_hd__fa_2_430/B sky130_fd_sc_hd__fa_2_434/CIN
+ sky130_fd_sc_hd__fa_2_433/A sky130_fd_sc_hd__fa_2_433/B sky130_fd_sc_hd__fa_2_433/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_296 vccd1 vssd1 sky130_fd_sc_hd__and3_4_16/X sky130_fd_sc_hd__buf_4_7/X
+ sky130_fd_sc_hd__buf_4_0/X sky130_fd_sc_hd__nor2_2_19/Y sky130_fd_sc_hd__buf_2_23/X
+ sky130_fd_sc_hd__o21ai_1_507/B1 sky130_fd_sc_hd__nor2b_2_3/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_444 sky130_fd_sc_hd__nor2_1_252/A sky130_fd_sc_hd__nor2_1_249/B
+ sky130_fd_sc_hd__fa_2_444/A sky130_fd_sc_hd__fa_2_444/B sky130_fd_sc_hd__ha_2_15/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_455 sky130_fd_sc_hd__fa_2_453/B sky130_fd_sc_hd__fa_2_459/B
+ sky130_fd_sc_hd__fa_2_455/A sky130_fd_sc_hd__fa_2_455/B sky130_fd_sc_hd__fa_2_455/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_466 sky130_fd_sc_hd__fa_2_464/CIN sky130_fd_sc_hd__fa_2_466/SUM
+ sky130_fd_sc_hd__fa_2_466/A sky130_fd_sc_hd__fa_2_466/B sky130_fd_sc_hd__fa_2_466/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_477 sky130_fd_sc_hd__or2_0_103/B sky130_fd_sc_hd__nor2_1_258/A
+ sky130_fd_sc_hd__fa_2_477/A sky130_fd_sc_hd__fa_2_477/B sky130_fd_sc_hd__nor2b_1_53/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_488 sky130_fd_sc_hd__nor2_1_263/B sky130_fd_sc_hd__or2_0_109/A
+ sky130_fd_sc_hd__fa_2_488/A sky130_fd_sc_hd__fa_2_488/B sky130_fd_sc_hd__nor2b_1_75/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor2_1_209 sky130_fd_sc_hd__nor2_1_209/B sky130_fd_sc_hd__nor2_1_209/Y
+ sky130_fd_sc_hd__nor2_1_209/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__and2_0_190 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_48/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_90/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_12_405 sky130_fd_sc_hd__buf_12_405/A sky130_fd_sc_hd__buf_12_476/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_416 sky130_fd_sc_hd__buf_12_66/X sky130_fd_sc_hd__buf_12_616/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_427 sky130_fd_sc_hd__buf_12_427/A sky130_fd_sc_hd__buf_12_534/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_438 sky130_fd_sc_hd__buf_12_438/A sky130_fd_sc_hd__buf_12_626/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_449 sky130_fd_sc_hd__buf_12_449/A sky130_fd_sc_hd__buf_12_641/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_605 sky130_fd_sc_hd__nand2_1_644/A sky130_fd_sc_hd__nor2_1_216/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_616 sky130_fd_sc_hd__nand2_1_633/A sky130_fd_sc_hd__nor2_1_212/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_627 sky130_fd_sc_hd__clkinv_1_627/Y sky130_fd_sc_hd__nand2_1_667/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_638 sky130_fd_sc_hd__nand2_1_688/A sky130_fd_sc_hd__nor2_1_227/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_649 sky130_fd_sc_hd__clkinv_1_649/Y sky130_fd_sc_hd__nand2_1_711/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_180 vssd1 vccd1 sky130_fd_sc_hd__inv_2_21/Y sky130_fd_sc_hd__nand2b_1_7/Y
+ sky130_fd_sc_hd__a222oi_1_59/Y sky130_fd_sc_hd__xor2_1_11/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_191 vssd1 vccd1 sky130_fd_sc_hd__inv_2_26/Y sky130_fd_sc_hd__nand2b_1_2/Y
+ sky130_fd_sc_hd__nand2_1_152/Y sky130_fd_sc_hd__ha_2_0/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_14 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_355/Q sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__o211ai_1_30/Y sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__a222oi_1_14/Y sky130_fd_sc_hd__dfxtp_1_306/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_601 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_25 vccd1 vssd1 sky130_fd_sc_hd__xnor2_1_187/Y sky130_fd_sc_hd__buf_2_17/X
+ sky130_fd_sc_hd__nor2_4_1/Y sky130_fd_sc_hd__xnor2_1_125/Y sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__a222oi_1_25/Y sky130_fd_sc_hd__xnor2_1_62/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_36 vccd1 vssd1 sky130_fd_sc_hd__xnor2_1_104/Y sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__xnor2_1_166/Y sky130_fd_sc_hd__xnor2_1_41/Y sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_36/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_612 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_623 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_47 vccd1 vssd1 sky130_fd_sc_hd__nor2_4_7/Y sky130_fd_sc_hd__xor2_2_1/X
+ sky130_fd_sc_hd__buf_6_3/X sky130_fd_sc_hd__nor2_4_1/Y sky130_fd_sc_hd__xor2_2_0/X
+ sky130_fd_sc_hd__a222oi_1_47/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_634 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_58 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__or2_0_9/B
+ sky130_fd_sc_hd__or2_0_9/A sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__or2_0_4/B
+ sky130_fd_sc_hd__a222oi_1_58/Y sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_69 vccd1 vssd1 sky130_fd_sc_hd__and3_4_6/X sky130_fd_sc_hd__buf_2_4/X
+ sky130_fd_sc_hd__buf_6_5/X sky130_fd_sc_hd__nor2_1_72/Y sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__a222oi_1_69/Y sky130_fd_sc_hd__nor2b_1_6/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_645 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_656 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_16 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_16/B sky130_fd_sc_hd__xnor2_1_16/Y
+ sky130_fd_sc_hd__xnor2_1_16/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_540 sky130_fd_sc_hd__nand2_1_540/Y sky130_fd_sc_hd__nand2_1_540/B
+ sky130_fd_sc_hd__nand2_1_546/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_667 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_27 vssd1 vccd1 sky130_fd_sc_hd__fa_2_97/A sky130_fd_sc_hd__and3_4_5/C
+ sky130_fd_sc_hd__xnor2_1_27/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_551 sky130_fd_sc_hd__or2_0_55/B sky130_fd_sc_hd__nor2_1_180/Y
+ sky130_fd_sc_hd__nor2_1_184/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_38 vssd1 vccd1 sky130_fd_sc_hd__fa_2_122/A sky130_fd_sc_hd__nor2_2_7/A
+ sky130_fd_sc_hd__xnor2_1_38/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_678 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_562 sky130_fd_sc_hd__nor2_1_182/A sky130_fd_sc_hd__or2_0_63/X
+ sky130_fd_sc_hd__or2_0_64/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_689 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_49 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_49/B sky130_fd_sc_hd__inv_2_17/A
+ sky130_fd_sc_hd__xnor2_1_49/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_573 sky130_fd_sc_hd__xnor2_1_156/A sky130_fd_sc_hd__nand2_1_574/Y
+ sky130_fd_sc_hd__or2_0_63/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_584 sky130_fd_sc_hd__nor2_1_188/A sky130_fd_sc_hd__nor2_1_189/Y
+ sky130_fd_sc_hd__nor2_1_192/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_595 sky130_fd_sc_hd__xnor2_1_165/A sky130_fd_sc_hd__nand2_1_596/Y
+ sky130_fd_sc_hd__nand2_1_595/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_1120 sky130_fd_sc_hd__clkinv_4_63/A sky130_fd_sc_hd__a22o_1_40/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1131 sky130_fd_sc_hd__clkinv_4_74/A sky130_fd_sc_hd__a22o_1_51/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1142 sky130_fd_sc_hd__buf_2_39/A sky130_fd_sc_hd__inv_4_16/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1600 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1611 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_2_5 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_5/Y sky130_fd_sc_hd__xnor2_2_5/A
+ sky130_fd_sc_hd__xnor2_2_5/B vssd1 vccd1 sky130_fd_sc_hd__xnor2_2
Xsky130_fd_sc_hd__decap_12_1622 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1633 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1644 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1655 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1666 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1677 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_380 sky130_fd_sc_hd__dfxtp_1_380/Q sky130_fd_sc_hd__dfxtp_1_380/CLK
+ sky130_fd_sc_hd__nor2b_1_103/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1688 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_0 sky130_fd_sc_hd__buf_2_27/A sky130_fd_sc_hd__nand2_1_0/B
+ sky130_fd_sc_hd__nand2_1_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_391 sky130_fd_sc_hd__dfxtp_1_391/Q sky130_fd_sc_hd__dfxtp_1_392/CLK
+ sky130_fd_sc_hd__nor2b_1_92/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1699 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__or4_1_2 sky130_fd_sc_hd__ha_2_3/A sky130_fd_sc_hd__ha_2_9/B sky130_fd_sc_hd__or4_1_2/X
+ sky130_fd_sc_hd__ha_2_5/A sky130_fd_sc_hd__ha_2_4/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__or4_1
Xsky130_fd_sc_hd__fa_2_230 sky130_fd_sc_hd__fa_2_226/B sky130_fd_sc_hd__fa_2_231/B
+ sky130_fd_sc_hd__fa_2_230/A sky130_fd_sc_hd__fa_2_230/B sky130_fd_sc_hd__xor2_1_331/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_241 sky130_fd_sc_hd__fa_2_238/CIN sky130_fd_sc_hd__fa_2_243/CIN
+ sky130_fd_sc_hd__fa_2_241/A sky130_fd_sc_hd__fa_2_241/B sky130_fd_sc_hd__xor2_1_347/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_252 sky130_fd_sc_hd__fa_2_248/A sky130_fd_sc_hd__fa_2_251/B
+ sky130_fd_sc_hd__fa_2_252/A sky130_fd_sc_hd__fa_2_252/B sky130_fd_sc_hd__fa_2_252/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_263 sky130_fd_sc_hd__nor2_1_142/A sky130_fd_sc_hd__nor2_1_145/B
+ sky130_fd_sc_hd__fa_2_263/A sky130_fd_sc_hd__fa_2_263/B sky130_fd_sc_hd__fa_2_263/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_274 sky130_fd_sc_hd__nor2_1_152/A sky130_fd_sc_hd__nor2_1_154/B
+ sky130_fd_sc_hd__fa_2_274/A sky130_fd_sc_hd__fa_2_274/B sky130_fd_sc_hd__xor2_1_400/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_285 sky130_fd_sc_hd__xor3_1_22/A sky130_fd_sc_hd__fa_2_286/B
+ sky130_fd_sc_hd__fa_2_285/A sky130_fd_sc_hd__fa_2_285/B sky130_fd_sc_hd__xor2_1_444/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_1 vccd1 vssd1 sky130_fd_sc_hd__and2_0_1/X la_data_out[36]
+ sky130_fd_sc_hd__nor2_2_0/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__fa_2_296 sky130_fd_sc_hd__fa_2_287/A sky130_fd_sc_hd__fa_2_297/B
+ sky130_fd_sc_hd__fa_2_296/A sky130_fd_sc_hd__fa_2_296/B sky130_fd_sc_hd__fa_2_296/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22oi_1_7 sky130_fd_sc_hd__nor2_4_0/Y sky130_fd_sc_hd__nor2_2_0/Y
+ sky130_fd_sc_hd__a22oi_1_7/B2 sky130_fd_sc_hd__or2_0_86/A sky130_fd_sc_hd__nand2_2_2/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_202 sky130_fd_sc_hd__buf_6_45/X sky130_fd_sc_hd__buf_12_413/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_213 sky130_fd_sc_hd__buf_6_53/X sky130_fd_sc_hd__buf_12_294/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_60 sky130_fd_sc_hd__nor2_1_96/Y sky130_fd_sc_hd__nand2_1_283/Y
+ sky130_fd_sc_hd__a21oi_1_60/Y sky130_fd_sc_hd__nand2_1_293/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_224 sky130_fd_sc_hd__buf_6_43/X sky130_fd_sc_hd__buf_12_445/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_71 sky130_fd_sc_hd__inv_2_42/A sky130_fd_sc_hd__o21ai_1_549/Y
+ sky130_fd_sc_hd__xnor2_2_0/A sky130_fd_sc_hd__nor2_1_132/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_235 sky130_fd_sc_hd__buf_6_71/X sky130_fd_sc_hd__buf_12_352/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_82 sky130_fd_sc_hd__o21ai_1_516/Y sky130_fd_sc_hd__nor2_1_122/A
+ sky130_fd_sc_hd__a21oi_1_82/Y sky130_fd_sc_hd__or2_0_47/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_246 sky130_fd_sc_hd__buf_6_30/X sky130_fd_sc_hd__buf_12_386/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_93 sky130_fd_sc_hd__nand2_1_443/Y sky130_fd_sc_hd__a21oi_1_93/B1
+ sky130_fd_sc_hd__a21oi_1_93/Y sky130_fd_sc_hd__nand2_1_444/A vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_1_105 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_181/Q sky130_fd_sc_hd__dfxtp_1_149/Q sky130_fd_sc_hd__o21ai_1_11/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_257 sky130_fd_sc_hd__buf_6_25/X sky130_fd_sc_hd__buf_12_427/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_116 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_170/Q sky130_fd_sc_hd__dfxtp_1_138/Q sky130_fd_sc_hd__o21ai_1_22/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_268 sky130_fd_sc_hd__buf_6_89/X sky130_fd_sc_hd__buf_12_563/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_127 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_161/Q sky130_fd_sc_hd__dfxtp_1_129/Q sky130_fd_sc_hd__o21ai_1_33/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_279 sky130_fd_sc_hd__buf_12_279/A sky130_fd_sc_hd__buf_12_509/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_138 sky130_fd_sc_hd__xnor2_1_78/Y sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xnor2_1_15/Y sky130_fd_sc_hd__o21ai_1_56/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_149 sky130_fd_sc_hd__xor2_1_313/X sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xor2_1_100/X sky130_fd_sc_hd__o21ai_1_77/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_402 sky130_fd_sc_hd__xnor2_1_3/A sky130_fd_sc_hd__nand2_1_312/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_413 sky130_fd_sc_hd__a21oi_1_85/B1 sky130_fd_sc_hd__nand2_1_420/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_424 sky130_fd_sc_hd__nor2_1_111/A sky130_fd_sc_hd__nand2_1_360/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_435 sky130_fd_sc_hd__o21ai_1_472/A2 sky130_fd_sc_hd__xnor2_1_79/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_446 sky130_fd_sc_hd__nand2_1_374/A sky130_fd_sc_hd__or2_0_32/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_457 sky130_fd_sc_hd__a21oi_1_70/B1 sky130_fd_sc_hd__nand2_1_394/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_468 sky130_fd_sc_hd__nor2_1_134/B sky130_fd_sc_hd__nor2_1_136/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_479 sky130_fd_sc_hd__nand2_1_434/A sky130_fd_sc_hd__nor2_1_144/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a222oi_1_2 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_343/Q sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__o211ai_1_18/Y sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__a222oi_1_2/Y sky130_fd_sc_hd__dfxtp_1_294/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_420 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_431 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_442 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_453 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_464 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_475 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_486 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_370 sky130_fd_sc_hd__xnor2_1_80/A sky130_fd_sc_hd__nand2_1_371/Y
+ sky130_fd_sc_hd__nand2_1_370/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_497 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_381 sky130_fd_sc_hd__xnor2_1_85/A sky130_fd_sc_hd__nand2_1_382/Y
+ sky130_fd_sc_hd__or2_0_41/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_980 sky130_fd_sc_hd__buf_2_167/A sky130_fd_sc_hd__clkinv_2_33/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xor2_1_209 sky130_fd_sc_hd__o21a_1_1/A1 sky130_fd_sc_hd__xor2_1_209/X
+ sky130_fd_sc_hd__xor2_1_209/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_392 sky130_fd_sc_hd__nand2_1_392/Y sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__buf_4_4/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_991 sky130_fd_sc_hd__clkinv_1_991/Y sky130_fd_sc_hd__inv_2_156/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1430 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1441 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1452 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1463 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1474 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_905 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_266/Y sky130_fd_sc_hd__xor2_1_688/B
+ sky130_fd_sc_hd__nand2_1_841/Y sky130_fd_sc_hd__xnor2_1_302/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1485 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_916 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_279/Y la_data_out[42]
+ sky130_fd_sc_hd__a21oi_1_190/Y sky130_fd_sc_hd__o21ai_1_916/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1496 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_9 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__buf_2_14 vccd1 vssd1 sky130_fd_sc_hd__or2_0_71/B sky130_fd_sc_hd__buf_2_14/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_25 vccd1 vssd1 sky130_fd_sc_hd__or2_0_72/A sky130_fd_sc_hd__buf_2_25/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_36 vccd1 vssd1 sky130_fd_sc_hd__buf_2_36/X sky130_fd_sc_hd__buf_2_36/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_47 vccd1 vssd1 sky130_fd_sc_hd__buf_2_47/X sky130_fd_sc_hd__buf_2_47/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_58 vccd1 vssd1 sky130_fd_sc_hd__buf_8_94/A sky130_fd_sc_hd__buf_8_3/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_69 vccd1 vssd1 sky130_fd_sc_hd__buf_2_69/X sky130_fd_sc_hd__buf_2_69/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o211ai_1_30 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_35/B1
+ sky130_fd_sc_hd__o211ai_1_30/Y sky130_fd_sc_hd__a22oi_1_92/Y sky130_fd_sc_hd__a22oi_1_93/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_41 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o22ai_1_22/B1
+ sky130_fd_sc_hd__fa_2_354/A sky130_fd_sc_hd__nand2_1_61/Y sky130_fd_sc_hd__a21oi_1_12/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_52 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o22ai_1_11/B1
+ sky130_fd_sc_hd__fa_2_401/A sky130_fd_sc_hd__nand2_1_72/Y sky130_fd_sc_hd__a21oi_1_23/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_63 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o22ai_1_2/B1
+ sky130_fd_sc_hd__nor2_1_219/A sky130_fd_sc_hd__nand2_1_83/Y sky130_fd_sc_hd__a21oi_1_34/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__diode_2_9 sky130_fd_sc_hd__conb_1_147/HI vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkinv_1_210 sky130_fd_sc_hd__o22ai_1_12/B1 sky130_fd_sc_hd__dfxtp_1_107/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_221 sky130_fd_sc_hd__nor2_1_12/A sky130_fd_sc_hd__dfxtp_1_135/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_232 sky130_fd_sc_hd__o22ai_1_4/A2 sky130_fd_sc_hd__dfxtp_1_163/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_243 sky130_fd_sc_hd__o22ai_1_1/B1 sky130_fd_sc_hd__dfxtp_1_96/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_254 sky130_fd_sc_hd__o21ai_1_105/A2 sky130_fd_sc_hd__xnor2_1_161/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_265 sky130_fd_sc_hd__o21ai_1_149/A2 sky130_fd_sc_hd__xnor2_1_185/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_276 sky130_fd_sc_hd__and2_0_131/A sky130_fd_sc_hd__a222oi_1_20/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_287 sky130_fd_sc_hd__and2_0_196/A sky130_fd_sc_hd__a222oi_1_31/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_298 sky130_fd_sc_hd__and2_0_231/A sky130_fd_sc_hd__a222oi_1_42/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xor3_1_5 sky130_fd_sc_hd__xor3_1_5/X sky130_fd_sc_hd__xor3_1_5/C
+ sky130_fd_sc_hd__xor3_1_5/B sky130_fd_sc_hd__xor3_1_5/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__a21oi_1_6 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_35/Y
+ sky130_fd_sc_hd__a21oi_1_6/Y sky130_fd_sc_hd__dfxtp_1_93/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__and3_4_12 sky130_fd_sc_hd__nor2_4_14/B sky130_fd_sc_hd__nor2_4_14/A
+ sky130_fd_sc_hd__and3_4_12/C sky130_fd_sc_hd__and3_4_12/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__clkbuf_4_19 sky130_fd_sc_hd__clkbuf_4_19/X sky130_fd_sc_hd__buf_6_8/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and3_4_23 sky130_fd_sc_hd__and3_4_23/A sky130_fd_sc_hd__and3_4_23/B
+ sky130_fd_sc_hd__and3_4_23/C sky130_fd_sc_hd__and3_4_23/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__a21oi_1_140 sky130_fd_sc_hd__xnor2_1_190/B sky130_fd_sc_hd__clkinv_1_629/Y
+ sky130_fd_sc_hd__xor2_1_641/A sky130_fd_sc_hd__or2_0_75/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_151 sky130_fd_sc_hd__or2_0_87/X sky130_fd_sc_hd__clkinv_1_662/Y
+ sky130_fd_sc_hd__a21oi_1_151/Y sky130_fd_sc_hd__clkinv_1_663/Y vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_162 sky130_fd_sc_hd__xnor2_1_215/B sky130_fd_sc_hd__clkinv_1_695/Y
+ sky130_fd_sc_hd__xor2_1_663/A sky130_fd_sc_hd__or2_0_93/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_173 sky130_fd_sc_hd__xnor2_1_294/B sky130_fd_sc_hd__clkinv_1_814/Y
+ sky130_fd_sc_hd__xor2_1_679/A sky130_fd_sc_hd__or2_0_103/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_184 sky130_fd_sc_hd__buf_6_91/X sky130_fd_sc_hd__nor2_1_267/Y
+ sky130_fd_sc_hd__a21oi_1_184/Y sky130_fd_sc_hd__nand3_1_5/C vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_195 sky130_fd_sc_hd__nor4b_1_0/D_N sky130_fd_sc_hd__maj3_1_2/X
+ sky130_fd_sc_hd__a21oi_1_195/Y sky130_fd_sc_hd__o211ai_1_65/Y vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_103 sky130_fd_sc_hd__inv_2_171/Y sky130_fd_sc_hd__buf_4_30/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_114 sky130_fd_sc_hd__buf_8_114/A sky130_fd_sc_hd__buf_6_75/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_125 sky130_fd_sc_hd__inv_4_9/Y sky130_fd_sc_hd__buf_6_76/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_136 sky130_fd_sc_hd__inv_2_84/Y sky130_fd_sc_hd__buf_8_136/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_147 sky130_fd_sc_hd__inv_2_121/Y sky130_fd_sc_hd__buf_8_161/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nor2_4_9 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__nor2_4_9/A
+ sky130_fd_sc_hd__nor2_4_9/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__buf_8_158 sky130_fd_sc_hd__buf_6_21/X sky130_fd_sc_hd__buf_6_89/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__decap_12_250 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_261 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_272 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_283 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_294 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1260 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1271 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_702 vssd1 vccd1 sky130_fd_sc_hd__inv_2_49/Y sky130_fd_sc_hd__nand2b_1_21/Y
+ sky130_fd_sc_hd__o21ai_1_702/B1 sky130_fd_sc_hd__xor2_1_481/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1282 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_713 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_713/A2 sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_713/B1 sky130_fd_sc_hd__xor2_1_491/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1293 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_724 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_10/X sky130_fd_sc_hd__nand2_1_546/Y
+ sky130_fd_sc_hd__a21oi_1_115/Y sky130_fd_sc_hd__xnor2_1_146/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_735 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_181/Y sky130_fd_sc_hd__nor2_1_180/A
+ sky130_fd_sc_hd__nor2_1_179/Y sky130_fd_sc_hd__o21ai_1_735/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_746 vssd1 vccd1 sky130_fd_sc_hd__nand2_2_13/Y sky130_fd_sc_hd__nand2b_1_20/Y
+ sky130_fd_sc_hd__a22oi_1_216/Y sky130_fd_sc_hd__xor2_1_521/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_757 vssd1 vccd1 sky130_fd_sc_hd__inv_2_51/Y sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__o21ai_1_757/B1 sky130_fd_sc_hd__xor2_1_532/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_768 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_10/X sky130_fd_sc_hd__nand2_1_567/Y
+ sky130_fd_sc_hd__a21oi_1_118/Y sky130_fd_sc_hd__xnor2_1_155/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_779 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_3/Y sky130_fd_sc_hd__nand2b_2_6/Y
+ sky130_fd_sc_hd__o21ai_1_779/B1 sky130_fd_sc_hd__xor2_1_553/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_20 sky130_fd_sc_hd__fa_2_97/A sky130_fd_sc_hd__fa_2_3/A sky130_fd_sc_hd__xor2_1_20/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_31 sky130_fd_sc_hd__xor2_1_6/B sky130_fd_sc_hd__fa_2_13/A
+ sky130_fd_sc_hd__xor2_1_31/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_42 sky130_fd_sc_hd__xor2_1_42/B sky130_fd_sc_hd__xor2_1_42/X
+ sky130_fd_sc_hd__xor2_1_42/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_53 sky130_fd_sc_hd__fa_2_97/A sky130_fd_sc_hd__fa_2_31/A
+ sky130_fd_sc_hd__xor2_1_53/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_64 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__fa_2_46/B
+ sky130_fd_sc_hd__xor2_1_64/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_75 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__xor2_1_75/X
+ sky130_fd_sc_hd__xor2_1_75/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_86 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__xor2_1_86/X
+ sky130_fd_sc_hd__xor2_1_86/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_97 sky130_fd_sc_hd__xor2_1_9/B sky130_fd_sc_hd__xor2_1_97/X
+ sky130_fd_sc_hd__xor2_1_97/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2b_1_3 sky130_fd_sc_hd__nand2b_1_3/Y sky130_fd_sc_hd__and3_1_0/C
+ sky130_fd_sc_hd__and3_1_0/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__o21ai_2_18 sky130_fd_sc_hd__a31oi_1_1/Y sky130_fd_sc_hd__o21ai_2_18/Y
+ sky130_fd_sc_hd__o21ai_2_18/A2 sky130_fd_sc_hd__o21ai_2_18/A1 vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__o21ai_2
Xsky130_fd_sc_hd__xor2_1_540 sky130_fd_sc_hd__fa_2_379/A sky130_fd_sc_hd__xor2_1_540/X
+ sky130_fd_sc_hd__xor2_1_540/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_551 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__xor2_1_551/X
+ sky130_fd_sc_hd__xor2_1_551/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_562 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__fa_2_380/A
+ sky130_fd_sc_hd__xor2_1_562/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_573 sky130_fd_sc_hd__fah_1_14/A sky130_fd_sc_hd__fa_2_391/B
+ sky130_fd_sc_hd__xor2_1_573/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_584 sky130_fd_sc_hd__fah_1_14/A sky130_fd_sc_hd__xor2_1_584/X
+ sky130_fd_sc_hd__xor2_1_584/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_595 sky130_fd_sc_hd__fah_1_14/A sky130_fd_sc_hd__fah_1_14/CI
+ sky130_fd_sc_hd__xor2_1_595/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a221oi_1_1 sky130_fd_sc_hd__nand4_1_1/B sky130_fd_sc_hd__o22ai_1_137/Y
+ sky130_fd_sc_hd__o31ai_2_0/A2 sky130_fd_sc_hd__nor2_4_19/B sky130_fd_sc_hd__nand4_1_0/C
+ sky130_fd_sc_hd__dfxtp_1_363/Q vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__a221oi_1
Xsky130_fd_sc_hd__a222oi_1_604 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_394/Q sky130_fd_sc_hd__and2b_4_13/X
+ sky130_fd_sc_hd__nor2_4_19/Y sky130_fd_sc_hd__dfxtp_1_458/Q sky130_fd_sc_hd__nor2_4_19/B
+ sky130_fd_sc_hd__clkinv_1_801/A sky130_fd_sc_hd__dfxtp_1_426/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__and2_0_14 vccd1 vssd1 sky130_fd_sc_hd__and2_0_14/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_14/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_25 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_2_6/D sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__and2_0_25/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_36 vccd1 vssd1 sky130_fd_sc_hd__and2_0_36/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__nor2_1_73/B vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_47 vccd1 vssd1 sky130_fd_sc_hd__and2_0_47/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__nor2_1_85/B vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_58 vccd1 vssd1 sky130_fd_sc_hd__and2_0_58/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__or2_0_4/B vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_69 vccd1 vssd1 sky130_fd_sc_hd__and2_0_69/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__or2_0_66/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nor2_2_6 sky130_fd_sc_hd__inv_6_0/Y sky130_fd_sc_hd__nor2_2_6/Y
+ sky130_fd_sc_hd__buf_8_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__buf_8_13 sky130_fd_sc_hd__inv_2_93/Y sky130_fd_sc_hd__buf_8_13/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_24 sky130_fd_sc_hd__buf_8_24/A sky130_fd_sc_hd__buf_8_24/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_35 sky130_fd_sc_hd__buf_8_35/A sky130_fd_sc_hd__buf_8_35/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_46 sky130_fd_sc_hd__buf_8_46/A sky130_fd_sc_hd__buf_8_46/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_57 sky130_fd_sc_hd__buf_8_57/A sky130_fd_sc_hd__buf_8_57/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xnor2_1_170 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_170/B sky130_fd_sc_hd__inv_2_45/A
+ sky130_fd_sc_hd__xnor2_1_170/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__buf_8_68 sky130_fd_sc_hd__inv_4_14/Y sky130_fd_sc_hd__buf_8_68/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xnor2_1_181 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_181/B sky130_fd_sc_hd__inv_2_48/A
+ sky130_fd_sc_hd__xnor2_1_181/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__buf_8_79 sky130_fd_sc_hd__buf_8_79/A sky130_fd_sc_hd__buf_8_79/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xnor2_1_192 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_192/B sky130_fd_sc_hd__and2_0_269/A
+ sky130_fd_sc_hd__xnor2_1_192/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__dfxtp_1_209 sky130_fd_sc_hd__fa_2_357/A sky130_fd_sc_hd__dfxtp_2_0/CLK
+ sky130_fd_sc_hd__and2_0_60/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_510 vssd1 vccd1 sky130_fd_sc_hd__inv_2_33/Y sky130_fd_sc_hd__nand2b_2_3/Y
+ sky130_fd_sc_hd__o21ai_1_510/B1 sky130_fd_sc_hd__xor2_1_309/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1090 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_521 vssd1 vccd1 sky130_fd_sc_hd__buf_2_11/X sky130_fd_sc_hd__nand2b_1_8/Y
+ sky130_fd_sc_hd__o21ai_1_521/B1 sky130_fd_sc_hd__xor2_1_320/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_532 vssd1 vccd1 sky130_fd_sc_hd__inv_2_36/Y sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_532/B1 sky130_fd_sc_hd__xor2_1_331/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_543 vssd1 vccd1 sky130_fd_sc_hd__inv_2_40/Y sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_543/B1 sky130_fd_sc_hd__xor2_1_341/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_554 vssd1 vccd1 sky130_fd_sc_hd__inv_2_29/Y sky130_fd_sc_hd__nand2b_1_9/Y
+ sky130_fd_sc_hd__o21ai_1_554/B1 sky130_fd_sc_hd__xor2_1_352/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_565 vssd1 vccd1 sky130_fd_sc_hd__inv_2_32/Y sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_565/B1 sky130_fd_sc_hd__xor2_1_363/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_576 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_145/Y sky130_fd_sc_hd__nand2_1_442/Y
+ sky130_fd_sc_hd__nand2_1_437/Y sky130_fd_sc_hd__o21ai_1_576/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_587 vssd1 vccd1 sky130_fd_sc_hd__buf_2_9/X sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_587/B1 sky130_fd_sc_hd__xor2_1_380/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_598 vssd1 vccd1 sky130_fd_sc_hd__nand2_2_12/Y sky130_fd_sc_hd__nand2b_2_3/Y
+ sky130_fd_sc_hd__a22oi_1_208/Y sky130_fd_sc_hd__xor2_1_392/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__buf_2_109 vccd1 vssd1 sky130_fd_sc_hd__buf_2_109/X sky130_fd_sc_hd__buf_2_109/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__xor2_1_370 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__fah_1_5/CI
+ sky130_fd_sc_hd__xor2_1_370/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_381 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__fa_2_260/B
+ sky130_fd_sc_hd__xor2_1_381/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_392 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__fa_2_267/B
+ sky130_fd_sc_hd__xor2_1_392/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__ha_2_9 vssd1 vccd1 sky130_fd_sc_hd__ha_2_9/A sky130_fd_sc_hd__ha_2_8/B
+ sky130_fd_sc_hd__ha_2_9/SUM sky130_fd_sc_hd__ha_2_9/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_330 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1_2/D sky130_fd_sc_hd__buf_2_175/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_401 vccd1 vssd1 sky130_fd_sc_hd__and3_4_23/X sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__buf_6_2/X sky130_fd_sc_hd__nor2_1_178/Y sky130_fd_sc_hd__buf_4_7/X
+ sky130_fd_sc_hd__o21ai_1_667/B1 sky130_fd_sc_hd__nor2b_1_15/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_341 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1_17/D sky130_fd_sc_hd__dfxtp_1_18/Q
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_412 vccd1 vssd1 sky130_fd_sc_hd__and3_4_20/X sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__buf_4_3/X sky130_fd_sc_hd__nor2_4_16/Y sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__o21ai_1_682/B1 sky130_fd_sc_hd__and2b_4_11/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_352 vssd1 vccd1 sky130_fd_sc_hd__inv_2_1/A sky130_fd_sc_hd__a222oi_1_4/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_423 vccd1 vssd1 sky130_fd_sc_hd__and3_4_26/X sky130_fd_sc_hd__buf_2_20/X
+ sky130_fd_sc_hd__buf_2_21/X sky130_fd_sc_hd__nor2_2_31/Y sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__o21ai_1_697/B1 sky130_fd_sc_hd__nor2b_1_12/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_434 vccd1 vssd1 sky130_fd_sc_hd__and3_4_21/X sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__buf_4_2/X sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__o21ai_1_708/B1 sky130_fd_sc_hd__and2b_4_12/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_445 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__or2_0_60/B sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__or2_0_60/A
+ sky130_fd_sc_hd__o21ai_1_723/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_456 vccd1 vssd1 sky130_fd_sc_hd__and3_4_20/X sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__nor2_1_85/B sky130_fd_sc_hd__nor2_4_16/Y sky130_fd_sc_hd__nor2_2_10/B
+ sky130_fd_sc_hd__o21ai_1_738/B1 sky130_fd_sc_hd__and2b_4_11/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_467 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__buf_4_4/X sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__o21ai_1_751/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_478 vccd1 vssd1 sky130_fd_sc_hd__and3_4_25/X sky130_fd_sc_hd__or2_0_72/B
+ sky130_fd_sc_hd__or2_0_72/A sky130_fd_sc_hd__nor2_1_186/Y sky130_fd_sc_hd__or2_0_71/B
+ sky130_fd_sc_hd__o21ai_1_765/B1 sky130_fd_sc_hd__nor2b_1_17/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_489 vccd1 vssd1 sky130_fd_sc_hd__and3_4_20/X sky130_fd_sc_hd__buf_2_27/X
+ sky130_fd_sc_hd__buf_2_15/X sky130_fd_sc_hd__nor2_4_16/Y sky130_fd_sc_hd__buf_2_4/A
+ sky130_fd_sc_hd__o21ai_1_779/B1 sky130_fd_sc_hd__and2b_4_11/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__and2_0_350 vccd1 vssd1 sky130_fd_sc_hd__and2_0_350/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__buf_2_188/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_361 vccd1 vssd1 sky130_fd_sc_hd__and2_0_361/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__and2_0_361/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_372 vccd1 vssd1 sky130_fd_sc_hd__and2_0_372/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_65/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_383 vccd1 vssd1 sky130_fd_sc_hd__and2_0_383/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_80/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_394 vccd1 vssd1 sky130_fd_sc_hd__and2_0_394/X sky130_fd_sc_hd__and2_0_401/B
+ sky130_fd_sc_hd__and2_0_394/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__conb_1_3 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__conb_1_3/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__inv_2_150 sky130_fd_sc_hd__inv_2_150/A sky130_fd_sc_hd__inv_2_150/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_12_9 sky130_fd_sc_hd__buf_12_9/A sky130_fd_sc_hd__buf_12_9/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_609 sky130_fd_sc_hd__buf_12_609/A sky130_fd_sc_hd__buf_12_609/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__inv_2_161 sky130_fd_sc_hd__inv_2_81/Y sky130_fd_sc_hd__inv_2_161/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_172 sky130_fd_sc_hd__inv_2_172/A sky130_fd_sc_hd__inv_2_173/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_183 sky130_fd_sc_hd__inv_2_183/A sky130_fd_sc_hd__inv_2_183/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_194 sky130_fd_sc_hd__nand2_1_8/B sky130_fd_sc_hd__nand2_1_7/B
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__o22ai_1_102 sky130_fd_sc_hd__xnor2_2_4/Y sky130_fd_sc_hd__xnor2_1_251/Y
+ sky130_fd_sc_hd__fa_2_444/A sky130_fd_sc_hd__xnor2_1_252/Y sky130_fd_sc_hd__o22ai_1_96/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_113 sky130_fd_sc_hd__xnor2_1_274/Y sky130_fd_sc_hd__xnor2_1_260/Y
+ sky130_fd_sc_hd__ha_2_16/A sky130_fd_sc_hd__inv_2_65/Y sky130_fd_sc_hd__o22ai_1_99/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_124 sky130_fd_sc_hd__xnor2_1_272/Y sky130_fd_sc_hd__xnor2_1_271/Y
+ sky130_fd_sc_hd__fa_2_455/A sky130_fd_sc_hd__nor2b_1_24/A sky130_fd_sc_hd__nand2_1_722/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_135 sky130_fd_sc_hd__a221o_1_0/A2 sky130_fd_sc_hd__a221o_1_0/B2
+ sky130_fd_sc_hd__a221o_1_0/C1 sky130_fd_sc_hd__a221o_1_0/A1 sky130_fd_sc_hd__a221o_1_0/B1
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_809 sky130_fd_sc_hd__nand2_1_796/A sky130_fd_sc_hd__nor2_1_255/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_2_13 sky130_fd_sc_hd__nor2_2_13/B sky130_fd_sc_hd__nor2_2_13/Y
+ sky130_fd_sc_hd__nor2_2_13/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__nor2_2_24 sky130_fd_sc_hd__nor2_2_24/B sky130_fd_sc_hd__nor2_2_24/Y
+ sky130_fd_sc_hd__nor2_2_24/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__o211ai_1_3 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_3/A2
+ sky130_fd_sc_hd__o211ai_1_3/Y sky130_fd_sc_hd__a22oi_1_38/Y sky130_fd_sc_hd__a22oi_1_39/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__a31oi_1_0 vssd1 vccd1 sky130_fd_sc_hd__a31oi_1_0/Y sky130_fd_sc_hd__a31oi_1_0/B1
+ sky130_fd_sc_hd__o31ai_1_1/A1 sky130_fd_sc_hd__nor2_1_273/A sky130_fd_sc_hd__a31oi_1_0/A3
+ vssd1 vccd1 sky130_fd_sc_hd__a31oi_1
Xsky130_fd_sc_hd__o21ai_1_340 vssd1 vccd1 sky130_fd_sc_hd__inv_2_16/Y sky130_fd_sc_hd__nand2b_2_0/Y
+ sky130_fd_sc_hd__o21ai_1_340/B1 sky130_fd_sc_hd__xor2_1_159/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_351 vssd1 vccd1 sky130_fd_sc_hd__buf_2_1/X sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__o21ai_1_351/B1 sky130_fd_sc_hd__xor2_1_166/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_362 vssd1 vccd1 sky130_fd_sc_hd__inv_2_15/Y sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__o21ai_1_362/B1 sky130_fd_sc_hd__xor2_1_178/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_373 vssd1 vccd1 sky130_fd_sc_hd__inv_2_18/Y sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__o21ai_1_373/B1 sky130_fd_sc_hd__xor2_1_188/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_384 vssd1 vccd1 sky130_fd_sc_hd__buf_2_2/X sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__o21ai_1_384/B1 sky130_fd_sc_hd__xor2_1_200/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_395 vssd1 vccd1 sky130_fd_sc_hd__a21oi_2_7/Y sky130_fd_sc_hd__nor2_1_110/Y
+ sky130_fd_sc_hd__nand2_1_345/Y sky130_fd_sc_hd__xnor2_2_1/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_805 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_816 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_700 sky130_fd_sc_hd__xor2_1_649/B sky130_fd_sc_hd__nand2_1_701/Y
+ sky130_fd_sc_hd__nand2_1_700/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_827 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_711 sky130_fd_sc_hd__nand2_1_711/Y sky130_fd_sc_hd__or2_0_83/A
+ la_data_out[67] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_838 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_722 sky130_fd_sc_hd__nand2_1_722/Y sky130_fd_sc_hd__nor2b_1_24/A
+ sky130_fd_sc_hd__xor2_1_673/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_849 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__mux2_2_20 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_20/A1 sky130_fd_sc_hd__buf_2_78/X
+ sky130_fd_sc_hd__mux2_8_0/S sky130_fd_sc_hd__mux2_2_20/X vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_733 sky130_fd_sc_hd__nand2_1_733/Y sky130_fd_sc_hd__nor2_1_237/A
+ sky130_fd_sc_hd__nor2_1_237/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_31 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_31/A1 sky130_fd_sc_hd__buf_6_13/X
+ sky130_fd_sc_hd__mux2_8_1/S sky130_fd_sc_hd__mux2_2_31/X vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_744 sky130_fd_sc_hd__nand2_1_744/Y sky130_fd_sc_hd__nor2_1_239/A
+ sky130_fd_sc_hd__xor2_1_664/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_42 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_42/A1 sky130_fd_sc_hd__buf_2_93/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__mux2_2_42/X vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_755 sky130_fd_sc_hd__xor2_1_659/B sky130_fd_sc_hd__nand2_1_770/Y
+ sky130_fd_sc_hd__nand2_1_755/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_53 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_53/A1 sky130_fd_sc_hd__buf_4_17/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__or2_0_82/A vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_766 sky130_fd_sc_hd__xnor2_1_217/A sky130_fd_sc_hd__nand2_1_783/Y
+ sky130_fd_sc_hd__or2_0_96/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_777 sky130_fd_sc_hd__nand2_1_777/Y sky130_fd_sc_hd__or2_0_94/A
+ sky130_fd_sc_hd__or2_0_94/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_788 sky130_fd_sc_hd__inv_2_68/A sky130_fd_sc_hd__ha_2_9/B
+ sky130_fd_sc_hd__o31ai_2_0/A2 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_799 sky130_fd_sc_hd__nand2_1_799/Y sky130_fd_sc_hd__or2_0_101/A
+ sky130_fd_sc_hd__or2_0_101/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_1804 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1815 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1826 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1837 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_540 wbs_dat_o[19] sky130_fd_sc_hd__dfxtp_1_544/CLK sky130_fd_sc_hd__nor2b_1_138/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1848 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_551 wbs_dat_o[30] sky130_fd_sc_hd__dfxtp_1_552/CLK sky130_fd_sc_hd__nor2b_1_127/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1859 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_sram_1kbyte_1rw1r_32x256_8_11 sky130_fd_sc_hd__clkbuf_1_249/X sky130_fd_sc_hd__clkbuf_1_249/X
+ sky130_fd_sc_hd__buf_12_543/X sky130_fd_sc_hd__buf_12_626/X sky130_fd_sc_hd__buf_12_561/X
+ sky130_fd_sc_hd__buf_12_546/X sky130_fd_sc_hd__buf_12_444/X sky130_fd_sc_hd__buf_12_615/X
+ sky130_fd_sc_hd__buf_12_658/X sky130_fd_sc_hd__clkinv_1_954/Y sky130_fd_sc_hd__buf_12_537/X
+ sky130_fd_sc_hd__buf_12_599/X sky130_fd_sc_hd__buf_12_577/X vccd1 sky130_fd_sc_hd__clkinv_8_28/Y
+ sky130_fd_sc_hd__buf_2_144/A sky130_fd_sc_hd__buf_2_154/A sky130_fd_sc_hd__buf_2_82/A
+ sky130_fd_sc_hd__buf_2_81/A sky130_fd_sc_hd__buf_2_80/A sky130_fd_sc_hd__buf_2_79/A
+ sky130_fd_sc_hd__buf_2_78/A sky130_fd_sc_hd__buf_2_77/A sky130_fd_sc_hd__buf_2_76/A
+ sky130_fd_sc_hd__buf_2_75/A sky130_fd_sc_hd__buf_2_74/A sky130_fd_sc_hd__buf_2_73/A
+ sky130_fd_sc_hd__buf_2_72/A sky130_fd_sc_hd__buf_2_71/A sky130_fd_sc_hd__buf_2_70/A
+ sky130_fd_sc_hd__buf_2_69/A sky130_fd_sc_hd__buf_12_562/X sky130_fd_sc_hd__buf_8_1/A
+ sky130_fd_sc_hd__inv_4_12/A sky130_fd_sc_hd__buf_6_12/A sky130_fd_sc_hd__buf_4_12/A
+ sky130_fd_sc_hd__buf_4_10/A sky130_fd_sc_hd__buf_4_9/A sky130_fd_sc_hd__buf_6_16/A
+ sky130_fd_sc_hd__buf_4_14/A sky130_fd_sc_hd__buf_6_15/A sky130_fd_sc_hd__buf_6_13/A
+ sky130_fd_sc_hd__buf_4_20/A sky130_fd_sc_hd__buf_4_22/A sky130_fd_sc_hd__buf_4_23/A
+ sky130_fd_sc_hd__buf_2_146/A sky130_fd_sc_hd__buf_2_145/A sky130_fd_sc_hd__buf_6_14/A
+ sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[10] sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[11]
+ sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[12] sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[13]
+ sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[14] sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[15]
+ sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[16] sky130_fd_sc_hd__buf_12_608/X sky130_fd_sc_hd__buf_12_155/X
+ sky130_fd_sc_hd__buf_12_123/X sky130_fd_sc_hd__buf_12_15/X sky130_fd_sc_hd__buf_12_139/X
+ sky130_fd_sc_hd__clkinv_8_75/Y sky130_fd_sc_hd__buf_4_40/X sky130_fd_sc_hd__inv_2_108/A
+ sky130_fd_sc_hd__clkinv_1_914/Y sky130_fd_sc_hd__clkinv_1_912/Y sky130_fd_sc_hd__clkinv_1_910/Y
+ sky130_fd_sc_hd__buf_6_93/X sky130_fd_sc_hd__clkinv_1_905/Y sky130_fd_sc_hd__clkbuf_1_278/X
+ sky130_fd_sc_hd__clkinv_1_898/Y sky130_fd_sc_hd__clkinv_1_895/Y sky130_fd_sc_hd__clkbuf_1_42/X
+ sky130_fd_sc_hd__clkinv_1_890/Y sky130_fd_sc_hd__clkinv_1_889/Y sky130_fd_sc_hd__clkinv_1_888/Y
+ sky130_fd_sc_hd__clkinv_1_887/Y sky130_fd_sc_hd__clkinv_1_886/Y sky130_fd_sc_hd__clkinv_1_883/Y
+ sky130_fd_sc_hd__clkinv_1_881/Y sky130_fd_sc_hd__clkinv_1_880/Y sky130_fd_sc_hd__clkinv_1_879/Y
+ sky130_fd_sc_hd__clkinv_1_876/Y wbs_dat_i[21] sky130_fd_sc_hd__buf_2_37/A sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[0]
+ sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[1] sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[2]
+ sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[3] sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[4]
+ sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[5] sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[6]
+ sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[7] sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[8]
+ sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[9] sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[25]
+ sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[26] sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[27]
+ sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[28] sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[29]
+ sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[30] sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[31]
+ sky130_fd_sc_hd__clkinv_1_845/Y sky130_fd_sc_hd__clkinv_1_869/Y sky130_fd_sc_hd__clkinv_1_867/Y
+ sky130_fd_sc_hd__clkinv_1_865/Y sky130_fd_sc_hd__clkinv_1_863/Y sky130_fd_sc_hd__clkinv_1_860/Y
+ sky130_fd_sc_hd__clkinv_1_857/Y sky130_fd_sc_hd__clkinv_1_853/Y sky130_fd_sc_hd__clkinv_1_849/Y
+ sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[17] sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[18]
+ sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[19] sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[20]
+ sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[21] sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[22]
+ sky130_fd_sc_hd__buf_12_552/X sky130_fd_sc_hd__buf_12_516/X sky130_fd_sc_hd__buf_12_532/X
+ sky130_fd_sc_hd__buf_12_665/X sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[23] sky130_sram_1kbyte_1rw1r_32x256_8_11/dout0[24]
+ sky130_sram_1kbyte_1rw1r_32x256_8_11/sky130_sram_1kbyte_1rw1r_32x256_8_bank_0/sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0/gnd_uq26
+ vssd1 sky130_sram_1kbyte_1rw1r_32x256_8
Xsky130_fd_sc_hd__a222oi_1_220 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__or2_0_42/B
+ sky130_fd_sc_hd__or2_0_39/B sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__or2_0_58/A
+ sky130_fd_sc_hd__o21ai_1_409/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_160 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_160/X sky130_fd_sc_hd__inv_12_0/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_231 vccd1 vssd1 sky130_fd_sc_hd__and3_4_10/X sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__buf_4_4/X sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__o21ai_1_424/B1 sky130_fd_sc_hd__and2b_4_7/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_171 vssd1 vccd1 sky130_fd_sc_hd__a22o_1_32/B2 sky130_fd_sc_hd__clkbuf_1_171/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_242 vccd1 vssd1 sky130_fd_sc_hd__and3_4_14/X sky130_fd_sc_hd__buf_4_0/X
+ sky130_fd_sc_hd__buf_2_23/X sky130_fd_sc_hd__nor2_1_127/Y sky130_fd_sc_hd__buf_2_31/X
+ sky130_fd_sc_hd__o21ai_1_438/B1 sky130_fd_sc_hd__nor2b_1_10/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_182 vssd1 vccd1 sky130_fd_sc_hd__a22o_1_22/B2 sky130_fd_sc_hd__clkbuf_1_182/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_253 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__or2_0_60/B sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__or2_0_60/A
+ sky130_fd_sc_hd__o21ai_1_452/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_193 vssd1 vccd1 sky130_fd_sc_hd__buf_12_19/A sky130_fd_sc_hd__clkbuf_1_53/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_401 sky130_fd_sc_hd__fa_2_398/CIN sky130_fd_sc_hd__fa_2_400/B
+ sky130_fd_sc_hd__fa_2_401/A sky130_fd_sc_hd__fa_2_401/B sky130_fd_sc_hd__xor2_1_599/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_264 vccd1 vssd1 sky130_fd_sc_hd__and3_4_17/X sky130_fd_sc_hd__and2_0_38/A
+ sky130_fd_sc_hd__and2_0_49/A sky130_fd_sc_hd__nor2_2_20/Y sky130_fd_sc_hd__and2_0_45/A
+ sky130_fd_sc_hd__o21ai_1_466/B1 sky130_fd_sc_hd__nor2b_2_4/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_412 sky130_fd_sc_hd__fa_2_411/CIN sky130_fd_sc_hd__or2_0_69/B
+ sky130_fd_sc_hd__fa_2_412/A sky130_fd_sc_hd__fa_2_412/B sky130_fd_sc_hd__xor2_1_625/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_275 vccd1 vssd1 sky130_fd_sc_hd__and3_4_14/X sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__buf_8_0/X sky130_fd_sc_hd__nor2_1_127/Y sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__o21ai_1_480/B1 sky130_fd_sc_hd__nor2b_1_10/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_423 sky130_fd_sc_hd__fah_1_17/A sky130_fd_sc_hd__fa_2_420/A
+ sky130_fd_sc_hd__fa_2_423/A sky130_fd_sc_hd__fa_2_423/B sky130_fd_sc_hd__fa_2_450/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_286 vccd1 vssd1 sky130_fd_sc_hd__and3_4_16/X sky130_fd_sc_hd__buf_2_23/X
+ sky130_fd_sc_hd__buf_2_31/X sky130_fd_sc_hd__nor2_2_19/Y sky130_fd_sc_hd__buf_2_19/X
+ sky130_fd_sc_hd__o21ai_1_494/B1 sky130_fd_sc_hd__nor2b_2_3/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_434 sky130_fd_sc_hd__nor2_1_246/A sky130_fd_sc_hd__nor2_1_247/B
+ sky130_fd_sc_hd__fa_2_434/A sky130_fd_sc_hd__fa_2_434/B sky130_fd_sc_hd__fa_2_434/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_297 vccd1 vssd1 sky130_fd_sc_hd__and3_4_15/X sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__buf_8_0/X sky130_fd_sc_hd__nor2_1_130/Y sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__o21ai_1_508/B1 sky130_fd_sc_hd__nor2b_1_11/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_445 sky130_fd_sc_hd__fa_2_439/B sky130_fd_sc_hd__fa_2_446/CIN
+ sky130_fd_sc_hd__fa_2_445/A sky130_fd_sc_hd__fa_2_445/B sky130_fd_sc_hd__o22ai_1_96/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_456 sky130_fd_sc_hd__fa_2_456/COUT sky130_fd_sc_hd__fa_2_453/A
+ sky130_fd_sc_hd__fa_2_456/A sky130_fd_sc_hd__fa_2_456/B sky130_fd_sc_hd__fa_2_456/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_467 sky130_fd_sc_hd__fa_2_464/B sky130_fd_sc_hd__fa_2_466/A
+ sky130_fd_sc_hd__fa_2_467/A sky130_fd_sc_hd__fa_2_467/B sky130_fd_sc_hd__nor2b_1_33/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_478 sky130_fd_sc_hd__nor2_1_258/B sky130_fd_sc_hd__or2_0_104/A
+ sky130_fd_sc_hd__fa_2_478/A sky130_fd_sc_hd__fa_2_478/B sky130_fd_sc_hd__nor2b_1_55/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_489 sky130_fd_sc_hd__or2_0_109/B sky130_fd_sc_hd__nor2_1_264/A
+ sky130_fd_sc_hd__fa_2_489/A sky130_fd_sc_hd__fa_2_489/B sky130_fd_sc_hd__nor2b_1_77/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_180 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_77/D sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__o21ai_1_97/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_191 vccd1 vssd1 sky130_fd_sc_hd__and2_0_191/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_191/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_12_406 sky130_fd_sc_hd__buf_12_406/A sky130_fd_sc_hd__buf_12_545/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_417 sky130_fd_sc_hd__buf_12_417/A sky130_fd_sc_hd__buf_12_627/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_428 sky130_fd_sc_hd__buf_12_428/A sky130_fd_sc_hd__buf_12_615/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_439 sky130_fd_sc_hd__buf_12_439/A sky130_fd_sc_hd__buf_12_613/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_606 sky130_fd_sc_hd__clkinv_1_606/Y sky130_fd_sc_hd__nand2_1_647/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_617 sky130_fd_sc_hd__o21ai_1_861/A2 sky130_fd_sc_hd__buf_2_28/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_628 sky130_fd_sc_hd__nand2_1_668/A sky130_fd_sc_hd__nor2_1_222/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_639 sky130_fd_sc_hd__clkinv_1_639/Y sky130_fd_sc_hd__nand2_1_691/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__or2_1_10 sky130_fd_sc_hd__or2_1_10/A sky130_fd_sc_hd__or2_1_10/X
+ sky130_fd_sc_hd__or2_1_10/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_1
Xsky130_fd_sc_hd__o21ai_1_170 vssd1 vccd1 sky130_fd_sc_hd__nand2_4_4/Y sky130_fd_sc_hd__nand2b_1_2/Y
+ sky130_fd_sc_hd__a22oi_1_191/Y sky130_fd_sc_hd__xor3_1_5/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_181 vssd1 vccd1 sky130_fd_sc_hd__buf_2_1/X sky130_fd_sc_hd__nand2b_1_4/Y
+ sky130_fd_sc_hd__a222oi_1_60/Y sky130_fd_sc_hd__xor2_1_12/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_192 vssd1 vccd1 sky130_fd_sc_hd__inv_2_20/Y sky130_fd_sc_hd__nand2b_1_6/Y
+ sky130_fd_sc_hd__a222oi_1_68/Y sky130_fd_sc_hd__xor2_1_20/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_15 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_356/Q sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__o211ai_1_31/Y sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__buf_2_203/A sky130_fd_sc_hd__dfxtp_1_307/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_602 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_26 vccd1 vssd1 sky130_fd_sc_hd__xnor2_1_187/Y sky130_fd_sc_hd__inv_2_5/A
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__xnor2_1_62/Y sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__a222oi_1_26/Y sky130_fd_sc_hd__xnor2_1_125/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_37 vccd1 vssd1 sky130_fd_sc_hd__nand2_1_123/A sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__xnor2_1_169/Y sky130_fd_sc_hd__xnor2_1_44/Y sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_37/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_613 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_624 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_48 vccd1 vssd1 sky130_fd_sc_hd__xnor2_2_1/Y sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__buf_2_22/X sky130_fd_sc_hd__o2bb2ai_1_0/Y sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_48/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_635 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_59 vccd1 vssd1 sky130_fd_sc_hd__and3_4_7/X sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__nor2_2_10/B sky130_fd_sc_hd__nor2_2_7/Y sky130_fd_sc_hd__buf_6_4/X
+ sky130_fd_sc_hd__a222oi_1_59/Y sky130_fd_sc_hd__nor2b_2_1/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_646 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_530 sky130_fd_sc_hd__nor2_1_172/A sky130_fd_sc_hd__nand2_1_542/A
+ sky130_fd_sc_hd__or2_0_61/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_17 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_17/B sky130_fd_sc_hd__xnor2_1_17/Y
+ sky130_fd_sc_hd__xnor2_1_17/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_657 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_541 sky130_fd_sc_hd__nor2_1_175/B sky130_fd_sc_hd__or2_0_60/X
+ sky130_fd_sc_hd__or2_0_59/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_668 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_28 vssd1 vccd1 sky130_fd_sc_hd__o21ai_2_8/Y sky130_fd_sc_hd__xnor2_1_28/Y
+ sky130_fd_sc_hd__xnor2_1_28/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_552 sky130_fd_sc_hd__nor2_1_180/A sky130_fd_sc_hd__or2_0_66/X
+ sky130_fd_sc_hd__or2_0_65/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_39 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_39/B sky130_fd_sc_hd__inv_2_21/A
+ sky130_fd_sc_hd__xnor2_1_39/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_679 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_563 sky130_fd_sc_hd__xnor2_1_152/A sky130_fd_sc_hd__nand2_1_564/Y
+ sky130_fd_sc_hd__or2_0_65/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_574 sky130_fd_sc_hd__nand2_1_574/Y sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__buf_4_2/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_585 sky130_fd_sc_hd__o21ai_2_16/A1 sky130_fd_sc_hd__or2_1_1/X
+ sky130_fd_sc_hd__nor2_2_28/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_596 sky130_fd_sc_hd__nand2_1_596/Y sky130_fd_sc_hd__buf_6_4/X
+ sky130_fd_sc_hd__nor2_2_10/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_1110 sky130_fd_sc_hd__clkinv_4_53/A sky130_fd_sc_hd__a22o_1_30/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1121 sky130_fd_sc_hd__clkinv_4_64/A sky130_fd_sc_hd__a22o_1_41/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1132 sky130_fd_sc_hd__clkinv_4_75/A sky130_fd_sc_hd__a22o_1_52/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1143 sky130_fd_sc_hd__clkbuf_4_7/A sky130_fd_sc_hd__clkinv_4_86/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1601 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1612 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_2_6 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_6/Y sky130_fd_sc_hd__mux2_4_4/X
+ la_data_out[77] vssd1 vccd1 sky130_fd_sc_hd__xnor2_2
Xsky130_fd_sc_hd__decap_12_1623 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1634 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1645 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1656 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1667 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_370 sky130_fd_sc_hd__dfxtp_1_370/Q sky130_fd_sc_hd__dfxtp_1_371/CLK
+ sky130_fd_sc_hd__nor2b_1_113/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1678 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_381 sky130_fd_sc_hd__dfxtp_1_381/Q sky130_fd_sc_hd__dfxtp_1_392/CLK
+ sky130_fd_sc_hd__nor2b_1_102/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1689 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_1 sky130_fd_sc_hd__buf_8_0/A sky130_fd_sc_hd__nand2_1_1/B
+ sky130_fd_sc_hd__nand2_1_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_392 sky130_fd_sc_hd__dfxtp_1_392/Q sky130_fd_sc_hd__dfxtp_1_392/CLK
+ sky130_fd_sc_hd__nor2b_1_91/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__or4_1_3 sky130_fd_sc_hd__or4_1_3/C sky130_fd_sc_hd__or4_1_3/A sky130_fd_sc_hd__or4_1_3/X
+ sky130_fd_sc_hd__or4_1_3/B sky130_fd_sc_hd__or4_1_3/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__or4_1
Xsky130_fd_sc_hd__fa_2_220 sky130_fd_sc_hd__fa_2_213/A sky130_fd_sc_hd__fa_2_218/B
+ sky130_fd_sc_hd__fa_2_220/A sky130_fd_sc_hd__fa_2_220/B sky130_fd_sc_hd__fa_2_220/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_231 sky130_fd_sc_hd__fa_2_228/B sky130_fd_sc_hd__fa_2_234/CIN
+ sky130_fd_sc_hd__fa_2_231/A sky130_fd_sc_hd__fa_2_231/B sky130_fd_sc_hd__fa_2_231/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_242 sky130_fd_sc_hd__fa_2_238/A sky130_fd_sc_hd__fa_2_243/B
+ sky130_fd_sc_hd__fa_2_242/A sky130_fd_sc_hd__fa_2_242/B sky130_fd_sc_hd__xor2_1_350/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_253 sky130_fd_sc_hd__fa_2_252/CIN sky130_fd_sc_hd__fah_1_5/B
+ sky130_fd_sc_hd__fa_2_253/A sky130_fd_sc_hd__fa_2_253/B sky130_fd_sc_hd__xor2_1_371/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_264 sky130_fd_sc_hd__fa_2_263/B sky130_fd_sc_hd__fa_2_266/CIN
+ sky130_fd_sc_hd__fa_2_264/A sky130_fd_sc_hd__fa_2_264/B sky130_fd_sc_hd__xor2_1_385/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_275 sky130_fd_sc_hd__fa_2_273/B sky130_fd_sc_hd__fa_2_276/A
+ sky130_fd_sc_hd__fa_2_275/A sky130_fd_sc_hd__fa_2_275/B sky130_fd_sc_hd__fa_2_275/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_286 sky130_fd_sc_hd__xor3_1_21/A sky130_fd_sc_hd__fa_2_287/B
+ sky130_fd_sc_hd__fa_2_286/A sky130_fd_sc_hd__fa_2_286/B sky130_fd_sc_hd__fa_2_286/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_2 vccd1 vssd1 sky130_fd_sc_hd__and2_0_2/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_2/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__fa_2_297 sky130_fd_sc_hd__fa_2_282/B sky130_fd_sc_hd__fa_2_299/CIN
+ sky130_fd_sc_hd__fa_2_297/A sky130_fd_sc_hd__fa_2_297/B sky130_fd_sc_hd__fa_2_298/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22oi_1_8 sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__a22oi_1_8/B2 sky130_fd_sc_hd__a22oi_1_8/A2 sky130_fd_sc_hd__a22oi_1_8/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_203 sky130_fd_sc_hd__buf_6_66/X sky130_fd_sc_hd__buf_12_331/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_50 sky130_fd_sc_hd__o21ai_1_335/Y sky130_fd_sc_hd__a21oi_1_50/B1
+ sky130_fd_sc_hd__o21ai_2_7/B1 sky130_fd_sc_hd__nand2_1_248/A vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_214 sky130_fd_sc_hd__buf_6_40/X sky130_fd_sc_hd__buf_12_394/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_61 sky130_fd_sc_hd__or2_0_16/X sky130_fd_sc_hd__a21oi_1_61/B1
+ sky130_fd_sc_hd__xor2_1_191/B sky130_fd_sc_hd__xnor2_1_54/A vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_225 sky130_fd_sc_hd__buf_6_33/X sky130_fd_sc_hd__buf_12_454/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_72 sky130_fd_sc_hd__o21ai_1_456/Y sky130_fd_sc_hd__o21ai_1_414/Y
+ sky130_fd_sc_hd__o21a_1_2/B1 sky130_fd_sc_hd__nor2_1_107/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_236 sky130_fd_sc_hd__buf_6_84/X sky130_fd_sc_hd__buf_12_442/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_83 sky130_fd_sc_hd__nand2_1_400/Y sky130_fd_sc_hd__nor2_1_125/A
+ sky130_fd_sc_hd__a21oi_1_83/Y sky130_fd_sc_hd__or2_0_44/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_247 sky130_fd_sc_hd__buf_6_54/X sky130_fd_sc_hd__buf_12_335/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_94 sky130_fd_sc_hd__nor2_1_151/Y sky130_fd_sc_hd__o21ai_1_601/Y
+ sky130_fd_sc_hd__xor2_1_389/A sky130_fd_sc_hd__o21ai_1_607/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_1_106 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_180/Q sky130_fd_sc_hd__dfxtp_1_148/Q sky130_fd_sc_hd__o21ai_1_12/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_258 sky130_fd_sc_hd__buf_6_68/X sky130_fd_sc_hd__buf_12_258/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_117 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_169/Q sky130_fd_sc_hd__dfxtp_1_137/Q sky130_fd_sc_hd__o21ai_1_23/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_269 sky130_fd_sc_hd__buf_12_269/A sky130_fd_sc_hd__buf_12_660/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_128 sky130_fd_sc_hd__xor2_2_1/X sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xor2_2_0/X sky130_fd_sc_hd__o21ai_1_36/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_139 sky130_fd_sc_hd__xnor2_1_78/Y sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2_6/Y sky130_fd_sc_hd__xnor2_1_15/Y sky130_fd_sc_hd__o21ai_1_57/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_403 sky130_fd_sc_hd__nand2_1_313/A sky130_fd_sc_hd__nor2_1_103/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_414 sky130_fd_sc_hd__a21oi_1_69/B1 sky130_fd_sc_hd__nand2_1_339/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_425 sky130_fd_sc_hd__a21oi_2_7/B1 sky130_fd_sc_hd__nand2_1_351/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_436 sky130_fd_sc_hd__nand2_1_366/A sky130_fd_sc_hd__nor2_2_13/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_447 sky130_fd_sc_hd__nand2_1_377/A sky130_fd_sc_hd__nor2_2_12/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_458 sky130_fd_sc_hd__nor2_1_125/A sky130_fd_sc_hd__nand2_1_402/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_469 sky130_fd_sc_hd__nand2_1_417/A sky130_fd_sc_hd__nor2_1_135/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_90 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_90 vccd1 vssd1 sky130_fd_sc_hd__buf_6_90/X sky130_fd_sc_hd__buf_6_90/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_70 la_data_out[63] vssd1 vccd1 vccd1 vssd1 sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a222oi_1_3 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_344/Q sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__o211ai_1_19/Y sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__a222oi_1_3/Y sky130_fd_sc_hd__dfxtp_1_295/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_410 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_421 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_432 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_443 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_454 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_465 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_476 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_360 sky130_fd_sc_hd__nand2_1_360/Y sky130_fd_sc_hd__or2_0_39/B
+ sky130_fd_sc_hd__or2_0_42/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_487 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_371 sky130_fd_sc_hd__nand2_1_371/Y sky130_fd_sc_hd__or2_0_60/A
+ sky130_fd_sc_hd__or2_0_61/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_498 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_970 sky130_fd_sc_hd__clkinv_1_970/Y sky130_fd_sc_hd__inv_2_153/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_382 sky130_fd_sc_hd__nand2_1_382/Y sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__or2_0_60/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_981 sky130_fd_sc_hd__clkinv_1_981/Y sky130_fd_sc_hd__clkinv_2_33/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_393 sky130_fd_sc_hd__xnor2_1_91/A sky130_fd_sc_hd__nand2_1_394/Y
+ sky130_fd_sc_hd__or2_0_34/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_992 sky130_fd_sc_hd__clkinv_1_992/Y sky130_fd_sc_hd__inv_2_157/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1420 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1431 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1442 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1453 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1464 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1475 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_906 vssd1 vccd1 sky130_fd_sc_hd__nand2_1_848/A sky130_fd_sc_hd__o21ai_1_908/Y
+ sky130_fd_sc_hd__nand2_1_848/Y sky130_fd_sc_hd__and2_0_400/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1486 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_917 vssd1 vccd1 sky130_fd_sc_hd__nand2_1_859/B la_data_out[43]
+ sky130_fd_sc_hd__a21oi_1_191/Y sky130_fd_sc_hd__nor3_1_3/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1497 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_15 vccd1 vssd1 sky130_fd_sc_hd__buf_2_15/X sky130_fd_sc_hd__buf_2_31/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_26 vccd1 vssd1 sky130_fd_sc_hd__buf_2_26/X sky130_fd_sc_hd__buf_4_7/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_37 vccd1 vssd1 sky130_fd_sc_hd__buf_2_37/X sky130_fd_sc_hd__buf_2_37/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_48 vccd1 vssd1 sky130_fd_sc_hd__buf_2_48/X sky130_fd_sc_hd__buf_2_48/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_59 vccd1 vssd1 sky130_fd_sc_hd__buf_8_84/A sky130_fd_sc_hd__buf_8_6/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o211ai_1_20 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_43/B1
+ sky130_fd_sc_hd__o211ai_1_20/Y sky130_fd_sc_hd__a22oi_1_72/Y sky130_fd_sc_hd__a22oi_1_73/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_31 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_39/B1
+ sky130_fd_sc_hd__o211ai_1_31/Y sky130_fd_sc_hd__a22oi_1_94/Y sky130_fd_sc_hd__a22oi_1_95/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_42 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o22ai_1_21/B1
+ sky130_fd_sc_hd__fa_2_357/B sky130_fd_sc_hd__nand2_1_62/Y sky130_fd_sc_hd__a21oi_1_13/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_53 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o22ai_1_10/B1
+ sky130_fd_sc_hd__fah_1_12/A sky130_fd_sc_hd__nand2_1_73/Y sky130_fd_sc_hd__a21oi_1_24/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_64 sky130_fd_sc_hd__xor2_1_694/X sky130_fd_sc_hd__nand2_1_859/Y
+ sky130_fd_sc_hd__o211ai_1_64/Y sky130_fd_sc_hd__o21ai_1_916/Y sky130_fd_sc_hd__nand2b_1_33/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__clkinv_1_200 sky130_fd_sc_hd__nor2_1_19/A sky130_fd_sc_hd__dfxtp_1_142/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_211 sky130_fd_sc_hd__o22ai_1_52/B1 sky130_fd_sc_hd__dfxtp_1_170/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_222 sky130_fd_sc_hd__o22ai_1_8/B1 sky130_fd_sc_hd__dfxtp_1_103/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_233 sky130_fd_sc_hd__nor2_1_8/A sky130_fd_sc_hd__dfxtp_1_131/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_244 sky130_fd_sc_hd__o22ai_1_2/A2 sky130_fd_sc_hd__dfxtp_1_161/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_255 sky130_fd_sc_hd__o21ai_1_109/A2 sky130_fd_sc_hd__xnor2_1_166/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_266 sky130_fd_sc_hd__o21ai_1_153/A2 sky130_fd_sc_hd__xor2_1_632/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_277 sky130_fd_sc_hd__and2_0_126/A sky130_fd_sc_hd__a222oi_1_21/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_288 sky130_fd_sc_hd__and2_0_191/A sky130_fd_sc_hd__a222oi_1_32/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_299 sky130_fd_sc_hd__and2_0_226/A sky130_fd_sc_hd__a222oi_1_43/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_2_0 sky130_fd_sc_hd__o21ai_2_0/B1 sky130_fd_sc_hd__o21ai_2_0/Y
+ sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__o21ai_2_1/A2 vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__o21ai_2
Xsky130_fd_sc_hd__xor3_1_6 sky130_fd_sc_hd__xor3_1_6/X sky130_fd_sc_hd__xor3_1_7/X
+ sky130_fd_sc_hd__xor3_1_6/B sky130_fd_sc_hd__xor3_1_9/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__a21oi_1_7 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_36/Y
+ sky130_fd_sc_hd__a21oi_1_7/Y sky130_fd_sc_hd__dfxtp_1_89/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__and3_4_13 sky130_fd_sc_hd__and3_4_13/A sky130_fd_sc_hd__nor2b_1_9/A
+ sky130_fd_sc_hd__and3_4_13/C sky130_fd_sc_hd__and3_4_13/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__and3_4_24 sky130_fd_sc_hd__and3_4_24/A sky130_fd_sc_hd__and3_4_24/B
+ sky130_fd_sc_hd__and3_4_24/C sky130_fd_sc_hd__and3_4_24/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__a21oi_1_130 sky130_fd_sc_hd__nor2_1_208/Y sky130_fd_sc_hd__nand2_1_625/Y
+ sky130_fd_sc_hd__o21ai_2_17/B1 sky130_fd_sc_hd__nand2_1_635/Y vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_141 sky130_fd_sc_hd__xnor2_1_191/B sky130_fd_sc_hd__clkinv_1_631/Y
+ sky130_fd_sc_hd__xor2_1_642/A sky130_fd_sc_hd__or2_0_76/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_152 sky130_fd_sc_hd__xnor2_1_206/B sky130_fd_sc_hd__clkinv_1_663/Y
+ sky130_fd_sc_hd__xor2_1_653/A sky130_fd_sc_hd__or2_0_86/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_163 sky130_fd_sc_hd__o21ai_1_885/Y sky130_fd_sc_hd__clkinv_1_693/Y
+ sky130_fd_sc_hd__a21oi_1_163/Y sky130_fd_sc_hd__or2_1_12/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_174 sky130_fd_sc_hd__xnor2_1_295/B sky130_fd_sc_hd__clkinv_1_816/Y
+ sky130_fd_sc_hd__xor2_1_680/A sky130_fd_sc_hd__or2_0_104/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_185 la_data_out[36] sky130_fd_sc_hd__nor2_1_277/B sky130_fd_sc_hd__o31ai_1_0/B1
+ sky130_fd_sc_hd__o31ai_1_1/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_196 sky130_fd_sc_hd__maj3_1_3/X sky130_fd_sc_hd__nor4b_1_0/B
+ sky130_fd_sc_hd__a21oi_1_196/Y sky130_fd_sc_hd__ha_2_55/SUM vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_104 sky130_fd_sc_hd__inv_2_165/Y sky130_fd_sc_hd__buf_8_104/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_115 sky130_fd_sc_hd__buf_8_115/A sky130_fd_sc_hd__buf_6_79/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_126 sky130_fd_sc_hd__buf_2_60/A sky130_fd_sc_hd__buf_6_73/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_137 sky130_fd_sc_hd__inv_2_183/Y sky130_fd_sc_hd__buf_8_137/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_148 sky130_fd_sc_hd__buf_8_148/A sky130_fd_sc_hd__buf_8_148/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_159 sky130_fd_sc_hd__buf_8_159/A sky130_fd_sc_hd__buf_8_159/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__decap_12_240 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_251 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_262 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_273 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_284 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_295 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_190 sky130_fd_sc_hd__xnor2_1_15/A sky130_fd_sc_hd__nand2_1_191/Y
+ sky130_fd_sc_hd__or2_0_2/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_1250 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1261 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1272 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_703 vssd1 vccd1 sky130_fd_sc_hd__xor2_2_2/X sky130_fd_sc_hd__nand2b_1_16/Y
+ sky130_fd_sc_hd__o21ai_1_703/B1 sky130_fd_sc_hd__xor2_1_482/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1283 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_714 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_10/X sky130_fd_sc_hd__nand2_1_540/Y
+ sky130_fd_sc_hd__a21oi_1_114/Y sky130_fd_sc_hd__xnor2_1_143/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1294 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_725 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_780/A2 sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__o21ai_1_725/B1 sky130_fd_sc_hd__xor2_1_501/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_736 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_126/Y sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__o21ai_1_736/B1 sky130_fd_sc_hd__xor2_1_512/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_747 vssd1 vccd1 sky130_fd_sc_hd__inv_2_47/Y sky130_fd_sc_hd__nand2b_2_6/Y
+ sky130_fd_sc_hd__o21ai_1_747/B1 sky130_fd_sc_hd__xor2_1_522/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_758 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_9/X sky130_fd_sc_hd__nand2b_1_15/Y
+ sky130_fd_sc_hd__o21ai_1_758/B1 sky130_fd_sc_hd__xor2_1_533/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_769 vssd1 vccd1 sky130_fd_sc_hd__inv_2_50/Y sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_769/B1 sky130_fd_sc_hd__xor2_1_544/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_10 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__xor3_1_9/A
+ sky130_fd_sc_hd__xor2_1_10/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_21 sky130_fd_sc_hd__xor2_1_21/B sky130_fd_sc_hd__xor2_1_21/X
+ sky130_fd_sc_hd__xor2_1_21/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_32 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__xor2_1_32/X
+ sky130_fd_sc_hd__xor2_1_32/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_43 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__xor2_1_43/X
+ sky130_fd_sc_hd__xor2_1_43/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_54 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__xor2_1_54/X
+ sky130_fd_sc_hd__xor2_1_54/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_65 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__fa_2_46/A
+ sky130_fd_sc_hd__xor2_1_65/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_76 sky130_fd_sc_hd__fa_2_75/A sky130_fd_sc_hd__fa_2_58/B
+ sky130_fd_sc_hd__xor2_1_76/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_87 sky130_fd_sc_hd__xor2_1_6/B sky130_fd_sc_hd__fa_2_65/B
+ sky130_fd_sc_hd__xor2_1_87/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_98 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__fa_2_71/B
+ sky130_fd_sc_hd__xor2_1_98/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2b_1_4 sky130_fd_sc_hd__nand2b_1_4/Y sky130_fd_sc_hd__and3_4_4/C
+ sky130_fd_sc_hd__and3_4_4/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a21o_2_0 sky130_fd_sc_hd__a21o_2_0/X sky130_fd_sc_hd__a21o_2_0/B1
+ sky130_fd_sc_hd__nor3_1_3/Y sky130_fd_sc_hd__a21o_2_0/A2 vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__xor2_1_530 sky130_fd_sc_hd__fa_2_357/A sky130_fd_sc_hd__and3_4_24/A
+ sky130_fd_sc_hd__xor2_1_530/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_541 sky130_fd_sc_hd__xor2_1_548/B sky130_fd_sc_hd__fa_2_367/A
+ sky130_fd_sc_hd__xor2_1_541/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_552 sky130_fd_sc_hd__fah_1_14/A sky130_fd_sc_hd__fa_2_377/B
+ sky130_fd_sc_hd__xor2_1_552/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_563 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__fah_1_11/CI
+ sky130_fd_sc_hd__xor2_1_563/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_574 sky130_fd_sc_hd__fa_2_389/A sky130_fd_sc_hd__xor2_1_574/X
+ sky130_fd_sc_hd__xor2_1_574/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_585 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__fa_2_392/A
+ sky130_fd_sc_hd__xor2_1_585/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_596 sky130_fd_sc_hd__fah_1_14/A sky130_fd_sc_hd__nor2_2_32/B
+ sky130_fd_sc_hd__xor2_1_596/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a221oi_1_2 sky130_fd_sc_hd__nand4_1_1/A sky130_fd_sc_hd__o22ai_1_138/Y
+ sky130_fd_sc_hd__nand4_1_0/B sky130_fd_sc_hd__dfxtp_1_358/Q sky130_fd_sc_hd__ha_2_9/B
+ sky130_fd_sc_hd__nor2_4_19/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__a221oi_1
Xsky130_fd_sc_hd__a222oi_1_605 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_395/Q sky130_fd_sc_hd__and2b_4_13/X
+ sky130_fd_sc_hd__nor2_4_19/Y sky130_fd_sc_hd__nor2_4_19/B sky130_fd_sc_hd__dfxtp_1_459/Q
+ sky130_fd_sc_hd__clkinv_1_802/A sky130_fd_sc_hd__dfxtp_1_427/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_0 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_6/B sky130_fd_sc_hd__fa_2_110/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkinv_1_0 la_data_out[127] sky130_fd_sc_hd__clkinv_1_0/A vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_190 sky130_fd_sc_hd__nor2_1_190/B sky130_fd_sc_hd__nor2_1_190/Y
+ sky130_fd_sc_hd__nor2_1_193/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__and2_0_15 vccd1 vssd1 sky130_fd_sc_hd__and2_0_15/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__buf_2_27/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_26 vccd1 vssd1 sky130_fd_sc_hd__and2_0_26/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__nor2_2_5/B vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_37 vccd1 vssd1 sky130_fd_sc_hd__and2_0_37/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__nor2_1_87/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_48 vccd1 vssd1 sky130_fd_sc_hd__and2_0_48/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__buf_6_1/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_59 vccd1 vssd1 sky130_fd_sc_hd__and2_0_59/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__or2_0_4/B vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nor2_2_7 sky130_fd_sc_hd__nor2_2_7/B sky130_fd_sc_hd__nor2_2_7/Y
+ sky130_fd_sc_hd__nor2_2_7/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__buf_8_14 sky130_fd_sc_hd__buf_8_14/A sky130_fd_sc_hd__buf_8_14/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_25 sky130_fd_sc_hd__buf_8_25/A sky130_fd_sc_hd__buf_8_25/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_36 sky130_fd_sc_hd__buf_8_36/A sky130_fd_sc_hd__buf_8_36/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_47 sky130_fd_sc_hd__ha_2_34/A sky130_fd_sc_hd__buf_8_47/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xnor2_1_160 vssd1 vccd1 sky130_fd_sc_hd__fa_2_389/A sky130_fd_sc_hd__and3_4_25/C
+ sky130_fd_sc_hd__xnor2_1_160/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__buf_8_58 sky130_fd_sc_hd__buf_8_58/A sky130_fd_sc_hd__buf_8_58/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xnor2_1_171 vssd1 vccd1 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__nor2_2_32/A
+ sky130_fd_sc_hd__xnor2_1_171/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__buf_8_69 sky130_fd_sc_hd__inv_4_10/Y sky130_fd_sc_hd__buf_8_69/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xnor2_1_182 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_182/B sky130_fd_sc_hd__xnor2_1_182/Y
+ sky130_fd_sc_hd__xnor2_1_182/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_193 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_193/B sky130_fd_sc_hd__and2_0_267/A
+ sky130_fd_sc_hd__xnor2_1_193/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__o21ai_1_500 vssd1 vccd1 sky130_fd_sc_hd__inv_2_34/Y sky130_fd_sc_hd__nand2b_1_8/Y
+ sky130_fd_sc_hd__o21ai_1_500/B1 sky130_fd_sc_hd__xor2_1_300/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1080 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_511 vssd1 vccd1 sky130_fd_sc_hd__inv_2_31/Y sky130_fd_sc_hd__nand2b_1_9/Y
+ sky130_fd_sc_hd__o21ai_1_511/B1 sky130_fd_sc_hd__xor2_1_310/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1091 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_522 vssd1 vccd1 sky130_fd_sc_hd__buf_2_9/X sky130_fd_sc_hd__nand2b_1_9/Y
+ sky130_fd_sc_hd__o21ai_1_522/B1 sky130_fd_sc_hd__xor2_1_321/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_533 vssd1 vccd1 sky130_fd_sc_hd__inv_2_33/Y sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_533/B1 sky130_fd_sc_hd__xor2_1_332/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_544 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_0/A sky130_fd_sc_hd__nor2_1_131/Y
+ sky130_fd_sc_hd__nand2_1_410/Y sky130_fd_sc_hd__xnor2_1_96/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_555 vssd1 vccd1 sky130_fd_sc_hd__buf_2_8/X sky130_fd_sc_hd__nand2b_2_3/Y
+ sky130_fd_sc_hd__o21ai_1_555/B1 sky130_fd_sc_hd__xor2_1_353/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_566 vssd1 vccd1 sky130_fd_sc_hd__inv_2_35/Y sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_566/B1 sky130_fd_sc_hd__xor2_1_364/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_577 vssd1 vccd1 sky130_fd_sc_hd__inv_2_31/Y sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_577/B1 sky130_fd_sc_hd__xor2_1_373/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_588 vssd1 vccd1 sky130_fd_sc_hd__buf_2_10/X sky130_fd_sc_hd__nand2b_2_3/Y
+ sky130_fd_sc_hd__o21ai_1_588/B1 sky130_fd_sc_hd__xor2_1_381/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_599 vssd1 vccd1 sky130_fd_sc_hd__inv_2_31/Y sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_599/B1 sky130_fd_sc_hd__xor2_1_393/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_360 sky130_fd_sc_hd__fa_2_262/A sky130_fd_sc_hd__fa_2_252/B
+ sky130_fd_sc_hd__xor2_1_360/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_371 sky130_fd_sc_hd__fa_2_262/A sky130_fd_sc_hd__xor2_1_371/X
+ sky130_fd_sc_hd__xor2_1_371/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_382 sky130_fd_sc_hd__fa_2_262/A sky130_fd_sc_hd__xor2_1_382/X
+ sky130_fd_sc_hd__xor2_1_382/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_393 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__fa_2_269/B
+ sky130_fd_sc_hd__xor2_1_393/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_320 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_320/X sky130_fd_sc_hd__clkinv_1_917/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_331 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1_4/D sky130_fd_sc_hd__ha_2_19/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_402 vccd1 vssd1 sky130_fd_sc_hd__and3_4_21/X sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__or2_0_66/A sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__or2_0_60/B
+ sky130_fd_sc_hd__o21ai_1_668/B1 sky130_fd_sc_hd__and2b_4_12/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_342 vssd1 vccd1 sky130_fd_sc_hd__inv_2_4/A sky130_fd_sc_hd__a222oi_1_14/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_413 vccd1 vssd1 sky130_fd_sc_hd__and3_4_24/X sky130_fd_sc_hd__buf_4_7/X
+ sky130_fd_sc_hd__buf_4_0/X sky130_fd_sc_hd__nor2_1_183/Y sky130_fd_sc_hd__buf_2_23/X
+ sky130_fd_sc_hd__o21ai_1_683/B1 sky130_fd_sc_hd__nor2b_1_16/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_353 vssd1 vccd1 sky130_fd_sc_hd__inv_4_1/A sky130_fd_sc_hd__a222oi_1_3/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_424 vccd1 vssd1 sky130_fd_sc_hd__and3_4_18/X sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__nor2_2_10/B sky130_fd_sc_hd__nor2_2_32/Y sky130_fd_sc_hd__buf_6_4/X
+ sky130_fd_sc_hd__o21ai_1_698/B1 sky130_fd_sc_hd__nor2b_2_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_435 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__or2_0_60/A
+ sky130_fd_sc_hd__or2_0_61/A sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__or2_0_61/B
+ sky130_fd_sc_hd__o21ai_1_709/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_446 vccd1 vssd1 sky130_fd_sc_hd__and3_4_21/X sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__nor2_1_73/B sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__o21ai_1_725/B1 sky130_fd_sc_hd__and2b_4_12/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_457 vccd1 vssd1 sky130_fd_sc_hd__and3_4_18/X sky130_fd_sc_hd__buf_2_4/A
+ sky130_fd_sc_hd__buf_2_20/X sky130_fd_sc_hd__nor2_2_32/Y sky130_fd_sc_hd__buf_2_21/X
+ sky130_fd_sc_hd__o21ai_1_739/B1 sky130_fd_sc_hd__nor2b_2_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_468 vccd1 vssd1 sky130_fd_sc_hd__and3_4_25/X sky130_fd_sc_hd__or2_0_72/A
+ sky130_fd_sc_hd__or2_0_71/B sky130_fd_sc_hd__nor2_1_186/Y sky130_fd_sc_hd__buf_2_29/X
+ sky130_fd_sc_hd__o21ai_1_754/B1 sky130_fd_sc_hd__nor2b_1_17/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_479 vccd1 vssd1 sky130_fd_sc_hd__and3_4_26/X sky130_fd_sc_hd__buf_2_29/X
+ sky130_fd_sc_hd__buf_2_30/X sky130_fd_sc_hd__nor2_2_31/Y sky130_fd_sc_hd__buf_2_26/X
+ sky130_fd_sc_hd__o21ai_1_766/B1 sky130_fd_sc_hd__nor2b_1_12/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__dfxtp_1_90 sky130_fd_sc_hd__dfxtp_1_90/Q sky130_fd_sc_hd__dfxtp_1_94/CLK
+ sky130_fd_sc_hd__dfxtp_1_90/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_340 vccd1 vssd1 sky130_fd_sc_hd__and2_0_393/A sky130_fd_sc_hd__ha_2_40/SUM
+ sky130_fd_sc_hd__and2_0_342/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_351 vccd1 vssd1 sky130_fd_sc_hd__and2_0_351/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__buf_2_51/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_362 vccd1 vssd1 sky130_fd_sc_hd__and2_0_362/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__buf_6_6/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_373 vccd1 vssd1 sky130_fd_sc_hd__and2_0_373/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_55/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_384 vccd1 vssd1 sky130_fd_sc_hd__and2_0_384/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_73/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_395 vccd1 vssd1 sky130_fd_sc_hd__and2_0_395/X sky130_fd_sc_hd__and2_0_401/B
+ sky130_fd_sc_hd__and2_0_395/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__conb_1_4 sky130_fd_sc_hd__conb_1_4/LO sky130_fd_sc_hd__conb_1_4/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__inv_2_140 sky130_fd_sc_hd__inv_2_140/A sky130_fd_sc_hd__buf_12_2/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_151 sky130_fd_sc_hd__inv_2_151/A sky130_fd_sc_hd__inv_2_151/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_162 sky130_fd_sc_hd__inv_2_162/A sky130_fd_sc_hd__buf_12_8/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_173 sky130_fd_sc_hd__inv_2_173/A sky130_fd_sc_hd__inv_2_174/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_184 sky130_fd_sc_hd__inv_2_184/A sky130_fd_sc_hd__inv_2_184/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_195 sky130_fd_sc_hd__inv_2_195/A sky130_fd_sc_hd__inv_2_195/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__o22ai_1_103 sky130_fd_sc_hd__nor2b_1_19/A sky130_fd_sc_hd__o22ai_1_103/B1
+ sky130_fd_sc_hd__ha_2_11/B sky130_fd_sc_hd__nand2b_1_27/Y sky130_fd_sc_hd__o22ai_1_66/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_114 sky130_fd_sc_hd__xnor2_2_5/Y sky130_fd_sc_hd__xnor2_1_266/Y
+ sky130_fd_sc_hd__fa_2_454/B sky130_fd_sc_hd__xnor2_1_276/Y sky130_fd_sc_hd__o22ai_1_95/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_125 sky130_fd_sc_hd__xnor2_1_280/Y sky130_fd_sc_hd__xnor2_1_273/Y
+ sky130_fd_sc_hd__fa_2_457/CIN sky130_fd_sc_hd__nor2b_1_19/A sky130_fd_sc_hd__o22ai_1_66/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_136 sky130_fd_sc_hd__dfxtp_1_360/Q sky130_fd_sc_hd__nand4_1_0/D
+ sky130_fd_sc_hd__o22ai_1_136/Y sky130_fd_sc_hd__a221oi_1_0/A1 sky130_fd_sc_hd__dfxtp_1_359/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_2_14 sky130_fd_sc_hd__nor2_2_14/B sky130_fd_sc_hd__nor2_2_14/Y
+ sky130_fd_sc_hd__nor2_2_14/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__nor2_2_25 sky130_fd_sc_hd__nor2_2_25/B sky130_fd_sc_hd__nor2_2_25/Y
+ sky130_fd_sc_hd__nor2_2_25/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__o211ai_1_4 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_4/A2
+ sky130_fd_sc_hd__o211ai_1_4/Y sky130_fd_sc_hd__a22oi_1_40/Y sky130_fd_sc_hd__a22oi_1_41/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__a31oi_1_1 vssd1 vccd1 sky130_fd_sc_hd__a31oi_1_1/Y sky130_fd_sc_hd__nor2_1_267/B
+ sky130_fd_sc_hd__o31ai_1_1/B1 la_data_out[36] sky130_fd_sc_hd__a31oi_1_1/A3 vssd1
+ vccd1 sky130_fd_sc_hd__a31oi_1
Xsky130_fd_sc_hd__o21ai_1_330 vssd1 vccd1 sky130_fd_sc_hd__inv_2_20/Y sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__o21ai_1_330/B1 sky130_fd_sc_hd__xor2_1_150/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_341 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_86/Y sky130_fd_sc_hd__nand2_1_271/Y
+ sky130_fd_sc_hd__nand2_1_266/Y sky130_fd_sc_hd__o21ai_1_341/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_352 vssd1 vccd1 sky130_fd_sc_hd__inv_2_19/Y sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__o21ai_1_352/B1 sky130_fd_sc_hd__xor2_1_167/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_363 vssd1 vccd1 sky130_fd_sc_hd__nand2_4_4/Y sky130_fd_sc_hd__nand2b_2_0/Y
+ sky130_fd_sc_hd__a22oi_1_198/Y sky130_fd_sc_hd__xor2_1_179/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_374 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_1/A sky130_fd_sc_hd__nor2_2_5/Y
+ sky130_fd_sc_hd__nand2_1_292/Y sky130_fd_sc_hd__xnor2_1_52/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_385 vssd1 vccd1 sky130_fd_sc_hd__inv_2_16/Y sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__o21ai_1_385/B1 sky130_fd_sc_hd__xor2_1_201/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_396 vssd1 vccd1 sky130_fd_sc_hd__a21oi_2_9/Y sky130_fd_sc_hd__nor2_2_13/Y
+ sky130_fd_sc_hd__nand2_1_367/Y sky130_fd_sc_hd__xnor2_1_78/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_806 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_817 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_701 sky130_fd_sc_hd__nand2_1_701/Y la_data_out[72] sky130_fd_sc_hd__mux2_2_49/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_828 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_712 sky130_fd_sc_hd__and2_0_284/B sky130_fd_sc_hd__or2_0_84/A
+ sky130_fd_sc_hd__or2_0_84/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_839 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__mux2_2_10 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_10/A1 sky130_fd_sc_hd__buf_2_74/X
+ sky130_fd_sc_hd__mux2_8_0/S sky130_fd_sc_hd__fa_2_419/A vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_723 sky130_fd_sc_hd__xnor2_1_205/A sky130_fd_sc_hd__nand2_1_724/Y
+ sky130_fd_sc_hd__nand2_1_723/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_21 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_21/A1 sky130_fd_sc_hd__buf_2_79/X
+ sky130_fd_sc_hd__mux2_8_0/S sky130_fd_sc_hd__or2_0_75/B vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_734 sky130_fd_sc_hd__xor2_1_654/B sky130_fd_sc_hd__nand2_1_735/Y
+ sky130_fd_sc_hd__nand2_1_734/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_32 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_32/A1 sky130_fd_sc_hd__buf_4_9/X
+ sky130_fd_sc_hd__mux2_8_1/S sky130_fd_sc_hd__mux2_2_32/X vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_745 sky130_fd_sc_hd__xnor2_1_210/B sky130_fd_sc_hd__nand2_1_746/Y
+ sky130_fd_sc_hd__or2_0_91/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_43 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_43/A1 sky130_fd_sc_hd__buf_2_91/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__mux2_2_43/X vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_756 sky130_fd_sc_hd__xor2_1_660/B sky130_fd_sc_hd__nand2_1_771/Y
+ sky130_fd_sc_hd__or2_1_12/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_54 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_54/A1 sky130_fd_sc_hd__buf_4_11/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__or2_0_84/B vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_767 sky130_fd_sc_hd__xor2_1_666/A sky130_fd_sc_hd__nand2_1_784/Y
+ sky130_fd_sc_hd__nand2_1_767/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_778 sky130_fd_sc_hd__nand2_1_778/Y sky130_fd_sc_hd__or2_0_93/A
+ sky130_fd_sc_hd__or2_0_93/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_789 sky130_fd_sc_hd__inv_2_67/A sky130_fd_sc_hd__o31ai_2_0/A2
+ sky130_fd_sc_hd__nand2_1_789/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__conb_1_140 sky130_fd_sc_hd__conb_1_140/LO sky130_fd_sc_hd__clkinv_1_2/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1805 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1816 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1827 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_530 wbs_dat_o[9] sky130_fd_sc_hd__dfxtp_1_533/CLK sky130_fd_sc_hd__nor2b_1_148/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_190 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__fa_2_134/A
+ sky130_fd_sc_hd__xor2_1_190/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1838 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_541 wbs_dat_o[20] sky130_fd_sc_hd__dfxtp_1_544/CLK sky130_fd_sc_hd__nor2b_1_137/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1849 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_552 wbs_dat_o[31] sky130_fd_sc_hd__dfxtp_1_552/CLK sky130_fd_sc_hd__nor2b_1_126/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a222oi_1_210 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__buf_4_6/X sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__buf_4_1/X
+ sky130_fd_sc_hd__o21ai_1_385/B1 sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_150 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_47/A1 sky130_fd_sc_hd__clkbuf_1_150/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_221 vccd1 vssd1 sky130_fd_sc_hd__and3_4_11/X sky130_fd_sc_hd__or2_0_60/B
+ sky130_fd_sc_hd__or2_0_60/A sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__or2_0_61/A
+ sky130_fd_sc_hd__o21ai_1_410/B1 sky130_fd_sc_hd__and2b_4_8/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_161 vssd1 vccd1 sky130_fd_sc_hd__buf_12_55/A sky130_fd_sc_hd__clkbuf_4_26/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_232 vccd1 vssd1 sky130_fd_sc_hd__and3_1_1/X sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__buf_2_32/X sky130_fd_sc_hd__nor2_1_117/Y sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__o21ai_1_425/B1 sky130_fd_sc_hd__nor2b_1_8/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_172 vssd1 vccd1 sky130_fd_sc_hd__a22o_1_31/B2 sky130_fd_sc_hd__clkbuf_1_309/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_243 vccd1 vssd1 sky130_fd_sc_hd__and3_4_16/X sky130_fd_sc_hd__and2_0_38/A
+ sky130_fd_sc_hd__and2_0_49/A sky130_fd_sc_hd__nor2_2_19/Y sky130_fd_sc_hd__and2_0_45/A
+ sky130_fd_sc_hd__o21ai_1_439/B1 sky130_fd_sc_hd__nor2b_2_3/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_183 vssd1 vccd1 sky130_fd_sc_hd__a22o_1_34/B2 sky130_fd_sc_hd__clkbuf_1_183/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_254 vccd1 vssd1 sky130_fd_sc_hd__and3_4_11/X sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__buf_4_4/X sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__o21ai_1_453/B1 sky130_fd_sc_hd__and2b_4_8/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_194 vssd1 vccd1 sky130_fd_sc_hd__buf_12_11/A sky130_fd_sc_hd__clkbuf_1_60/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_402 sky130_fd_sc_hd__fah_1_10/B sky130_fd_sc_hd__fa_2_403/CIN
+ sky130_fd_sc_hd__fa_2_402/A sky130_fd_sc_hd__fa_2_402/B sky130_fd_sc_hd__xor2_1_603/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_265 vccd1 vssd1 sky130_fd_sc_hd__and3_4_16/X sky130_fd_sc_hd__buf_2_19/X
+ sky130_fd_sc_hd__buf_6_5/X sky130_fd_sc_hd__nor2_2_19/Y sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__o21ai_1_467/B1 sky130_fd_sc_hd__nor2b_2_3/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_413 sky130_fd_sc_hd__fa_2_412/B sky130_fd_sc_hd__or2_0_68/A
+ sky130_fd_sc_hd__fa_2_413/A sky130_fd_sc_hd__fa_2_413/B sky130_fd_sc_hd__fa_2_413/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_276 vccd1 vssd1 sky130_fd_sc_hd__and3_4_17/X sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__and2_0_38/A sky130_fd_sc_hd__nor2_2_20/Y sky130_fd_sc_hd__and2_0_49/A
+ sky130_fd_sc_hd__o21ai_1_482/B1 sky130_fd_sc_hd__nor2b_2_4/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_424 sky130_fd_sc_hd__nor2_1_243/A sky130_fd_sc_hd__nor2_1_244/B
+ sky130_fd_sc_hd__fa_2_424/A sky130_fd_sc_hd__fa_2_424/B sky130_fd_sc_hd__fa_2_424/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_287 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__buf_4_2/X sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__o21ai_1_495/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_435 sky130_fd_sc_hd__fa_2_434/B sky130_fd_sc_hd__fa_2_437/CIN
+ sky130_fd_sc_hd__fa_2_435/A sky130_fd_sc_hd__fa_2_435/B sky130_fd_sc_hd__fa_2_435/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_298 vccd1 vssd1 sky130_fd_sc_hd__and3_4_10/X sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__and2_0_38/A sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__and2_0_49/A
+ sky130_fd_sc_hd__o21ai_1_510/B1 sky130_fd_sc_hd__and2b_4_7/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_446 sky130_fd_sc_hd__nor2_1_251/A sky130_fd_sc_hd__nor2_1_252/B
+ sky130_fd_sc_hd__fa_2_446/A sky130_fd_sc_hd__fa_2_446/B sky130_fd_sc_hd__fa_2_446/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_457 sky130_fd_sc_hd__fa_2_452/CIN sky130_fd_sc_hd__fa_2_459/A
+ sky130_fd_sc_hd__fa_2_457/A sky130_fd_sc_hd__fa_2_457/B sky130_fd_sc_hd__fa_2_457/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_468 sky130_fd_sc_hd__fa_2_466/B sky130_fd_sc_hd__or2_0_99/A
+ sky130_fd_sc_hd__fa_2_468/A sky130_fd_sc_hd__fa_2_468/B sky130_fd_sc_hd__nor2b_1_35/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_479 sky130_fd_sc_hd__or2_0_104/B sky130_fd_sc_hd__nor2_1_259/A
+ sky130_fd_sc_hd__fa_2_479/A sky130_fd_sc_hd__fa_2_479/B sky130_fd_sc_hd__nor2b_1_57/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_170 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_76/D sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_170/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_181 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_45/D sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__o21ai_1_96/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_192 vccd1 vssd1 sky130_fd_sc_hd__and2_0_192/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__o21ai_1_89/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_12_407 sky130_fd_sc_hd__buf_12_407/A sky130_fd_sc_hd__buf_12_630/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_418 sky130_fd_sc_hd__buf_12_418/A sky130_fd_sc_hd__buf_12_622/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_429 sky130_fd_sc_hd__buf_12_429/A sky130_fd_sc_hd__buf_12_621/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_607 sky130_fd_sc_hd__xnor2_1_182/B sky130_fd_sc_hd__a21oi_1_136/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_618 sky130_fd_sc_hd__nand2_1_599/A sky130_fd_sc_hd__nand2_1_604/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_629 sky130_fd_sc_hd__clkinv_1_629/Y sky130_fd_sc_hd__nand2_1_671/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__or2_1_11 sky130_fd_sc_hd__or2_1_11/A sky130_fd_sc_hd__or2_1_11/X
+ sky130_fd_sc_hd__or2_1_11/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_1
Xsky130_fd_sc_hd__o21ai_1_160 vssd1 vccd1 sky130_fd_sc_hd__nand2_2_9/Y sky130_fd_sc_hd__o21ai_1_160/A1
+ sky130_fd_sc_hd__a22oi_1_190/Y sky130_fd_sc_hd__and2_0_102/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_171 vssd1 vccd1 sky130_fd_sc_hd__inv_2_12/Y sky130_fd_sc_hd__nand2b_1_6/Y
+ sky130_fd_sc_hd__a222oi_1_52/Y sky130_fd_sc_hd__xor2_1_4/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_182 vssd1 vccd1 sky130_fd_sc_hd__inv_2_19/Y sky130_fd_sc_hd__nand2b_1_5/Y
+ sky130_fd_sc_hd__a222oi_1_61/Y sky130_fd_sc_hd__xor2_1_13/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_193 vssd1 vccd1 sky130_fd_sc_hd__inv_2_9/Y sky130_fd_sc_hd__nand2b_1_6/Y
+ sky130_fd_sc_hd__a222oi_1_69/Y sky130_fd_sc_hd__xor2_1_22/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_16 vccd1 vssd1 sky130_fd_sc_hd__nand2_1_129/A sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__xnor2_1_175/Y sky130_fd_sc_hd__xnor2_1_50/Y sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_16/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_603 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_27 vccd1 vssd1 sky130_fd_sc_hd__xnor2_1_86/Y sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__inv_2_57/A sky130_fd_sc_hd__xnor2_1_23/Y sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_27/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_38 vccd1 vssd1 sky130_fd_sc_hd__xor2_1_384/X sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__xor2_1_597/X sky130_fd_sc_hd__xor2_1_171/X sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_38/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_614 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_625 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_49 vccd1 vssd1 sky130_fd_sc_hd__and3_4_1/X sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__buf_4_5/X sky130_fd_sc_hd__nor2_2_9/Y sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__a222oi_1_49/Y sky130_fd_sc_hd__and2b_4_3/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_636 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_520 sky130_fd_sc_hd__xnor2_1_135/A sky130_fd_sc_hd__nand2_1_521/Y
+ sky130_fd_sc_hd__or2_0_57/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_647 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_531 sky130_fd_sc_hd__xnor2_1_139/A sky130_fd_sc_hd__nand2_1_532/Y
+ sky130_fd_sc_hd__nand2_1_531/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_658 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_18 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_78/A sky130_fd_sc_hd__and3_4_4/B
+ sky130_fd_sc_hd__xnor2_1_21/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_542 sky130_fd_sc_hd__xnor2_1_143/A sky130_fd_sc_hd__nand2_1_543/Y
+ sky130_fd_sc_hd__nand2_1_542/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_669 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_29 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_29/B sky130_fd_sc_hd__xnor2_1_29/Y
+ sky130_fd_sc_hd__xnor2_1_29/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_553 sky130_fd_sc_hd__xnor2_1_148/A sky130_fd_sc_hd__nand2_1_554/Y
+ sky130_fd_sc_hd__or2_0_59/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_564 sky130_fd_sc_hd__nand2_1_564/Y sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__buf_4_4/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_0 sky130_fd_sc_hd__nor2b_1_0/B_N sky130_fd_sc_hd__nor2b_1_0/Y
+ la_data_out[32] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nand2_1_575 sky130_fd_sc_hd__xnor2_1_158/A sky130_fd_sc_hd__nand2_1_576/Y
+ sky130_fd_sc_hd__or2_1_2/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_586 sky130_fd_sc_hd__xnor2_1_161/A sky130_fd_sc_hd__nand2_1_587/Y
+ sky130_fd_sc_hd__or2_1_3/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_597 sky130_fd_sc_hd__xor2_1_580/B sky130_fd_sc_hd__nand2_1_598/Y
+ sky130_fd_sc_hd__nand2_1_597/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_1100 sky130_fd_sc_hd__nand2_1_865/B wbs_adr_i[8] vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1111 sky130_fd_sc_hd__clkinv_4_54/A sky130_fd_sc_hd__a22o_1_31/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1122 sky130_fd_sc_hd__clkinv_4_65/A sky130_fd_sc_hd__a22o_1_42/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1133 sky130_fd_sc_hd__clkinv_4_76/A sky130_fd_sc_hd__a22o_1_53/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1144 sky130_fd_sc_hd__clkbuf_4_8/A sky130_fd_sc_hd__clkinv_4_87/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1602 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1613 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1624 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1635 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1646 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1657 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_360 sky130_fd_sc_hd__dfxtp_1_360/Q sky130_fd_sc_hd__dfxtp_1_29/CLK
+ sky130_fd_sc_hd__ha_2_6/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1668 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_371 sky130_fd_sc_hd__dfxtp_1_371/Q sky130_fd_sc_hd__dfxtp_1_371/CLK
+ sky130_fd_sc_hd__nor2b_1_112/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1679 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_382 sky130_fd_sc_hd__dfxtp_1_382/Q sky130_fd_sc_hd__dfxtp_1_392/CLK
+ sky130_fd_sc_hd__nor2b_1_101/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_2 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__nand2_1_7/B
+ sky130_fd_sc_hd__mux2_4_2/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_393 sky130_fd_sc_hd__dfxtp_1_393/Q sky130_fd_sc_hd__dfxtp_1_395/CLK
+ sky130_fd_sc_hd__nor2b_1_90/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_210 sky130_fd_sc_hd__fa_2_205/B sky130_fd_sc_hd__fa_2_212/B
+ sky130_fd_sc_hd__fa_2_210/A sky130_fd_sc_hd__fa_2_210/B sky130_fd_sc_hd__xor2_1_305/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_221 sky130_fd_sc_hd__fa_2_209/B sky130_fd_sc_hd__fa_2_221/SUM
+ sky130_fd_sc_hd__fa_2_221/A sky130_fd_sc_hd__fa_2_221/B sky130_fd_sc_hd__xor2_1_319/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_232 sky130_fd_sc_hd__fa_2_224/B sky130_fd_sc_hd__fa_2_233/A
+ sky130_fd_sc_hd__fa_2_232/A sky130_fd_sc_hd__fa_2_232/B sky130_fd_sc_hd__fa_2_232/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_243 sky130_fd_sc_hd__fa_2_240/B sky130_fd_sc_hd__fa_2_245/CIN
+ sky130_fd_sc_hd__fa_2_243/A sky130_fd_sc_hd__fa_2_243/B sky130_fd_sc_hd__fa_2_243/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_254 sky130_fd_sc_hd__fah_1_2/B sky130_fd_sc_hd__fa_2_255/CIN
+ sky130_fd_sc_hd__fa_2_254/A sky130_fd_sc_hd__fa_2_254/B sky130_fd_sc_hd__fa_2_254/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_265 sky130_fd_sc_hd__fa_2_260/CIN sky130_fd_sc_hd__fa_2_264/B
+ sky130_fd_sc_hd__fa_2_265/A sky130_fd_sc_hd__fa_2_265/B sky130_fd_sc_hd__xor2_1_386/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_276 sky130_fd_sc_hd__nor2_1_154/A sky130_fd_sc_hd__nor2_1_155/B
+ sky130_fd_sc_hd__fa_2_276/A sky130_fd_sc_hd__fa_2_276/B sky130_fd_sc_hd__xor2_1_404/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_287 sky130_fd_sc_hd__xor3_1_20/B sky130_fd_sc_hd__fa_2_287/SUM
+ sky130_fd_sc_hd__fa_2_287/A sky130_fd_sc_hd__fa_2_287/B sky130_fd_sc_hd__fa_2_287/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_3 vccd1 vssd1 sky130_fd_sc_hd__and2_0_3/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_3/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__fa_2_298 sky130_fd_sc_hd__fa_2_282/A sky130_fd_sc_hd__fa_2_298/SUM
+ sky130_fd_sc_hd__fa_2_298/A sky130_fd_sc_hd__fa_2_298/B sky130_fd_sc_hd__fa_2_298/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22oi_1_9 sky130_fd_sc_hd__nor2_4_0/Y sky130_fd_sc_hd__nor2_2_0/Y
+ sky130_fd_sc_hd__a22oi_1_9/B2 sky130_fd_sc_hd__nor2_1_237/A sky130_fd_sc_hd__a22oi_1_9/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__fa_2_90 sky130_fd_sc_hd__fa_2_82/B sky130_fd_sc_hd__fa_2_91/A sky130_fd_sc_hd__fa_2_90/A
+ sky130_fd_sc_hd__fa_2_90/B sky130_fd_sc_hd__fa_2_90/CIN vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a21oi_1_40 sky130_fd_sc_hd__a21oi_1_45/A1 sky130_fd_sc_hd__o21ai_1_201/Y
+ sky130_fd_sc_hd__a21oi_1_40/Y sky130_fd_sc_hd__nor2_1_50/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_204 sky130_fd_sc_hd__buf_6_64/X sky130_fd_sc_hd__buf_12_437/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_51 sky130_fd_sc_hd__a21oi_1_54/A1 sky130_fd_sc_hd__o21ai_1_327/Y
+ sky130_fd_sc_hd__a21oi_1_51/Y sky130_fd_sc_hd__nor2_1_76/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_215 sky130_fd_sc_hd__buf_6_35/X sky130_fd_sc_hd__buf_12_457/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_62 sky130_fd_sc_hd__xnor2_1_56/B sky130_fd_sc_hd__nand2_1_293/Y
+ sky130_fd_sc_hd__xnor2_1_1/A sky130_fd_sc_hd__nor2_1_44/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_226 sky130_fd_sc_hd__buf_6_31/X sky130_fd_sc_hd__buf_12_419/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_73 sky130_fd_sc_hd__a21oi_1_80/A1 sky130_fd_sc_hd__o21ai_1_423/Y
+ sky130_fd_sc_hd__a21oi_1_73/Y sky130_fd_sc_hd__nor2_1_108/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_237 sky130_fd_sc_hd__buf_6_81/X sky130_fd_sc_hd__buf_12_279/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_84 sky130_fd_sc_hd__nand2_1_421/Y sky130_fd_sc_hd__nand2_1_411/Y
+ sky130_fd_sc_hd__a21oi_1_84/Y sky130_fd_sc_hd__nor2_1_133/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_248 sky130_fd_sc_hd__buf_6_28/X sky130_fd_sc_hd__buf_12_444/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_95 sky130_fd_sc_hd__nor2_1_153/Y sky130_fd_sc_hd__nand2_1_454/Y
+ sky130_fd_sc_hd__a21oi_1_95/Y sky130_fd_sc_hd__nand2_1_464/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_1_107 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_179/Q sky130_fd_sc_hd__dfxtp_1_147/Q sky130_fd_sc_hd__o21ai_1_13/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_259 sky130_fd_sc_hd__buf_6_70/X sky130_fd_sc_hd__buf_12_259/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_118 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_168/Q sky130_fd_sc_hd__dfxtp_1_136/Q sky130_fd_sc_hd__o21ai_1_24/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_129 sky130_fd_sc_hd__xor2_2_1/X sky130_fd_sc_hd__xor2_2_0/X
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__nor2_1_2/A sky130_fd_sc_hd__o21ai_1_37/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_404 sky130_fd_sc_hd__a21oi_1_68/B1 sky130_fd_sc_hd__nand2_1_321/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_415 sky130_fd_sc_hd__o21ai_1_412/A2 sky130_fd_sc_hd__xnor2_1_69/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_426 sky130_fd_sc_hd__o21ai_1_442/A2 sky130_fd_sc_hd__xnor2_1_74/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_437 sky130_fd_sc_hd__o21ai_1_476/A2 sky130_fd_sc_hd__xnor2_1_80/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_448 sky130_fd_sc_hd__o21ai_1_496/A2 sky130_fd_sc_hd__xnor2_1_85/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_459 sky130_fd_sc_hd__nand2_1_398/A sky130_fd_sc_hd__nor2_2_15/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_80 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_91 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_80 vccd1 vssd1 sky130_fd_sc_hd__buf_6_80/X sky130_fd_sc_hd__buf_8_67/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_91 vccd1 vssd1 sky130_fd_sc_hd__buf_6_91/X la_data_out[38]
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_60 sky130_fd_sc_hd__buf_2_192/A vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_71 la_data_out[36] vssd1 vccd1 vccd1 vssd1 sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a222oi_1_4 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_345/Q sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__o211ai_1_20/Y sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__a222oi_1_4/Y sky130_fd_sc_hd__dfxtp_1_296/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_400 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_411 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_422 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_433 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_444 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_455 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_466 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_350 sky130_fd_sc_hd__xnor2_1_73/A sky130_fd_sc_hd__nand2_1_351/Y
+ sky130_fd_sc_hd__or2_0_28/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_477 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_361 sky130_fd_sc_hd__xnor2_1_78/A sky130_fd_sc_hd__nand2_1_362/Y
+ sky130_fd_sc_hd__or2_0_29/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_488 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_960 sky130_fd_sc_hd__clkinv_1_961/A sky130_fd_sc_hd__buf_4_8/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_372 sky130_fd_sc_hd__xnor2_1_82/A sky130_fd_sc_hd__nand2_1_373/Y
+ sky130_fd_sc_hd__or2_0_30/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_499 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_971 sky130_fd_sc_hd__clkinv_1_971/Y sky130_fd_sc_hd__inv_8_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_383 sky130_fd_sc_hd__xnor2_1_86/A sky130_fd_sc_hd__nand2_1_384/Y
+ sky130_fd_sc_hd__or2_0_33/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_982 sky130_fd_sc_hd__clkinv_1_982/Y sky130_fd_sc_hd__clkinv_4_27/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_394 sky130_fd_sc_hd__nand2_1_394/Y sky130_fd_sc_hd__or2_0_34/A
+ sky130_fd_sc_hd__or2_0_34/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_993 sky130_fd_sc_hd__clkinv_1_994/A sky130_fd_sc_hd__inv_2_3/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1410 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1421 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1432 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1443 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1454 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1465 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1476 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_907 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_278/B sky130_fd_sc_hd__nor2_1_275/Y
+ sky130_fd_sc_hd__a22o_1_71/B1 sky130_fd_sc_hd__o21ai_1_907/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1487 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_190 sky130_fd_sc_hd__dfxtp_1_190/Q sky130_fd_sc_hd__dfxtp_1_190/CLK
+ sky130_fd_sc_hd__and2_0_4/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_918 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_918/A2 la_data_out[45]
+ sky130_fd_sc_hd__xnor2_1_307/Y sky130_fd_sc_hd__o21ai_1_918/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1498 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_16 vccd1 vssd1 sky130_fd_sc_hd__buf_2_16/X sky130_fd_sc_hd__buf_2_16/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_27 vccd1 vssd1 sky130_fd_sc_hd__buf_2_27/X sky130_fd_sc_hd__buf_2_27/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_38 vccd1 vssd1 sky130_fd_sc_hd__buf_2_38/X wbs_dat_i[21] vssd1
+ vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_49 vccd1 vssd1 sky130_fd_sc_hd__buf_2_49/X sky130_fd_sc_hd__buf_2_49/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o211ai_1_10 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_53/B1
+ sky130_fd_sc_hd__o211ai_1_10/Y sky130_fd_sc_hd__a22oi_1_52/Y sky130_fd_sc_hd__a22oi_1_53/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_21 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_42/B1
+ sky130_fd_sc_hd__o211ai_1_21/Y sky130_fd_sc_hd__a22oi_1_74/Y sky130_fd_sc_hd__a22oi_1_75/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_32 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o21ai_1_2/A2
+ sky130_fd_sc_hd__fa_2_294/A sky130_fd_sc_hd__nand2_1_52/Y sky130_fd_sc_hd__a21oi_1_3/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_43 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o22ai_1_20/B1
+ sky130_fd_sc_hd__fa_2_364/A sky130_fd_sc_hd__nand2_1_63/Y sky130_fd_sc_hd__a21oi_1_14/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_54 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o22ai_1_9/B1
+ sky130_fd_sc_hd__fah_1_15/B sky130_fd_sc_hd__nand2_1_74/Y sky130_fd_sc_hd__a21oi_1_25/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_65 sky130_fd_sc_hd__xor2_1_696/X sky130_fd_sc_hd__nand2_1_861/Y
+ sky130_fd_sc_hd__o211ai_1_65/Y sky130_fd_sc_hd__o21ai_1_920/Y sky130_fd_sc_hd__nand2b_1_34/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__clkinv_1_201 sky130_fd_sc_hd__o22ai_1_15/B1 sky130_fd_sc_hd__dfxtp_1_110/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_212 sky130_fd_sc_hd__nor2_1_15/A sky130_fd_sc_hd__dfxtp_1_138/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_223 sky130_fd_sc_hd__o22ai_1_7/A2 sky130_fd_sc_hd__dfxtp_1_166/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_234 sky130_fd_sc_hd__o22ai_1_4/B1 sky130_fd_sc_hd__dfxtp_1_99/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_245 sky130_fd_sc_hd__nor2_1_6/A sky130_fd_sc_hd__dfxtp_1_129/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_256 sky130_fd_sc_hd__o21ai_1_113/A2 sky130_fd_sc_hd__xnor2_1_169/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_267 sky130_fd_sc_hd__o21ai_1_157/A2 sky130_fd_sc_hd__xor2_1_634/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_278 sky130_fd_sc_hd__and2_0_121/A sky130_fd_sc_hd__a222oi_1_22/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_289 sky130_fd_sc_hd__and2_0_186/A sky130_fd_sc_hd__a222oi_1_33/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_2_1 sky130_fd_sc_hd__buf_2_16/A sky130_fd_sc_hd__o21ai_2_1/Y
+ sky130_fd_sc_hd__o21ai_2_1/A2 sky130_fd_sc_hd__a21oi_1_1/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__o21ai_2
Xsky130_fd_sc_hd__xor3_1_7 sky130_fd_sc_hd__xor3_1_7/X sky130_fd_sc_hd__xor3_1_8/X
+ sky130_fd_sc_hd__xor3_1_7/B sky130_fd_sc_hd__xor3_1_7/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__a21oi_1_8 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_37/Y
+ sky130_fd_sc_hd__a21oi_1_8/Y sky130_fd_sc_hd__dfxtp_1_88/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__and3_4_14 sky130_fd_sc_hd__and3_4_14/A sky130_fd_sc_hd__and3_4_14/B
+ sky130_fd_sc_hd__and3_4_14/C sky130_fd_sc_hd__and3_4_14/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__and3_4_25 sky130_fd_sc_hd__and3_4_25/A sky130_fd_sc_hd__and3_4_25/B
+ sky130_fd_sc_hd__and3_4_25/C sky130_fd_sc_hd__and3_4_25/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__a21oi_1_120 sky130_fd_sc_hd__o21ai_1_633/Y sky130_fd_sc_hd__clkinv_1_574/Y
+ sky130_fd_sc_hd__o21ai_2_16/B1 sky130_fd_sc_hd__or2_1_1/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_131 sky130_fd_sc_hd__or2_0_62/X sky130_fd_sc_hd__clkinv_1_599/Y
+ sky130_fd_sc_hd__xor2_1_616/B sky130_fd_sc_hd__xnor2_1_179/A vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_142 sky130_fd_sc_hd__xnor2_1_192/B sky130_fd_sc_hd__clkinv_1_633/Y
+ sky130_fd_sc_hd__xor2_1_643/A sky130_fd_sc_hd__or2_1_11/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_153 sky130_fd_sc_hd__nor2_1_236/Y sky130_fd_sc_hd__o21ai_1_876/Y
+ sky130_fd_sc_hd__a21oi_1_153/Y sky130_fd_sc_hd__o21ai_1_878/Y vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_164 sky130_fd_sc_hd__o21ai_1_887/Y sky130_fd_sc_hd__o21ai_1_886/Y
+ sky130_fd_sc_hd__a21oi_1_164/Y sky130_fd_sc_hd__nor2_1_245/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_175 sky130_fd_sc_hd__xnor2_1_296/B sky130_fd_sc_hd__clkinv_1_818/Y
+ sky130_fd_sc_hd__xor2_1_681/A sky130_fd_sc_hd__or2_0_105/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_186 sky130_fd_sc_hd__nor2_1_278/Y sky130_fd_sc_hd__a21oi_1_187/Y
+ sky130_fd_sc_hd__and2_0_342/A sky130_fd_sc_hd__nand2_1_855/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_197 sky130_fd_sc_hd__ha_2_56/B la_data_out[48] sky130_fd_sc_hd__a21oi_1_197/Y
+ la_data_out[49] vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_105 sky130_fd_sc_hd__buf_8_105/A sky130_fd_sc_hd__buf_8_105/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_116 sky130_fd_sc_hd__buf_8_116/A sky130_fd_sc_hd__buf_8_116/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_127 sky130_fd_sc_hd__buf_8_127/A sky130_fd_sc_hd__buf_8_127/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_138 sky130_fd_sc_hd__buf_8_138/A sky130_fd_sc_hd__buf_8_138/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_149 sky130_fd_sc_hd__buf_8_149/A sky130_fd_sc_hd__buf_8_149/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_12_590 sky130_fd_sc_hd__buf_12_590/A sky130_fd_sc_hd__buf_12_590/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_230 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_241 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_252 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_263 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_274 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_285 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_296 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_180 sky130_fd_sc_hd__nand2_1_180/Y sky130_fd_sc_hd__or2_0_1/A
+ sky130_fd_sc_hd__or2_0_1/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_191 sky130_fd_sc_hd__nand2_1_191/Y sky130_fd_sc_hd__or2_0_2/A
+ sky130_fd_sc_hd__or2_0_2/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_790 sky130_fd_sc_hd__and2_0_317/A sky130_fd_sc_hd__clkinv_1_790/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1240 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1251 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1262 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1273 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_704 vssd1 vccd1 sky130_fd_sc_hd__inv_2_43/Y sky130_fd_sc_hd__nand2b_1_15/Y
+ sky130_fd_sc_hd__o21ai_1_704/B1 sky130_fd_sc_hd__xor2_1_483/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1284 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_715 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_771/A2 sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__o21ai_1_715/B1 sky130_fd_sc_hd__xor2_1_492/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1295 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_726 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_2/Y sky130_fd_sc_hd__nand2b_1_20/Y
+ sky130_fd_sc_hd__o21ai_1_726/B1 sky130_fd_sc_hd__xor2_1_502/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_737 vssd1 vccd1 sky130_fd_sc_hd__inv_2_49/Y sky130_fd_sc_hd__nand2b_1_15/Y
+ sky130_fd_sc_hd__o21ai_1_737/B1 sky130_fd_sc_hd__xor2_1_513/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_748 vssd1 vccd1 sky130_fd_sc_hd__inv_2_44/Y sky130_fd_sc_hd__nand2b_1_16/Y
+ sky130_fd_sc_hd__o21ai_1_748/B1 sky130_fd_sc_hd__xor2_1_523/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_759 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_3/Y sky130_fd_sc_hd__nand2b_1_16/Y
+ sky130_fd_sc_hd__o21ai_1_759/B1 sky130_fd_sc_hd__xor2_1_534/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_11 sky130_fd_sc_hd__xor2_1_6/B sky130_fd_sc_hd__fa_2_7/CIN
+ sky130_fd_sc_hd__xor2_1_11/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_22 sky130_fd_sc_hd__fa_2_97/A sky130_fd_sc_hd__fa_2_9/CIN
+ sky130_fd_sc_hd__xor2_1_22/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_33 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__fa_2_20/B
+ sky130_fd_sc_hd__xor2_1_33/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_44 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__fa_2_27/B
+ sky130_fd_sc_hd__xor2_1_44/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_55 sky130_fd_sc_hd__fa_2_97/A sky130_fd_sc_hd__fa_2_38/B
+ sky130_fd_sc_hd__xor2_1_55/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_66 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__xor2_1_66/X
+ sky130_fd_sc_hd__xor2_1_66/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_77 sky130_fd_sc_hd__fa_2_56/A sky130_fd_sc_hd__xor2_1_77/X
+ sky130_fd_sc_hd__xor2_1_77/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_88 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__fa_2_65/A
+ sky130_fd_sc_hd__xor2_1_88/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_99 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__fa_2_67/A
+ sky130_fd_sc_hd__xor2_1_99/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2b_1_5 sky130_fd_sc_hd__nand2b_1_5/Y sky130_fd_sc_hd__and3_4_5/C
+ sky130_fd_sc_hd__and3_4_5/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a21o_2_1 sky130_fd_sc_hd__a21o_2_1/X sky130_fd_sc_hd__a21o_2_1/B1
+ wbs_adr_i[2] wbs_adr_i[3] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__xor2_1_520 sky130_fd_sc_hd__fa_2_379/A sky130_fd_sc_hd__fa_2_351/B
+ sky130_fd_sc_hd__xor2_1_520/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_531 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__fa_2_358/A
+ sky130_fd_sc_hd__xor2_1_531/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_542 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__fa_2_363/B
+ sky130_fd_sc_hd__xor2_1_542/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_553 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__fa_2_377/A
+ sky130_fd_sc_hd__xor2_1_553/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_564 sky130_fd_sc_hd__fa_2_389/A sky130_fd_sc_hd__xor2_1_564/X
+ sky130_fd_sc_hd__xor2_1_564/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_575 sky130_fd_sc_hd__fa_2_389/A sky130_fd_sc_hd__nor2_2_31/B
+ sky130_fd_sc_hd__xor2_1_575/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_586 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__xor2_1_586/X
+ sky130_fd_sc_hd__xor2_1_586/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_597 sky130_fd_sc_hd__xor2_1_597/B sky130_fd_sc_hd__xor2_1_597/X
+ sky130_fd_sc_hd__xor2_1_597/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a221oi_1_3 sky130_fd_sc_hd__a31oi_1_0/B1 sky130_fd_sc_hd__nor2_1_278/B
+ sky130_fd_sc_hd__nor2_4_0/A sky130_fd_sc_hd__nand2_1_855/Y sky130_fd_sc_hd__a221oi_1_3/B2
+ sky130_fd_sc_hd__nor2_2_0/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__a221oi_1
Xsky130_fd_sc_hd__a222oi_1_606 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_424/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_456/Q sky130_fd_sc_hd__nor2_4_19/B
+ sky130_fd_sc_hd__clkinv_1_803/A sky130_fd_sc_hd__dfxtp_1_392/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__and2b_4_0 sky130_fd_sc_hd__nor2b_1_1/Y sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_4_4/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__and2b_4
Xsky130_fd_sc_hd__ha_2_60 vssd1 vccd1 sky130_fd_sc_hd__ha_2_60/A sky130_fd_sc_hd__ha_2_59/B
+ sky130_fd_sc_hd__ha_2_60/SUM sky130_fd_sc_hd__ha_2_60/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_9/B sky130_fd_sc_hd__fa_2_122/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkinv_1_1 la_data_out[126] sky130_fd_sc_hd__clkinv_1_1/A vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_180 sky130_fd_sc_hd__nor2_1_182/A sky130_fd_sc_hd__nor2_1_180/Y
+ sky130_fd_sc_hd__nor2_1_180/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_191 sky130_fd_sc_hd__buf_6_4/X sky130_fd_sc_hd__nor2_1_191/Y
+ sky130_fd_sc_hd__buf_6_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__and2_0_16 vccd1 vssd1 sky130_fd_sc_hd__and2_0_16/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__buf_4_0/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_27 vccd1 vssd1 sky130_fd_sc_hd__and2_0_27/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__buf_8_0/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_38 vccd1 vssd1 sky130_fd_sc_hd__and2_0_38/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__and2_0_38/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_49 vccd1 vssd1 sky130_fd_sc_hd__and2_0_49/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__and2_0_49/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nor2_2_8 sky130_fd_sc_hd__nor2_2_8/B sky130_fd_sc_hd__nor2_2_8/Y
+ sky130_fd_sc_hd__nor2_2_8/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__buf_8_15 sky130_fd_sc_hd__buf_8_15/A sky130_fd_sc_hd__buf_8_15/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_26 sky130_fd_sc_hd__buf_8_26/A sky130_fd_sc_hd__buf_8_26/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_37 sky130_fd_sc_hd__inv_2_91/Y sky130_fd_sc_hd__buf_8_37/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xnor2_1_150 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_150/B sky130_fd_sc_hd__xnor2_1_150/Y
+ sky130_fd_sc_hd__xnor2_1_150/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__buf_8_48 sky130_fd_sc_hd__buf_8_48/A sky130_fd_sc_hd__buf_8_48/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xnor2_1_161 vssd1 vccd1 sky130_fd_sc_hd__o21ai_2_16/Y sky130_fd_sc_hd__xnor2_1_161/Y
+ sky130_fd_sc_hd__xnor2_1_161/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__buf_8_59 sky130_fd_sc_hd__buf_8_59/A sky130_fd_sc_hd__buf_8_59/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xnor2_1_172 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_172/B sky130_fd_sc_hd__inv_2_43/A
+ sky130_fd_sc_hd__xnor2_1_172/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_183 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_183/B sky130_fd_sc_hd__inv_2_46/A
+ sky130_fd_sc_hd__xnor2_1_183/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_194 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_194/B sky130_fd_sc_hd__and2_0_265/A
+ sky130_fd_sc_hd__xnor2_1_194/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_1070 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_501 vssd1 vccd1 sky130_fd_sc_hd__inv_2_38/Y sky130_fd_sc_hd__nand2b_2_3/Y
+ sky130_fd_sc_hd__o21ai_1_501/B1 sky130_fd_sc_hd__xor2_1_301/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1081 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_512 vssd1 vccd1 sky130_fd_sc_hd__inv_2_36/Y sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_512/B1 sky130_fd_sc_hd__xor2_1_311/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1092 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_523 vssd1 vccd1 sky130_fd_sc_hd__inv_2_40/Y sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_523/B1 sky130_fd_sc_hd__xor2_1_322/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_534 vssd1 vccd1 sky130_fd_sc_hd__inv_2_39/Y sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_534/B1 sky130_fd_sc_hd__xor2_1_333/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_545 vssd1 vccd1 sky130_fd_sc_hd__buf_2_10/X sky130_fd_sc_hd__nand2b_1_8/Y
+ sky130_fd_sc_hd__o21ai_1_545/B1 sky130_fd_sc_hd__xor2_1_342/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_556 vssd1 vccd1 sky130_fd_sc_hd__inv_2_28/Y sky130_fd_sc_hd__nand2b_1_9/Y
+ sky130_fd_sc_hd__o21ai_1_556/B1 sky130_fd_sc_hd__xor2_1_354/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_567 vssd1 vccd1 sky130_fd_sc_hd__inv_2_42/Y sky130_fd_sc_hd__nand2_1_422/Y
+ sky130_fd_sc_hd__a21oi_1_87/Y sky130_fd_sc_hd__xnor2_1_102/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_578 vssd1 vccd1 sky130_fd_sc_hd__inv_2_33/Y sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_578/B1 sky130_fd_sc_hd__xor2_1_374/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_589 vssd1 vccd1 sky130_fd_sc_hd__inv_2_27/Y sky130_fd_sc_hd__nand2b_1_9/Y
+ sky130_fd_sc_hd__nand2_1_328/Y sky130_fd_sc_hd__xor2_1_382/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_350 sky130_fd_sc_hd__dfxtp_2_5/Q sky130_fd_sc_hd__xor2_1_350/X
+ sky130_fd_sc_hd__xor2_1_350/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_361 sky130_fd_sc_hd__fa_2_250/A sky130_fd_sc_hd__xor2_1_361/X
+ sky130_fd_sc_hd__xor2_1_361/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_372 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__fah_1_5/A
+ sky130_fd_sc_hd__xor2_1_372/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_383 sky130_fd_sc_hd__xor2_1_383/B sky130_fd_sc_hd__nor2_2_20/B
+ sky130_fd_sc_hd__xor2_1_383/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_394 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__fa_2_271/B
+ sky130_fd_sc_hd__xor2_1_394/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_310 vssd1 vccd1 sky130_fd_sc_hd__buf_2_161/A sky130_fd_sc_hd__buf_8_17/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_321 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_321/X sky130_fd_sc_hd__clkinv_1_901/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_332 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1_12/D sky130_fd_sc_hd__ha_2_23/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_403 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__or2_0_60/A
+ sky130_fd_sc_hd__or2_0_61/A sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__or2_0_61/B
+ sky130_fd_sc_hd__o21ai_1_669/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_343 vssd1 vccd1 sky130_fd_sc_hd__inv_2_3/A sky130_fd_sc_hd__a222oi_1_13/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_414 vccd1 vssd1 sky130_fd_sc_hd__and3_4_23/X sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__buf_8_0/X sky130_fd_sc_hd__nor2_1_178/Y sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__o21ai_1_684/B1 sky130_fd_sc_hd__nor2b_1_15/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_354 vssd1 vccd1 sky130_fd_sc_hd__inv_4_0/A sky130_fd_sc_hd__a222oi_1_2/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_425 vccd1 vssd1 sky130_fd_sc_hd__and3_4_24/X sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__buf_4_7/X sky130_fd_sc_hd__nor2_1_183/Y sky130_fd_sc_hd__buf_4_0/X
+ sky130_fd_sc_hd__o21ai_1_699/B1 sky130_fd_sc_hd__nor2b_1_16/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_436 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__buf_4_5/X sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__o21ai_1_712/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_447 vccd1 vssd1 sky130_fd_sc_hd__and3_4_24/X sky130_fd_sc_hd__or2_0_72/A
+ sky130_fd_sc_hd__or2_0_71/B sky130_fd_sc_hd__nor2_1_183/Y sky130_fd_sc_hd__buf_2_29/X
+ sky130_fd_sc_hd__o21ai_1_726/B1 sky130_fd_sc_hd__nor2b_1_16/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_458 vccd1 vssd1 sky130_fd_sc_hd__and3_4_24/X sky130_fd_sc_hd__or2_0_72/B
+ sky130_fd_sc_hd__or2_0_72/A sky130_fd_sc_hd__nor2_1_183/Y sky130_fd_sc_hd__or2_0_71/B
+ sky130_fd_sc_hd__o21ai_1_740/B1 sky130_fd_sc_hd__nor2b_1_16/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_469 vccd1 vssd1 sky130_fd_sc_hd__and3_4_20/X sky130_fd_sc_hd__buf_2_20/X
+ sky130_fd_sc_hd__buf_2_21/X sky130_fd_sc_hd__nor2_4_16/Y sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__o21ai_1_756/B1 sky130_fd_sc_hd__and2b_4_11/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__dfxtp_1_80 sky130_fd_sc_hd__dfxtp_1_80/Q sky130_fd_sc_hd__dfxtp_1_85/CLK
+ sky130_fd_sc_hd__dfxtp_1_80/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_91 sky130_fd_sc_hd__dfxtp_1_91/Q sky130_fd_sc_hd__dfxtp_1_94/CLK
+ sky130_fd_sc_hd__dfxtp_1_91/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_330 vccd1 vssd1 sky130_fd_sc_hd__and2_0_330/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_330/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_341 vccd1 vssd1 sky130_fd_sc_hd__and2_0_392/A sky130_fd_sc_hd__ha_2_44/SUM
+ sky130_fd_sc_hd__and2_0_342/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_352 vccd1 vssd1 sky130_fd_sc_hd__and2_0_352/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__and2_0_352/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_363 vccd1 vssd1 sky130_fd_sc_hd__and2_0_363/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_68/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_374 vccd1 vssd1 sky130_fd_sc_hd__and2_0_374/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_66/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_385 vccd1 vssd1 sky130_fd_sc_hd__and2_0_385/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_75/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_396 vccd1 vssd1 sky130_fd_sc_hd__and2_0_396/X sky130_fd_sc_hd__and2_0_401/B
+ sky130_fd_sc_hd__and2_0_396/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__conb_1_5 sky130_fd_sc_hd__conb_1_5/LO sky130_fd_sc_hd__conb_1_5/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__inv_2_130 sky130_fd_sc_hd__inv_2_130/A sky130_fd_sc_hd__buf_8_35/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_141 sky130_fd_sc_hd__inv_2_141/A sky130_fd_sc_hd__inv_2_141/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_152 sky130_fd_sc_hd__inv_2_152/A sky130_fd_sc_hd__inv_2_152/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_163 sky130_fd_sc_hd__buf_6_17/X sky130_fd_sc_hd__inv_2_164/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_174 sky130_fd_sc_hd__inv_2_174/A sky130_fd_sc_hd__inv_2_174/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_185 sky130_fd_sc_hd__inv_2_185/A sky130_fd_sc_hd__inv_2_185/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_196 sky130_fd_sc_hd__inv_2_196/A sky130_fd_sc_hd__inv_2_196/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__o22ai_1_104 sky130_fd_sc_hd__xnor2_1_259/Y sky130_fd_sc_hd__xnor2_1_253/Y
+ sky130_fd_sc_hd__ha_2_11/A sky130_fd_sc_hd__inv_2_65/Y sky130_fd_sc_hd__o22ai_1_99/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_115 sky130_fd_sc_hd__xnor2_2_4/Y sky130_fd_sc_hd__xnor2_1_262/Y
+ sky130_fd_sc_hd__fa_2_454/A sky130_fd_sc_hd__xnor2_1_275/Y sky130_fd_sc_hd__o22ai_1_96/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_126 sky130_fd_sc_hd__xnor2_1_288/Y sky130_fd_sc_hd__xnor2_1_274/Y
+ sky130_fd_sc_hd__fa_2_457/B sky130_fd_sc_hd__inv_2_65/Y sky130_fd_sc_hd__o22ai_1_99/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_137 sky130_fd_sc_hd__nor2_4_19/B sky130_fd_sc_hd__nand4_1_0/C
+ sky130_fd_sc_hd__o22ai_1_137/Y sky130_fd_sc_hd__o31ai_2_0/A2 sky130_fd_sc_hd__dfxtp_1_363/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_2_15 sky130_fd_sc_hd__nor2_2_15/B sky130_fd_sc_hd__nor2_2_15/Y
+ sky130_fd_sc_hd__nor2_2_15/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__nor2_2_26 sky130_fd_sc_hd__nor2_2_26/B sky130_fd_sc_hd__nor2_2_26/Y
+ sky130_fd_sc_hd__nor2_2_26/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__o211ai_1_5 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_5/A2
+ sky130_fd_sc_hd__o211ai_1_5/Y sky130_fd_sc_hd__a22oi_1_42/Y sky130_fd_sc_hd__a22oi_1_43/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__a31oi_1_2 vssd1 vccd1 sky130_fd_sc_hd__a31oi_1_2/Y sky130_fd_sc_hd__nor2_1_267/B
+ sky130_fd_sc_hd__nor2_1_273/B sky130_fd_sc_hd__o31ai_1_1/A1 la_data_out[36] vssd1
+ vccd1 sky130_fd_sc_hd__a31oi_1
Xsky130_fd_sc_hd__o21ai_1_320 vssd1 vccd1 sky130_fd_sc_hd__buf_2_5/X sky130_fd_sc_hd__nand2b_2_0/Y
+ sky130_fd_sc_hd__o21ai_1_320/B1 sky130_fd_sc_hd__xor2_1_140/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_331 vssd1 vccd1 sky130_fd_sc_hd__inv_2_21/Y sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__o21ai_1_331/B1 sky130_fd_sc_hd__xor2_1_151/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_342 vssd1 vccd1 sky130_fd_sc_hd__inv_2_17/Y sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__o21ai_1_342/B1 sky130_fd_sc_hd__xor2_1_160/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_353 vssd1 vccd1 sky130_fd_sc_hd__buf_2_3/X sky130_fd_sc_hd__nand2b_2_0/Y
+ sky130_fd_sc_hd__o21ai_1_353/B1 sky130_fd_sc_hd__xor2_1_168/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_364 vssd1 vccd1 sky130_fd_sc_hd__inv_2_17/Y sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__o21ai_1_364/B1 sky130_fd_sc_hd__xor2_1_180/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_375 vssd1 vccd1 sky130_fd_sc_hd__buf_2_2/X sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__o21ai_1_375/B1 sky130_fd_sc_hd__xor2_1_189/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_386 vssd1 vccd1 sky130_fd_sc_hd__inv_2_15/Y sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__o21ai_1_386/B1 sky130_fd_sc_hd__xor2_1_202/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_397 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_296/A sky130_fd_sc_hd__nor2_2_12/Y
+ sky130_fd_sc_hd__nand2_1_378/Y sky130_fd_sc_hd__xnor2_1_82/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_807 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_818 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_702 sky130_fd_sc_hd__xnor2_1_198/A sky130_fd_sc_hd__nand2_1_703/Y
+ sky130_fd_sc_hd__or2_0_81/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_829 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_713 sky130_fd_sc_hd__nand2_1_713/Y sky130_fd_sc_hd__nor2_1_233/B
+ sky130_fd_sc_hd__buf_6_91/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_11 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_11/A1 sky130_fd_sc_hd__buf_4_21/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__or2_0_79/A vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_724 sky130_fd_sc_hd__nand2_1_724/Y sky130_fd_sc_hd__nor2_1_234/A
+ sky130_fd_sc_hd__xor2_1_659/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_22 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_22/A1 sky130_fd_sc_hd__buf_2_80/X
+ sky130_fd_sc_hd__mux2_8_1/S sky130_fd_sc_hd__mux2_2_22/X vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_735 sky130_fd_sc_hd__nand2_1_735/Y sky130_fd_sc_hd__nor2_1_238/A
+ sky130_fd_sc_hd__xor2_1_662/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_33 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_33/A1 sky130_fd_sc_hd__buf_4_12/X
+ sky130_fd_sc_hd__mux2_8_1/S sky130_fd_sc_hd__buf_4_41/A vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_746 sky130_fd_sc_hd__nand2_1_746/Y sky130_fd_sc_hd__or2_0_91/A
+ sky130_fd_sc_hd__or2_0_91/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_44 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_44/A1 sky130_fd_sc_hd__buf_2_83/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__fa_2_415/B vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_757 sky130_fd_sc_hd__xor2_1_661/B sky130_fd_sc_hd__nand2_1_772/Y
+ sky130_fd_sc_hd__nand2_1_757/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_55 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_55/A1 sky130_fd_sc_hd__buf_6_14/X
+ sky130_fd_sc_hd__mux2_8_0/S sky130_fd_sc_hd__mux2_2_55/X vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_768 sky130_fd_sc_hd__xnor2_1_218/B sky130_fd_sc_hd__nand2_1_785/Y
+ sky130_fd_sc_hd__or2_0_97/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_779 sky130_fd_sc_hd__nand2_1_779/Y sky130_fd_sc_hd__or2_0_93/X
+ sky130_fd_sc_hd__or2_0_94/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__conb_1_130 sky130_fd_sc_hd__conb_1_130/LO sky130_fd_sc_hd__conb_1_130/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_141 sky130_fd_sc_hd__conb_1_141/LO sky130_fd_sc_hd__clkinv_1_1/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1806 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1817 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_520 sky130_fd_sc_hd__ha_2_58/A sky130_fd_sc_hd__dfxtp_1_520/CLK
+ sky130_fd_sc_hd__and2_0_357/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_180 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__fa_2_129/B
+ sky130_fd_sc_hd__xor2_1_180/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1828 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_531 wbs_dat_o[10] sky130_fd_sc_hd__dfxtp_1_532/CLK sky130_fd_sc_hd__nor2b_1_147/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_191 sky130_fd_sc_hd__xor2_1_191/B sky130_fd_sc_hd__xor2_1_191/X
+ sky130_fd_sc_hd__xor2_1_191/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1839 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_542 wbs_dat_o[21] sky130_fd_sc_hd__dfxtp_1_544/CLK sky130_fd_sc_hd__nor2b_1_136/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_553 sky130_fd_sc_hd__or2_0_113/A sky130_fd_sc_hd__clkinv_8_75/Y
+ sky130_fd_sc_hd__dfxtp_1_553/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a222oi_1_200 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__buf_4_6/X
+ sky130_fd_sc_hd__buf_4_1/X sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__nor2_2_5/A
+ sky130_fd_sc_hd__o21ai_1_370/B1 sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_140 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_140/X sky130_fd_sc_hd__clkinv_1_874/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_211 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__inv_6_0/Y
+ sky130_fd_sc_hd__buf_8_0/X sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__buf_4_6/X
+ sky130_fd_sc_hd__o21ai_1_386/B1 sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_151 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_12/A1 sky130_fd_sc_hd__clkbuf_1_151/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_222 vccd1 vssd1 sky130_fd_sc_hd__and3_4_17/X sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__buf_4_3/X sky130_fd_sc_hd__nor2_2_20/Y sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__o21ai_1_411/B1 sky130_fd_sc_hd__nor2b_2_4/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_162 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1_931/A sky130_fd_sc_hd__buf_8_67/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_233 vccd1 vssd1 sky130_fd_sc_hd__and3_4_15/X sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__buf_6_1/X sky130_fd_sc_hd__nor2_1_130/Y sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__o21ai_1_427/B1 sky130_fd_sc_hd__nor2b_1_11/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_173 vssd1 vccd1 sky130_fd_sc_hd__a22o_1_30/B2 sky130_fd_sc_hd__clkbuf_1_173/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_244 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__or2_0_60/B
+ sky130_fd_sc_hd__or2_0_60/A sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__or2_0_61/A
+ sky130_fd_sc_hd__o21ai_1_440/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_184 vssd1 vccd1 sky130_fd_sc_hd__buf_12_13/A sky130_fd_sc_hd__clkbuf_1_50/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_255 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__or2_0_61/A
+ sky130_fd_sc_hd__or2_0_42/B sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__or2_0_39/B
+ sky130_fd_sc_hd__o21ai_1_454/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_195 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_195/X sky130_fd_sc_hd__clkbuf_1_60/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_403 sky130_fd_sc_hd__nor2_1_200/A sky130_fd_sc_hd__nor2_1_203/B
+ sky130_fd_sc_hd__fa_2_403/A sky130_fd_sc_hd__fa_2_403/B sky130_fd_sc_hd__fa_2_403/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_266 vccd1 vssd1 sky130_fd_sc_hd__and3_4_13/X sky130_fd_sc_hd__or2_0_52/B
+ sky130_fd_sc_hd__or2_0_53/A sky130_fd_sc_hd__nor2_1_121/Y sky130_fd_sc_hd__buf_2_32/X
+ sky130_fd_sc_hd__o21ai_1_468/B1 sky130_fd_sc_hd__nor2b_1_9/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_414 sky130_fd_sc_hd__fa_2_413/CIN sky130_fd_sc_hd__or2_0_67/A
+ sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__fa_2_414/B sky130_fd_sc_hd__xor2_1_630/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_277 vccd1 vssd1 sky130_fd_sc_hd__and3_4_16/X sky130_fd_sc_hd__buf_2_31/X
+ sky130_fd_sc_hd__buf_2_19/X sky130_fd_sc_hd__nor2_2_19/Y sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__o21ai_1_483/B1 sky130_fd_sc_hd__nor2b_2_3/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_425 sky130_fd_sc_hd__fa_2_422/CIN sky130_fd_sc_hd__fa_2_430/A
+ sky130_fd_sc_hd__fa_2_425/A sky130_fd_sc_hd__fa_2_425/B sky130_fd_sc_hd__ha_2_11/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_288 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__or2_0_66/A sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__or2_0_60/B
+ sky130_fd_sc_hd__o21ai_1_496/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_436 sky130_fd_sc_hd__fa_2_434/A sky130_fd_sc_hd__fa_2_437/A
+ sky130_fd_sc_hd__fa_2_436/A sky130_fd_sc_hd__fa_2_436/B sky130_fd_sc_hd__o22ai_1_77/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_299 vccd1 vssd1 sky130_fd_sc_hd__and3_4_17/X sky130_fd_sc_hd__buf_2_31/X
+ sky130_fd_sc_hd__buf_2_19/X sky130_fd_sc_hd__nor2_2_20/Y sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__o21ai_1_511/B1 sky130_fd_sc_hd__nor2b_2_4/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_447 sky130_fd_sc_hd__fa_2_447/COUT sky130_fd_sc_hd__nor2_1_253/B
+ sky130_fd_sc_hd__fa_2_447/A sky130_fd_sc_hd__fa_2_447/B sky130_fd_sc_hd__fa_2_451/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_458 sky130_fd_sc_hd__fa_2_458/COUT sky130_fd_sc_hd__fa_2_451/A
+ sky130_fd_sc_hd__fa_2_458/A sky130_fd_sc_hd__fa_2_458/B sky130_fd_sc_hd__fa_2_458/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_469 sky130_fd_sc_hd__or2_0_99/B sky130_fd_sc_hd__nor2_1_254/A
+ sky130_fd_sc_hd__fa_2_469/A sky130_fd_sc_hd__fa_2_469/B sky130_fd_sc_hd__nor2b_1_37/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_160 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_74/D sky130_fd_sc_hd__o21ai_2_0/B1
+ sky130_fd_sc_hd__and2_0_160/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_171 vccd1 vssd1 sky130_fd_sc_hd__and2_0_171/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_171/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_182 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_78/D sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__o21ai_1_95/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_90 io_out[11] sky130_fd_sc_hd__conb_1_52/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_193 vccd1 vssd1 sky130_fd_sc_hd__and2_0_193/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__o21ai_1_88/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_12_408 sky130_fd_sc_hd__buf_12_408/A sky130_fd_sc_hd__buf_12_671/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_419 sky130_fd_sc_hd__buf_12_419/A sky130_fd_sc_hd__buf_12_595/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_608 sky130_fd_sc_hd__clkinv_1_608/Y sky130_fd_sc_hd__nand2_1_651/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_619 sky130_fd_sc_hd__nor2_1_188/B sky130_fd_sc_hd__nand2_1_599/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__or2_1_12 sky130_fd_sc_hd__or2_1_12/A sky130_fd_sc_hd__or2_1_12/X
+ sky130_fd_sc_hd__or2_1_12/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_1
Xsky130_fd_sc_hd__o21ai_1_150 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_153/A2 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_142/Y sky130_fd_sc_hd__and2_0_114/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_161 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_21/A sky130_fd_sc_hd__nor2_2_2/Y
+ sky130_fd_sc_hd__nand2_1_174/Y sky130_fd_sc_hd__o21ai_1_161/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_172 vssd1 vccd1 sky130_fd_sc_hd__inv_2_17/Y sky130_fd_sc_hd__nand2b_1_5/Y
+ sky130_fd_sc_hd__a222oi_1_53/Y sky130_fd_sc_hd__xor2_1_5/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_183 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_219/A2 sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__a222oi_1_62/Y sky130_fd_sc_hd__xor2_1_14/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_194 vssd1 vccd1 sky130_fd_sc_hd__buf_2_2/X sky130_fd_sc_hd__nand2b_1_3/Y
+ sky130_fd_sc_hd__a222oi_1_70/Y sky130_fd_sc_hd__xor2_1_23/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_17 vccd1 vssd1 sky130_fd_sc_hd__nand2_1_131/A sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__xor2_1_612/X sky130_fd_sc_hd__xor2_1_187/X sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_17/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_604 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_28 vccd1 vssd1 sky130_fd_sc_hd__xor2_1_313/X sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__inv_2_61/A sky130_fd_sc_hd__xor2_1_100/X sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_28/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_615 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_39 vccd1 vssd1 sky130_fd_sc_hd__nand2_1_127/A sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__xor2_1_602/X sky130_fd_sc_hd__xor2_1_176/X sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_39/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_626 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_510 sky130_fd_sc_hd__nand2_1_510/Y sky130_fd_sc_hd__or2_0_9/A
+ sky130_fd_sc_hd__or2_0_4/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_637 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_521 sky130_fd_sc_hd__nand2_1_521/Y sky130_fd_sc_hd__or2_0_58/A
+ sky130_fd_sc_hd__or2_0_9/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_648 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_532 sky130_fd_sc_hd__nand2_1_532/Y sky130_fd_sc_hd__or2_0_58/B
+ sky130_fd_sc_hd__or2_0_61/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_659 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_19 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_19/B sky130_fd_sc_hd__xnor2_1_19/Y
+ sky130_fd_sc_hd__xnor2_1_19/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_543 sky130_fd_sc_hd__nand2_1_543/Y sky130_fd_sc_hd__or2_0_60/A
+ sky130_fd_sc_hd__or2_0_61/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_554 sky130_fd_sc_hd__nand2_1_554/Y sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__or2_0_60/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_565 sky130_fd_sc_hd__xnor2_1_154/A sky130_fd_sc_hd__nand2_1_566/Y
+ sky130_fd_sc_hd__or2_1_4/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_1 sky130_fd_sc_hd__nor3_2_0/Y sky130_fd_sc_hd__nor2b_1_1/Y
+ sky130_fd_sc_hd__ha_2_8/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nand2_1_576 sky130_fd_sc_hd__nand2_1_576/Y sky130_fd_sc_hd__or2_1_2/A
+ sky130_fd_sc_hd__or2_1_2/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_587 sky130_fd_sc_hd__nand2_1_587/Y sky130_fd_sc_hd__or2_1_3/A
+ sky130_fd_sc_hd__or2_1_3/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_598 sky130_fd_sc_hd__nand2_1_598/Y sky130_fd_sc_hd__nor2_2_29/A
+ sky130_fd_sc_hd__nor2_2_29/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_1101 sky130_fd_sc_hd__nand2_1_866/B wbs_adr_i[6] vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1112 sky130_fd_sc_hd__clkinv_4_55/A sky130_fd_sc_hd__a22o_1_32/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1123 sky130_fd_sc_hd__clkinv_4_66/A sky130_fd_sc_hd__a22o_1_43/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1134 la_data_out[40] sky130_fd_sc_hd__inv_2_92/A vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1145 sky130_fd_sc_hd__clkbuf_4_9/A sky130_fd_sc_hd__inv_4_17/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1603 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1614 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1625 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1636 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1647 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_350 sky130_fd_sc_hd__dfxtp_1_350/Q sky130_fd_sc_hd__dfxtp_1_356/CLK
+ sky130_fd_sc_hd__and2_0_307/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1658 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_361 sky130_fd_sc_hd__a221o_1_0/A2 sky130_fd_sc_hd__dfxtp_1_29/CLK
+ sky130_fd_sc_hd__ha_2_4/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1669 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_372 sky130_fd_sc_hd__dfxtp_1_372/Q sky130_fd_sc_hd__dfxtp_1_375/CLK
+ sky130_fd_sc_hd__nor2b_1_111/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_383 sky130_fd_sc_hd__dfxtp_1_383/Q sky130_fd_sc_hd__dfxtp_1_392/CLK
+ sky130_fd_sc_hd__nor2b_1_100/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_3 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_1_7/B
+ la_data_out[67] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_394 sky130_fd_sc_hd__dfxtp_1_394/Q sky130_fd_sc_hd__dfxtp_1_395/CLK
+ sky130_fd_sc_hd__nor2b_1_88/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_200 sky130_fd_sc_hd__fa_2_192/A sky130_fd_sc_hd__fa_2_199/B
+ sky130_fd_sc_hd__fa_2_200/A sky130_fd_sc_hd__fa_2_200/B sky130_fd_sc_hd__fa_2_200/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_211 sky130_fd_sc_hd__fa_2_204/A sky130_fd_sc_hd__fa_2_210/B
+ sky130_fd_sc_hd__fa_2_211/A sky130_fd_sc_hd__fa_2_211/B sky130_fd_sc_hd__xor2_1_306/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_222 sky130_fd_sc_hd__or2_0_33/A sky130_fd_sc_hd__nor2_1_124/B
+ sky130_fd_sc_hd__fa_2_222/A sky130_fd_sc_hd__fa_2_222/B sky130_fd_sc_hd__fa_2_222/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_233 sky130_fd_sc_hd__fa_2_223/A sky130_fd_sc_hd__fa_2_229/B
+ sky130_fd_sc_hd__fa_2_233/A sky130_fd_sc_hd__fa_2_233/B sky130_fd_sc_hd__xor2_1_334/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_244 sky130_fd_sc_hd__fa_2_236/CIN sky130_fd_sc_hd__fa_2_242/B
+ sky130_fd_sc_hd__fa_2_244/A sky130_fd_sc_hd__fa_2_244/B sky130_fd_sc_hd__xor2_1_351/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_255 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__nor2_1_139/B
+ sky130_fd_sc_hd__fa_2_255/A sky130_fd_sc_hd__fa_2_255/B sky130_fd_sc_hd__fa_2_255/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_266 sky130_fd_sc_hd__nor2_1_145/A sky130_fd_sc_hd__nor2_1_147/B
+ sky130_fd_sc_hd__fa_2_266/A sky130_fd_sc_hd__fa_2_266/B sky130_fd_sc_hd__fa_2_266/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_277 sky130_fd_sc_hd__fa_2_275/CIN sky130_fd_sc_hd__fa_2_278/A
+ sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__fa_2_277/B sky130_fd_sc_hd__xor2_1_408/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_288 sky130_fd_sc_hd__xor3_1_28/A sky130_fd_sc_hd__fa_2_285/B
+ sky130_fd_sc_hd__ha_2_2/SUM sky130_fd_sc_hd__fa_2_288/B sky130_fd_sc_hd__fa_2_288/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_4 vccd1 vssd1 sky130_fd_sc_hd__and2_0_4/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_4/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__fa_2_299 sky130_fd_sc_hd__or2_1_9/A sky130_fd_sc_hd__nor2_2_22/A
+ sky130_fd_sc_hd__fa_2_299/A sky130_fd_sc_hd__fa_2_299/B sky130_fd_sc_hd__fa_2_299/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_80 sky130_fd_sc_hd__or2_0_6/A sky130_fd_sc_hd__nor2_1_65/B
+ sky130_fd_sc_hd__fa_2_80/A sky130_fd_sc_hd__fa_2_80/B sky130_fd_sc_hd__fa_2_80/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_91 sky130_fd_sc_hd__fa_2_81/A sky130_fd_sc_hd__fa_2_87/B sky130_fd_sc_hd__fa_2_91/A
+ sky130_fd_sc_hd__fa_2_91/B sky130_fd_sc_hd__fa_2_91/CIN vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a21oi_1_30 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_59/Y
+ sky130_fd_sc_hd__a21oi_1_30/Y sky130_fd_sc_hd__dfxtp_1_67/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_41 sky130_fd_sc_hd__a21oi_1_45/A1 sky130_fd_sc_hd__o21ai_1_209/Y
+ sky130_fd_sc_hd__a21oi_1_41/Y sky130_fd_sc_hd__nor2_1_51/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_205 sky130_fd_sc_hd__buf_6_82/X sky130_fd_sc_hd__buf_12_381/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_52 sky130_fd_sc_hd__a21oi_1_54/A1 sky130_fd_sc_hd__nand2_1_250/Y
+ sky130_fd_sc_hd__a21oi_1_52/Y sky130_fd_sc_hd__nor2_1_78/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_216 sky130_fd_sc_hd__buf_6_34/X sky130_fd_sc_hd__buf_12_453/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_63 sky130_fd_sc_hd__xnor2_1_56/B sky130_fd_sc_hd__a21oi_1_63/B1
+ sky130_fd_sc_hd__xnor2_1_2/A sky130_fd_sc_hd__nand2_1_302/A vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_227 sky130_fd_sc_hd__buf_6_27/X sky130_fd_sc_hd__buf_12_418/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_74 sky130_fd_sc_hd__a21oi_1_74/A1 sky130_fd_sc_hd__nor2_1_106/A
+ sky130_fd_sc_hd__a21oi_1_74/Y sky130_fd_sc_hd__or2_0_38/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_238 sky130_fd_sc_hd__buf_6_62/X sky130_fd_sc_hd__buf_12_351/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_85 sky130_fd_sc_hd__o21ai_1_570/Y sky130_fd_sc_hd__a21oi_1_85/B1
+ sky130_fd_sc_hd__a21oi_1_85/Y sky130_fd_sc_hd__or2_1_0/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_249 sky130_fd_sc_hd__buf_6_48/X sky130_fd_sc_hd__buf_12_344/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_96 sky130_fd_sc_hd__or2_0_43/X sky130_fd_sc_hd__a21oi_1_96/B1
+ sky130_fd_sc_hd__xor2_1_403/B sky130_fd_sc_hd__xnor2_1_117/A vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_1_108 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_178/Q sky130_fd_sc_hd__dfxtp_1_146/Q sky130_fd_sc_hd__o21ai_1_14/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_119 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_167/Q sky130_fd_sc_hd__dfxtp_1_135/Q sky130_fd_sc_hd__o21ai_1_25/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor3_1_0 sky130_fd_sc_hd__nor3_1_0/C sky130_fd_sc_hd__nor3_1_0/Y
+ sky130_fd_sc_hd__nor3_1_0/A sky130_fd_sc_hd__nor3_1_0/B vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__clkinv_1_405 sky130_fd_sc_hd__nand2_1_317/A sky130_fd_sc_hd__o21a_1_1/A2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_416 sky130_fd_sc_hd__nor2_1_106/B sky130_fd_sc_hd__nand2_1_343/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_427 sky130_fd_sc_hd__o21ai_1_444/A2 sky130_fd_sc_hd__o21ai_1_456/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_438 sky130_fd_sc_hd__a21oi_1_79/B1 sky130_fd_sc_hd__nor2_1_119/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_449 sky130_fd_sc_hd__nor2_1_122/B sky130_fd_sc_hd__nand2_1_387/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_70 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_81 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_92 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_70 vccd1 vssd1 sky130_fd_sc_hd__buf_6_70/X sky130_fd_sc_hd__buf_8_50/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_81 vccd1 vssd1 sky130_fd_sc_hd__buf_6_81/X sky130_fd_sc_hd__buf_6_81/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_92 vccd1 vssd1 sky130_fd_sc_hd__buf_6_92/X sky130_fd_sc_hd__buf_6_92/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_50 sky130_fd_sc_hd__buf_2_189/A vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_61 sky130_fd_sc_hd__dfxtp_1_12/Q vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a222oi_1_5 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_346/Q sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__o211ai_1_21/Y sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__a222oi_1_5/Y sky130_fd_sc_hd__dfxtp_1_297/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_401 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_412 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_423 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_434 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_445 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_456 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_340 sky130_fd_sc_hd__nand2_1_340/Y sky130_fd_sc_hd__nor2_1_108/Y
+ sky130_fd_sc_hd__nand2_1_374/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_467 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_351 sky130_fd_sc_hd__nand2_1_351/Y sky130_fd_sc_hd__or2_0_28/A
+ sky130_fd_sc_hd__or2_0_28/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_478 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_950 sky130_fd_sc_hd__clkbuf_1_60/A sky130_fd_sc_hd__clkinv_4_20/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_362 sky130_fd_sc_hd__nand2_1_362/Y sky130_fd_sc_hd__or2_0_29/A
+ sky130_fd_sc_hd__or2_0_29/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_489 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_961 sky130_fd_sc_hd__buf_2_157/A sky130_fd_sc_hd__clkinv_1_961/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_373 sky130_fd_sc_hd__nand2_1_373/Y sky130_fd_sc_hd__or2_0_30/A
+ sky130_fd_sc_hd__or2_0_30/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_972 sky130_fd_sc_hd__clkinv_1_972/Y sky130_fd_sc_hd__clkinv_4_23/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_384 sky130_fd_sc_hd__nand2_1_384/Y sky130_fd_sc_hd__or2_0_33/A
+ sky130_fd_sc_hd__or2_0_33/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_983 sky130_fd_sc_hd__clkinv_1_983/Y sky130_fd_sc_hd__clkinv_4_27/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_395 sky130_fd_sc_hd__nand2_1_395/Y sky130_fd_sc_hd__or2_0_44/X
+ sky130_fd_sc_hd__nor2_1_128/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_994 sky130_fd_sc_hd__clkinv_1_994/Y sky130_fd_sc_hd__clkinv_1_994/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1400 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1411 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1422 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1433 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1444 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1455 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1466 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1477 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_180 sky130_fd_sc_hd__dfxtp_1_180/Q sky130_fd_sc_hd__clkinv_4_2/Y
+ sky130_fd_sc_hd__and2_0_207/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_908 vssd1 vccd1 sky130_fd_sc_hd__o31ai_1_0/A1 sky130_fd_sc_hd__nor2_1_277/Y
+ sky130_fd_sc_hd__o21ai_2_18/A1 sky130_fd_sc_hd__o21ai_1_908/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1488 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_191 sky130_fd_sc_hd__dfxtp_1_191/Q sky130_fd_sc_hd__dfxtp_4_3/CLK
+ sky130_fd_sc_hd__and2_0_9/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_919 vssd1 vccd1 sky130_fd_sc_hd__ha_2_58/SUM sky130_fd_sc_hd__o21ai_1_919/A1
+ sky130_fd_sc_hd__a21oi_1_195/Y sky130_fd_sc_hd__o21ai_1_919/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1499 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_17 vccd1 vssd1 sky130_fd_sc_hd__buf_2_17/X sky130_fd_sc_hd__nor2_1_1/Y
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_28 vccd1 vssd1 sky130_fd_sc_hd__or2_0_72/B sky130_fd_sc_hd__buf_2_28/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_39 vccd1 vssd1 sky130_fd_sc_hd__buf_2_39/X sky130_fd_sc_hd__buf_2_39/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_990 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o211ai_1_11 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_52/B1
+ sky130_fd_sc_hd__a22oi_1_8/A2 sky130_fd_sc_hd__a22oi_1_54/Y sky130_fd_sc_hd__a22oi_1_55/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_22 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_41/B1
+ sky130_fd_sc_hd__o211ai_1_22/Y sky130_fd_sc_hd__a22oi_1_76/Y sky130_fd_sc_hd__a22oi_1_77/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_33 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o21ai_1_3/A2
+ sky130_fd_sc_hd__fa_2_301/A sky130_fd_sc_hd__nand2_1_53/Y sky130_fd_sc_hd__a21oi_1_4/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_44 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o22ai_1_19/B1
+ sky130_fd_sc_hd__fa_2_372/A sky130_fd_sc_hd__nand2_1_64/Y sky130_fd_sc_hd__a21oi_1_15/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_55 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o22ai_1_8/B1
+ sky130_fd_sc_hd__fa_2_406/A sky130_fd_sc_hd__nand2_1_75/Y sky130_fd_sc_hd__a21oi_1_26/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__clkinv_1_202 sky130_fd_sc_hd__o22ai_1_49/B1 sky130_fd_sc_hd__dfxtp_1_173/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_213 sky130_fd_sc_hd__o22ai_1_11/B1 sky130_fd_sc_hd__dfxtp_1_106/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_224 sky130_fd_sc_hd__nor2_1_11/A sky130_fd_sc_hd__dfxtp_1_134/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_235 sky130_fd_sc_hd__o22ai_1_3/A2 sky130_fd_sc_hd__dfxtp_1_162/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_246 sky130_fd_sc_hd__o22ai_1_2/B1 sky130_fd_sc_hd__dfxtp_1_97/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_257 sky130_fd_sc_hd__o21ai_1_117/A2 sky130_fd_sc_hd__xor2_1_597/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_268 sky130_fd_sc_hd__nand2_1_147/A sky130_fd_sc_hd__ha_2_9/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_279 sky130_fd_sc_hd__and2_0_120/A sky130_fd_sc_hd__a222oi_1_23/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_2_2 sky130_fd_sc_hd__buf_2_16/A sky130_fd_sc_hd__o21ai_2_2/Y
+ sky130_fd_sc_hd__o21ai_2_4/A2 sky130_fd_sc_hd__o21ai_2_2/A1 vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__o21ai_2
Xsky130_fd_sc_hd__xor3_1_8 sky130_fd_sc_hd__xor3_1_8/X sky130_fd_sc_hd__xor3_1_8/C
+ sky130_fd_sc_hd__xor3_1_8/B sky130_fd_sc_hd__xor3_1_8/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__a21oi_1_9 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_38/Y
+ sky130_fd_sc_hd__a21oi_1_9/Y sky130_fd_sc_hd__dfxtp_1_87/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__and3_4_15 sky130_fd_sc_hd__and3_4_15/A sky130_fd_sc_hd__and3_4_15/B
+ sky130_fd_sc_hd__and3_4_15/C sky130_fd_sc_hd__and3_4_15/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__and3_4_26 sky130_fd_sc_hd__nor2_2_31/B sky130_fd_sc_hd__and3_4_26/B
+ sky130_fd_sc_hd__nor2_2_31/A sky130_fd_sc_hd__and3_4_26/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__a21oi_1_110 sky130_fd_sc_hd__clkinv_1_549/Y sky130_fd_sc_hd__o21ai_1_673/Y
+ sky130_fd_sc_hd__a21oi_1_110/Y sky130_fd_sc_hd__nor2_1_169/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_121 sky130_fd_sc_hd__clkinv_1_580/Y sky130_fd_sc_hd__o21ai_1_799/Y
+ sky130_fd_sc_hd__a21oi_1_121/Y sky130_fd_sc_hd__nor2_1_190/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_132 sky130_fd_sc_hd__xnor2_1_181/B sky130_fd_sc_hd__nand2_1_635/Y
+ sky130_fd_sc_hd__xnor2_1_127/A sky130_fd_sc_hd__nor2_1_213/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_143 sky130_fd_sc_hd__xnor2_1_193/B sky130_fd_sc_hd__clkinv_1_635/Y
+ sky130_fd_sc_hd__xor2_1_644/A sky130_fd_sc_hd__or2_0_77/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_154 sky130_fd_sc_hd__or2_0_90/X sky130_fd_sc_hd__clkinv_1_668/Y
+ sky130_fd_sc_hd__a21oi_1_154/Y sky130_fd_sc_hd__clkinv_1_669/Y vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_165 sky130_fd_sc_hd__or2_0_94/X sky130_fd_sc_hd__clkinv_1_694/Y
+ sky130_fd_sc_hd__a21oi_1_165/Y sky130_fd_sc_hd__clkinv_1_695/Y vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_176 sky130_fd_sc_hd__xnor2_1_297/B sky130_fd_sc_hd__clkinv_1_820/Y
+ sky130_fd_sc_hd__xor2_1_682/A sky130_fd_sc_hd__or2_0_106/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_187 sky130_fd_sc_hd__nor2_1_273/Y sky130_fd_sc_hd__nor2_4_0/A
+ sky130_fd_sc_hd__a21oi_1_187/Y sky130_fd_sc_hd__nor2_1_278/B vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_198 sky130_fd_sc_hd__ha_2_58/SUM sky130_fd_sc_hd__ha_2_58/COUT
+ sky130_fd_sc_hd__nand2_1_860/A sky130_fd_sc_hd__o21ai_1_919/A1 vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_106 sky130_fd_sc_hd__buf_12_9/X sky130_fd_sc_hd__buf_8_106/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_117 sky130_fd_sc_hd__buf_8_117/A sky130_fd_sc_hd__buf_6_84/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_128 sky130_fd_sc_hd__buf_8_128/A sky130_fd_sc_hd__buf_6_77/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_139 sky130_fd_sc_hd__buf_8_73/A sky130_fd_sc_hd__buf_8_139/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_12_580 sky130_fd_sc_hd__buf_12_580/A sky130_fd_sc_hd__buf_12_580/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_591 sky130_fd_sc_hd__buf_12_591/A sky130_fd_sc_hd__buf_12_591/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_220 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_231 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_242 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_253 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_264 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_275 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_310 vssd1 vccd1 sky130_fd_sc_hd__maj3_1_3/A sky130_fd_sc_hd__nand4_1_3/B
+ la_data_out[50] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_286 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_170 sky130_fd_sc_hd__nor2_1_47/A sky130_fd_sc_hd__or2_0_10/X
+ sky130_fd_sc_hd__nand2_1_170/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_297 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_181 sky130_fd_sc_hd__nand2_1_181/Y sky130_fd_sc_hd__nor2_1_51/Y
+ sky130_fd_sc_hd__nand2_1_203/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_780 sky130_fd_sc_hd__and2_0_327/A sky130_fd_sc_hd__clkinv_1_780/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_192 sky130_fd_sc_hd__nand2_1_192/Y sky130_fd_sc_hd__nor2_1_57/Y
+ sky130_fd_sc_hd__nand2_1_203/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_791 sky130_fd_sc_hd__and2_0_316/A sky130_fd_sc_hd__clkinv_1_791/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1230 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1241 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1252 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1263 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1274 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_705 vssd1 vccd1 sky130_fd_sc_hd__buf_2_13/X sky130_fd_sc_hd__nand2b_1_19/Y
+ sky130_fd_sc_hd__o21ai_1_705/B1 sky130_fd_sc_hd__xor2_1_484/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1285 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_716 vssd1 vccd1 sky130_fd_sc_hd__buf_2_12/X sky130_fd_sc_hd__nand2b_1_21/Y
+ sky130_fd_sc_hd__o21ai_1_716/B1 sky130_fd_sc_hd__xor2_1_493/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1296 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_727 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_861/A2 sky130_fd_sc_hd__nand2b_1_19/Y
+ sky130_fd_sc_hd__nand2_1_494/Y sky130_fd_sc_hd__xor2_1_503/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_738 vssd1 vccd1 sky130_fd_sc_hd__xor2_2_2/X sky130_fd_sc_hd__nand2b_2_6/Y
+ sky130_fd_sc_hd__o21ai_1_738/B1 sky130_fd_sc_hd__xor2_1_514/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_749 vssd1 vccd1 sky130_fd_sc_hd__inv_2_50/Y sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__o21ai_1_749/B1 sky130_fd_sc_hd__xor2_1_524/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_12 sky130_fd_sc_hd__fa_2_56/A sky130_fd_sc_hd__fa_2_7/B sky130_fd_sc_hd__xor2_1_12/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_23 sky130_fd_sc_hd__fa_2_28/A sky130_fd_sc_hd__xor2_1_23/X
+ sky130_fd_sc_hd__xor2_1_23/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_34 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__fa_2_20/A
+ sky130_fd_sc_hd__xor2_1_34/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_45 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__fa_2_27/A
+ sky130_fd_sc_hd__xor2_1_45/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_56 sky130_fd_sc_hd__xor2_1_9/B sky130_fd_sc_hd__fa_2_38/A
+ sky130_fd_sc_hd__xor2_1_56/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_67 sky130_fd_sc_hd__fa_2_97/A sky130_fd_sc_hd__xor2_1_67/X
+ sky130_fd_sc_hd__xor2_1_67/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_78 sky130_fd_sc_hd__fa_2_56/A sky130_fd_sc_hd__and3_4_4/A
+ sky130_fd_sc_hd__xor2_1_78/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_89 sky130_fd_sc_hd__xor2_1_9/B sky130_fd_sc_hd__xor2_1_89/X
+ sky130_fd_sc_hd__xor2_1_89/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2b_1_6 sky130_fd_sc_hd__nand2b_1_6/Y sky130_fd_sc_hd__and3_4_6/C
+ sky130_fd_sc_hd__and3_4_6/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a21o_2_2 sky130_fd_sc_hd__a21o_2_2/X sky130_fd_sc_hd__a21o_2_2/B1
+ wbs_adr_i[5] sky130_fd_sc_hd__or3_1_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__xor2_1_510 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__xor2_1_510/X
+ sky130_fd_sc_hd__xor2_1_510/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_521 sky130_fd_sc_hd__fa_2_357/A sky130_fd_sc_hd__fa_2_354/B
+ sky130_fd_sc_hd__xor2_1_521/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_532 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__xor2_1_532/X
+ sky130_fd_sc_hd__xor2_1_532/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_543 sky130_fd_sc_hd__xor2_1_543/B sky130_fd_sc_hd__xor2_1_543/X
+ sky130_fd_sc_hd__xor2_1_543/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_554 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__xor2_1_554/X
+ sky130_fd_sc_hd__xor2_1_554/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_565 sky130_fd_sc_hd__fah_1_14/A sky130_fd_sc_hd__fah_1_11/A
+ sky130_fd_sc_hd__xor2_1_565/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_576 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__fa_2_390/A
+ sky130_fd_sc_hd__xor2_1_576/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_587 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__fa_2_397/B
+ sky130_fd_sc_hd__xor2_1_587/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_598 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__xor2_1_598/X
+ sky130_fd_sc_hd__xor2_1_598/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a222oi_1_607 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_393/Q sky130_fd_sc_hd__and2b_4_13/X
+ sky130_fd_sc_hd__nor2_4_19/Y sky130_fd_sc_hd__dfxtp_1_457/Q sky130_fd_sc_hd__nor2_4_19/B
+ sky130_fd_sc_hd__clkinv_1_804/A sky130_fd_sc_hd__dfxtp_1_425/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__and2b_4_1 sky130_fd_sc_hd__or2b_2_0/A sky130_fd_sc_hd__and2b_4_1/X
+ sky130_fd_sc_hd__and3_4_0/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__and2b_4
Xsky130_fd_sc_hd__ha_2_50 vssd1 vccd1 sky130_fd_sc_hd__ha_2_50/A sky130_fd_sc_hd__ha_2_52/B
+ sky130_fd_sc_hd__ha_2_50/SUM sky130_fd_sc_hd__ha_2_50/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_2 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_2/X sky130_fd_sc_hd__xnor2_1_0/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a221o_1_0 sky130_fd_sc_hd__nor3b_1_0/B sky130_fd_sc_hd__a221o_1_0/B1
+ sky130_fd_sc_hd__a221o_1_0/A1 sky130_fd_sc_hd__a221o_1_0/B2 sky130_fd_sc_hd__a221o_1_0/A2
+ vssd1 vccd1 sky130_fd_sc_hd__a221o_1_0/C1 vssd1 vccd1 sky130_fd_sc_hd__a221o_1
Xsky130_fd_sc_hd__clkinv_1_2 la_data_out[125] sky130_fd_sc_hd__clkinv_1_2/A vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_170 sky130_fd_sc_hd__nor2_1_170/B sky130_fd_sc_hd__nor2_1_170/Y
+ sky130_fd_sc_hd__nor2_1_173/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_181 sky130_fd_sc_hd__nor2_1_181/B sky130_fd_sc_hd__nor2_1_181/Y
+ sky130_fd_sc_hd__nor2_1_181/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_192 sky130_fd_sc_hd__nor2_1_194/Y sky130_fd_sc_hd__nor2_1_192/Y
+ sky130_fd_sc_hd__nor2_1_198/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_90 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__nor2_4_3/Y
+ sky130_fd_sc_hd__nand2_1_52/B sky130_fd_sc_hd__dfxtp_1_156/Q sky130_fd_sc_hd__a22oi_1_90/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__and2_0_17 vccd1 vssd1 sky130_fd_sc_hd__and2_0_17/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__buf_6_2/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_28 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_4_0/D sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__buf_2_26/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_39 vccd1 vssd1 sky130_fd_sc_hd__and2_0_39/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__buf_6_1/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nor2_2_9 sky130_fd_sc_hd__nor2_2_9/B sky130_fd_sc_hd__nor2_2_9/Y
+ sky130_fd_sc_hd__nor2_2_9/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__buf_8_16 sky130_fd_sc_hd__buf_8_16/A sky130_fd_sc_hd__buf_8_16/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_27 sky130_fd_sc_hd__buf_8_27/A sky130_fd_sc_hd__buf_8_27/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xnor2_1_140 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_140/B sky130_fd_sc_hd__and3_1_2/C
+ sky130_fd_sc_hd__fa_2_338/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__buf_8_38 sky130_fd_sc_hd__inv_2_79/Y sky130_fd_sc_hd__buf_8_38/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xnor2_1_151 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_530/A sky130_fd_sc_hd__and3_4_24/B
+ sky130_fd_sc_hd__xnor2_1_153/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__buf_8_49 sky130_fd_sc_hd__buf_8_49/A sky130_fd_sc_hd__buf_8_49/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xnor2_1_162 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_575/A sky130_fd_sc_hd__and3_4_26/B
+ sky130_fd_sc_hd__xnor2_1_164/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_173 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_609/A sky130_fd_sc_hd__and3_4_20/C
+ sky130_fd_sc_hd__xnor2_1_176/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_184 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_186/A sky130_fd_sc_hd__and3_4_22/C
+ sky130_fd_sc_hd__xor2_1_631/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_195 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_195/B sky130_fd_sc_hd__and2_0_263/A
+ sky130_fd_sc_hd__xnor2_1_195/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_4_90 wbs_dat_i[7] sky130_fd_sc_hd__clkinv_4_90/Y vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_1060 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1071 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_502 vssd1 vccd1 sky130_fd_sc_hd__inv_2_30/Y sky130_fd_sc_hd__nand2b_1_9/Y
+ sky130_fd_sc_hd__o21ai_1_502/B1 sky130_fd_sc_hd__xor2_1_302/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1082 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_513 vssd1 vccd1 sky130_fd_sc_hd__inv_2_39/Y sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_513/B1 sky130_fd_sc_hd__xor2_1_312/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1093 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_524 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_0/Y sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_524/B1 sky130_fd_sc_hd__xor2_1_323/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_535 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_7/X sky130_fd_sc_hd__nor2_1_126/B
+ sky130_fd_sc_hd__o21ai_1_535/B1 sky130_fd_sc_hd__xnor2_1_93/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_546 vssd1 vccd1 sky130_fd_sc_hd__inv_2_27/Y sky130_fd_sc_hd__nand2b_1_14/Y
+ sky130_fd_sc_hd__nand2_1_326/Y sky130_fd_sc_hd__xor2_1_343/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_557 vssd1 vccd1 sky130_fd_sc_hd__nand2_2_12/Y sky130_fd_sc_hd__nand2b_1_8/Y
+ sky130_fd_sc_hd__a22oi_1_207/Y sky130_fd_sc_hd__xor2_1_355/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_568 vssd1 vccd1 sky130_fd_sc_hd__buf_2_11/X sky130_fd_sc_hd__nand2b_2_3/Y
+ sky130_fd_sc_hd__o21ai_1_568/B1 sky130_fd_sc_hd__xor2_1_365/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_579 vssd1 vccd1 sky130_fd_sc_hd__inv_2_42/Y sky130_fd_sc_hd__nor2_1_132/B
+ sky130_fd_sc_hd__a21oi_1_92/Y sky130_fd_sc_hd__xnor2_1_105/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_340 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__fa_2_237/A
+ sky130_fd_sc_hd__xor2_1_340/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_351 sky130_fd_sc_hd__fa_2_250/A sky130_fd_sc_hd__xor2_1_351/X
+ sky130_fd_sc_hd__xor2_1_351/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_362 sky130_fd_sc_hd__xor2_1_362/B sky130_fd_sc_hd__nor2_2_19/B
+ sky130_fd_sc_hd__xor2_1_362/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_373 sky130_fd_sc_hd__fa_2_281/A sky130_fd_sc_hd__xor2_1_373/X
+ sky130_fd_sc_hd__xor2_1_373/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_384 sky130_fd_sc_hd__xor2_1_384/B sky130_fd_sc_hd__xor2_1_384/X
+ sky130_fd_sc_hd__xor2_1_384/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_395 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__xor2_1_395/X
+ sky130_fd_sc_hd__xor2_1_395/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_300 vssd1 vccd1 sky130_fd_sc_hd__bufinv_8_0/A sky130_fd_sc_hd__inv_2_191/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_311 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_311/X sky130_fd_sc_hd__clkinv_1_870/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_322 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_322/X sky130_fd_sc_hd__clkinv_1_903/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_333 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1_14/D sky130_fd_sc_hd__ha_2_24/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_404 vccd1 vssd1 sky130_fd_sc_hd__and3_4_20/X sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__buf_4_2/X sky130_fd_sc_hd__nor2_4_16/Y sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__o21ai_1_670/B1 sky130_fd_sc_hd__and2b_4_11/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_344 vssd1 vccd1 sky130_fd_sc_hd__inv_4_6/A sky130_fd_sc_hd__a222oi_1_12/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_415 vccd1 vssd1 sky130_fd_sc_hd__and3_4_18/X sky130_fd_sc_hd__nor2_2_10/B
+ sky130_fd_sc_hd__buf_6_4/X sky130_fd_sc_hd__nor2_2_32/Y sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__o21ai_1_686/B1 sky130_fd_sc_hd__nor2b_2_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_355 vssd1 vccd1 sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__a222oi_1_1/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_426 vccd1 vssd1 sky130_fd_sc_hd__and3_4_25/X sky130_fd_sc_hd__buf_2_27/X
+ sky130_fd_sc_hd__buf_2_15/X sky130_fd_sc_hd__nor2_1_186/Y sky130_fd_sc_hd__buf_2_4/A
+ sky130_fd_sc_hd__o21ai_1_700/B1 sky130_fd_sc_hd__nor2b_1_17/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_437 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__or2_0_60/B
+ sky130_fd_sc_hd__or2_0_60/A sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__or2_0_61/A
+ sky130_fd_sc_hd__o21ai_1_713/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_448 vccd1 vssd1 sky130_fd_sc_hd__and3_4_18/X sky130_fd_sc_hd__buf_2_20/X
+ sky130_fd_sc_hd__buf_2_21/X sky130_fd_sc_hd__nor2_2_32/Y sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__o21ai_1_728/B1 sky130_fd_sc_hd__nor2b_2_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_459 vccd1 vssd1 sky130_fd_sc_hd__and3_4_25/X sky130_fd_sc_hd__buf_2_29/X
+ sky130_fd_sc_hd__buf_2_30/X sky130_fd_sc_hd__nor2_1_186/Y sky130_fd_sc_hd__buf_2_26/X
+ sky130_fd_sc_hd__o21ai_1_741/B1 sky130_fd_sc_hd__nor2b_1_17/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__dfxtp_1_70 sky130_fd_sc_hd__dfxtp_1_70/Q sky130_fd_sc_hd__dfxtp_1_72/CLK
+ sky130_fd_sc_hd__dfxtp_1_70/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_81 sky130_fd_sc_hd__dfxtp_1_81/Q sky130_fd_sc_hd__dfxtp_1_81/CLK
+ sky130_fd_sc_hd__dfxtp_1_81/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_92 sky130_fd_sc_hd__dfxtp_1_92/Q sky130_fd_sc_hd__dfxtp_1_94/CLK
+ sky130_fd_sc_hd__and2_0_7/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_320 vccd1 vssd1 sky130_fd_sc_hd__and2_0_320/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_320/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_331 vccd1 vssd1 sky130_fd_sc_hd__and2_0_331/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_331/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_342 vccd1 vssd1 sky130_fd_sc_hd__and2_0_390/A sky130_fd_sc_hd__ha_2_43/SUM
+ sky130_fd_sc_hd__and2_0_342/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_353 vccd1 vssd1 sky130_fd_sc_hd__and2_0_353/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__buf_2_46/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_364 vccd1 vssd1 sky130_fd_sc_hd__and2_0_364/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_62/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_375 vccd1 vssd1 sky130_fd_sc_hd__and2_0_375/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_69/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_386 vccd1 vssd1 sky130_fd_sc_hd__and2_0_386/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_77/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_397 vccd1 vssd1 sky130_fd_sc_hd__and2_0_397/X sky130_fd_sc_hd__and2_0_401/B
+ sky130_fd_sc_hd__and2_0_397/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__conb_1_6 sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__conb_1_6/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__or2_0_0 sky130_fd_sc_hd__or2_0_0/A sky130_fd_sc_hd__or2_0_0/X sky130_fd_sc_hd__or2_0_0/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__inv_2_120 sky130_fd_sc_hd__inv_2_120/A sky130_fd_sc_hd__buf_6_19/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_131 sky130_fd_sc_hd__inv_4_11/Y sky130_fd_sc_hd__buf_8_36/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_142 sky130_fd_sc_hd__buf_8_98/A sky130_fd_sc_hd__inv_2_143/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_153 sky130_fd_sc_hd__inv_2_153/A sky130_fd_sc_hd__inv_2_153/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_164 sky130_fd_sc_hd__inv_2_164/A sky130_fd_sc_hd__inv_2_164/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_175 sky130_fd_sc_hd__inv_2_175/A sky130_fd_sc_hd__buf_8_70/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_186 sky130_fd_sc_hd__inv_2_186/A sky130_fd_sc_hd__inv_2_186/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_197 sky130_fd_sc_hd__inv_2_94/A sky130_fd_sc_hd__inv_2_197/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__o22ai_1_105 sky130_fd_sc_hd__xnor2_2_4/Y sky130_fd_sc_hd__xnor2_1_254/Y
+ sky130_fd_sc_hd__fa_2_429/A sky130_fd_sc_hd__xnor2_1_261/Y sky130_fd_sc_hd__o22ai_1_96/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_116 sky130_fd_sc_hd__xnor2_2_4/Y sky130_fd_sc_hd__xnor2_1_261/Y
+ sky130_fd_sc_hd__fa_2_449/CIN sky130_fd_sc_hd__xnor2_1_262/Y sky130_fd_sc_hd__o22ai_1_96/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_127 sky130_fd_sc_hd__xnor2_2_4/Y sky130_fd_sc_hd__xnor2_1_275/Y
+ sky130_fd_sc_hd__fa_2_458/CIN sky130_fd_sc_hd__xnor2_1_284/Y sky130_fd_sc_hd__o22ai_1_96/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_138 sky130_fd_sc_hd__dfxtp_1_358/Q sky130_fd_sc_hd__ha_2_9/B
+ sky130_fd_sc_hd__o22ai_1_138/Y sky130_fd_sc_hd__nand4_1_0/B sky130_fd_sc_hd__nor2_4_19/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_2_16 sky130_fd_sc_hd__buf_2_31/X sky130_fd_sc_hd__nor2_2_16/Y
+ sky130_fd_sc_hd__buf_2_23/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__nor2_2_27 sky130_fd_sc_hd__nor2_2_27/B sky130_fd_sc_hd__nor2_2_27/Y
+ sky130_fd_sc_hd__nor2_2_27/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__o211ai_1_6 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_6/A2
+ sky130_fd_sc_hd__o211ai_1_6/Y sky130_fd_sc_hd__a22oi_1_44/Y sky130_fd_sc_hd__a22oi_1_45/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o21ai_1_310 vssd1 vccd1 sky130_fd_sc_hd__buf_2_3/X sky130_fd_sc_hd__nand2b_1_7/Y
+ sky130_fd_sc_hd__o21ai_1_310/B1 sky130_fd_sc_hd__xor2_1_129/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_321 vssd1 vccd1 sky130_fd_sc_hd__inv_2_15/Y sky130_fd_sc_hd__nand2b_1_1/Y
+ sky130_fd_sc_hd__o21ai_1_321/B1 sky130_fd_sc_hd__xor2_1_141/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_332 vssd1 vccd1 sky130_fd_sc_hd__inv_2_11/Y sky130_fd_sc_hd__nand2_1_251/Y
+ sky130_fd_sc_hd__a21oi_1_52/Y sky130_fd_sc_hd__xnor2_1_39/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_343 vssd1 vccd1 sky130_fd_sc_hd__inv_2_12/Y sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__o21ai_1_343/B1 sky130_fd_sc_hd__xor2_1_161/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_354 vssd1 vccd1 sky130_fd_sc_hd__inv_2_26/Y sky130_fd_sc_hd__nand2b_1_1/Y
+ sky130_fd_sc_hd__nand2_1_158/Y sky130_fd_sc_hd__xor2_1_169/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_365 vssd1 vccd1 sky130_fd_sc_hd__inv_2_11/Y sky130_fd_sc_hd__nor2_1_95/Y
+ sky130_fd_sc_hd__nand2_1_282/Y sky130_fd_sc_hd__xnor2_1_49/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_376 vssd1 vccd1 sky130_fd_sc_hd__inv_2_16/Y sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__o21ai_1_376/B1 sky130_fd_sc_hd__xor2_1_190/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_387 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_3/A sky130_fd_sc_hd__nor2_2_6/Y
+ sky130_fd_sc_hd__nand2_1_311/Y sky130_fd_sc_hd__xnor2_1_58/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_398 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_313/A sky130_fd_sc_hd__nor2_1_124/Y
+ sky130_fd_sc_hd__nand2_1_389/Y sky130_fd_sc_hd__xnor2_1_86/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_808 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_819 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_703 sky130_fd_sc_hd__nand2_1_703/Y sky130_fd_sc_hd__or2_0_81/A
+ la_data_out[71] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_714 sky130_fd_sc_hd__inv_2_66/A sky130_fd_sc_hd__and2_0_1/X
+ sky130_fd_sc_hd__nor3_1_1/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_12 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_12/A1 sky130_fd_sc_hd__buf_2_148/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__or2_0_78/A vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_725 sky130_fd_sc_hd__xor2_1_652/B sky130_fd_sc_hd__nand2_1_726/Y
+ sky130_fd_sc_hd__nand2_1_725/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_23 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_23/A1 sky130_fd_sc_hd__buf_2_84/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__fa_2_416/A vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_736 sky130_fd_sc_hd__nand2_1_736/Y sky130_fd_sc_hd__or2_0_89/X
+ sky130_fd_sc_hd__or2_0_90/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_34 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_34/A1 sky130_fd_sc_hd__inv_8_2/Y
+ sky130_fd_sc_hd__mux2_8_1/S sky130_fd_sc_hd__mux2_2_34/X vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_747 sky130_fd_sc_hd__xor2_1_657/B sky130_fd_sc_hd__nand2_1_748/Y
+ sky130_fd_sc_hd__nand2_1_747/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_45 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_45/A1 sky130_fd_sc_hd__buf_2_85/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__fa_2_417/B vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_758 sky130_fd_sc_hd__xnor2_1_213/A sky130_fd_sc_hd__nand2_1_773/Y
+ sky130_fd_sc_hd__nand2_1_758/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_769 sky130_fd_sc_hd__and2_0_301/B sky130_fd_sc_hd__or2_0_85/A
+ sky130_fd_sc_hd__or2_0_85/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__conb_1_120 sky130_fd_sc_hd__conb_1_120/LO sky130_fd_sc_hd__conb_1_120/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_131 sky130_fd_sc_hd__conb_1_131/LO sky130_fd_sc_hd__conb_1_131/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_142 sky130_fd_sc_hd__conb_1_142/LO sky130_fd_sc_hd__clkinv_1_0/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_1807 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_510 la_data_out[33] sky130_fd_sc_hd__dfxtp_1_520/CLK sky130_fd_sc_hd__and2_0_351/X
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_170 sky130_fd_sc_hd__fa_2_122/A sky130_fd_sc_hd__nor2_2_8/B
+ sky130_fd_sc_hd__xor2_1_170/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1818 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_521 wbs_dat_o[0] sky130_fd_sc_hd__dfxtp_1_533/CLK sky130_fd_sc_hd__nor2b_1_157/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_181 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__fa_2_131/B
+ sky130_fd_sc_hd__xor2_1_181/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1829 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_532 wbs_dat_o[11] sky130_fd_sc_hd__dfxtp_1_532/CLK sky130_fd_sc_hd__nor2b_1_146/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_192 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__xor2_1_192/X
+ sky130_fd_sc_hd__xor2_1_192/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_543 wbs_dat_o[22] sky130_fd_sc_hd__dfxtp_1_544/CLK sky130_fd_sc_hd__nor2b_1_135/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_554 wbs_ack_o sky130_fd_sc_hd__clkinv_4_77/Y sky130_fd_sc_hd__nor2b_1_125/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_130 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_130/X sky130_fd_sc_hd__inv_2_0/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_201 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__nor2_2_5/B
+ sky130_fd_sc_hd__nor2_2_4/B sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__buf_2_4/A
+ sky130_fd_sc_hd__o21ai_1_371/B1 sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_141 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_141/X sky130_fd_sc_hd__clkinv_1_868/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_212 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__buf_2_32/X sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__o21ai_1_389/B1 sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_152 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_38/A1 sky130_fd_sc_hd__clkbuf_1_152/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_223 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__or2_0_9/B
+ sky130_fd_sc_hd__or2_0_9/A sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__or2_0_4/B
+ sky130_fd_sc_hd__o21ai_1_412/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_163 vssd1 vccd1 sky130_fd_sc_hd__buf_8_4/A sky130_fd_sc_hd__buf_8_2/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_234 vccd1 vssd1 sky130_fd_sc_hd__and3_4_15/X sky130_fd_sc_hd__buf_2_19/X
+ sky130_fd_sc_hd__buf_6_5/X sky130_fd_sc_hd__nor2_1_130/Y sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__o21ai_1_428/B1 sky130_fd_sc_hd__nor2b_1_11/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_174 vssd1 vccd1 sky130_fd_sc_hd__a22o_1_29/B2 sky130_fd_sc_hd__clkbuf_1_174/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_245 vccd1 vssd1 sky130_fd_sc_hd__and3_4_11/X sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__buf_4_5/X sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__o21ai_1_441/B1 sky130_fd_sc_hd__and2b_4_8/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_185 vssd1 vccd1 sky130_fd_sc_hd__buf_2_142/A sky130_fd_sc_hd__buf_6_93/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_256 vccd1 vssd1 sky130_fd_sc_hd__and3_4_10/X sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__nor2_1_73/B sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__o21ai_1_457/B1 sky130_fd_sc_hd__and2b_4_7/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_196 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_277/A sky130_fd_sc_hd__clkbuf_1_49/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_404 sky130_fd_sc_hd__fa_2_403/A sky130_fd_sc_hd__fa_2_405/CIN
+ sky130_fd_sc_hd__fa_2_404/A sky130_fd_sc_hd__fa_2_404/B sky130_fd_sc_hd__fa_2_404/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_267 vccd1 vssd1 sky130_fd_sc_hd__and3_4_14/X sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__buf_6_2/X sky130_fd_sc_hd__nor2_1_127/Y sky130_fd_sc_hd__buf_4_7/X
+ sky130_fd_sc_hd__o21ai_1_469/B1 sky130_fd_sc_hd__nor2b_1_10/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_415 sky130_fd_sc_hd__xor2_1_638/B sky130_fd_sc_hd__fa_2_415/SUM
+ sky130_fd_sc_hd__fa_2_415/A sky130_fd_sc_hd__fa_2_415/B sky130_fd_sc_hd__fa_2_415/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_278 vccd1 vssd1 sky130_fd_sc_hd__and3_4_10/X sky130_fd_sc_hd__and2_0_45/A
+ sky130_fd_sc_hd__and2_0_87/A sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__buf_6_0/X
+ sky130_fd_sc_hd__o21ai_1_484/B1 sky130_fd_sc_hd__and2b_4_7/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_426 sky130_fd_sc_hd__fa_2_422/B sky130_fd_sc_hd__fa_2_428/B
+ sky130_fd_sc_hd__fa_2_426/A sky130_fd_sc_hd__fa_2_426/B sky130_fd_sc_hd__o22ai_1_64/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_289 vccd1 vssd1 sky130_fd_sc_hd__and3_4_11/X sky130_fd_sc_hd__and2_0_87/A
+ sky130_fd_sc_hd__buf_6_0/X sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__o21ai_1_499/B1 sky130_fd_sc_hd__and2b_4_8/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_437 sky130_fd_sc_hd__nor2_1_247/A sky130_fd_sc_hd__or2_0_94/B
+ sky130_fd_sc_hd__fa_2_437/A sky130_fd_sc_hd__fa_2_437/B sky130_fd_sc_hd__fa_2_437/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_448 sky130_fd_sc_hd__fa_2_423/B sky130_fd_sc_hd__fa_2_448/SUM
+ sky130_fd_sc_hd__fa_2_448/A sky130_fd_sc_hd__fa_2_448/B sky130_fd_sc_hd__fa_2_448/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_459 sky130_fd_sc_hd__fa_2_447/A sky130_fd_sc_hd__fah_1_18/CI
+ sky130_fd_sc_hd__fa_2_459/A sky130_fd_sc_hd__fa_2_459/B sky130_fd_sc_hd__fa_2_459/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_4_20 sky130_fd_sc_hd__inv_4_20/Y wbs_dat_i[12] vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__and2_0_150 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_40/D sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_150/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_161 vccd1 vssd1 sky130_fd_sc_hd__and2_0_161/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_161/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_172 vccd1 vssd1 sky130_fd_sc_hd__and2_0_172/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_172/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_80 io_out[21] sky130_fd_sc_hd__conb_1_62/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_183 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_46/D sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__o21ai_1_94/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_91 io_out[10] sky130_fd_sc_hd__conb_1_51/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_194 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_81/D sky130_fd_sc_hd__o21ai_2_0/B1
+ sky130_fd_sc_hd__o21ai_1_87/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_12_409 sky130_fd_sc_hd__buf_12_409/A sky130_fd_sc_hd__buf_12_629/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__sdlclkp_1_0 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_4_1/Y
+ sky130_fd_sc_hd__dfxtp_1_43/CLK sky130_fd_sc_hd__o21ai_1_0/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__sdlclkp_1
Xsky130_fd_sc_hd__clkinv_1_609 sky130_fd_sc_hd__nand2_1_648/A sky130_fd_sc_hd__nor2_1_217/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_140 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_141/A2 sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__a22oi_1_180/Y sky130_fd_sc_hd__and2_0_128/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_151 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_153/A2 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_143/Y sky130_fd_sc_hd__and2_0_113/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_162 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_83/A sky130_fd_sc_hd__nor2_1_62/Y
+ sky130_fd_sc_hd__nand2_1_207/Y sky130_fd_sc_hd__xnor2_1_19/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_173 vssd1 vccd1 sky130_fd_sc_hd__inv_2_22/Y sky130_fd_sc_hd__nand2b_1_7/Y
+ sky130_fd_sc_hd__a222oi_1_54/Y sky130_fd_sc_hd__xor2_1_6/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_184 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_251/A2 sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__a222oi_1_63/Y sky130_fd_sc_hd__xor2_1_15/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_195 vssd1 vccd1 sky130_fd_sc_hd__inv_2_16/Y sky130_fd_sc_hd__nand2b_1_4/Y
+ sky130_fd_sc_hd__a222oi_1_71/Y sky130_fd_sc_hd__xor2_1_24/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_18 vccd1 vssd1 sky130_fd_sc_hd__nand2_1_133/A sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__xor2_1_616/X sky130_fd_sc_hd__xor2_1_191/X sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_18/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_605 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__a222oi_1_29 vccd1 vssd1 sky130_fd_sc_hd__xnor2_1_91/Y sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__xnor2_1_154/Y sky130_fd_sc_hd__xnor2_1_28/Y sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_29/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_616 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_500 sky130_fd_sc_hd__nand2_1_500/Y sky130_fd_sc_hd__nor2_4_17/Y
+ sky130_fd_sc_hd__buf_2_28/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_627 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_511 sky130_fd_sc_hd__xnor2_1_132/A sky130_fd_sc_hd__nand2_1_512/Y
+ sky130_fd_sc_hd__or2_1_9/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_638 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_522 sky130_fd_sc_hd__xnor2_1_136/A sky130_fd_sc_hd__nand2_1_523/Y
+ sky130_fd_sc_hd__or2_1_8/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_649 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_533 sky130_fd_sc_hd__xnor2_1_141/A sky130_fd_sc_hd__nand2_1_534/Y
+ sky130_fd_sc_hd__or2_1_7/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_544 sky130_fd_sc_hd__xnor2_1_145/A sky130_fd_sc_hd__nand2_1_545/Y
+ sky130_fd_sc_hd__or2_1_6/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_555 sky130_fd_sc_hd__xnor2_1_149/A sky130_fd_sc_hd__nand2_1_556/Y
+ sky130_fd_sc_hd__or2_1_5/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_566 sky130_fd_sc_hd__nand2_1_566/Y sky130_fd_sc_hd__or2_1_4/A
+ sky130_fd_sc_hd__or2_1_4/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_2 sky130_fd_sc_hd__xnor2_1_8/Y sky130_fd_sc_hd__nor2b_1_2/Y
+ sky130_fd_sc_hd__xnor2_1_5/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nand2_1_577 sky130_fd_sc_hd__xnor2_1_159/A sky130_fd_sc_hd__nand2_1_578/Y
+ sky130_fd_sc_hd__nand2_1_577/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_588 sky130_fd_sc_hd__nand2_1_588/Y sky130_fd_sc_hd__nor2_1_190/Y
+ sky130_fd_sc_hd__nand2_1_599/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_599 sky130_fd_sc_hd__nand2_1_599/Y sky130_fd_sc_hd__nand2_1_605/A
+ sky130_fd_sc_hd__nand2_1_599/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_1102 sky130_fd_sc_hd__clkinv_4_45/A sky130_fd_sc_hd__a22o_1_22/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1113 sky130_fd_sc_hd__clkinv_4_56/A sky130_fd_sc_hd__a22o_1_33/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1124 sky130_fd_sc_hd__clkinv_4_67/A sky130_fd_sc_hd__a22o_1_44/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1135 sky130_fd_sc_hd__clkinv_1_846/A wbs_dat_i[31] vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1146 sky130_fd_sc_hd__buf_2_186/A sky130_fd_sc_hd__inv_4_18/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1604 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1615 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1626 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1637 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_340 sky130_fd_sc_hd__a22oi_1_1/B2 sky130_fd_sc_hd__dfxtp_1_343/CLK
+ sky130_fd_sc_hd__and2_0_331/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1648 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_351 sky130_fd_sc_hd__dfxtp_1_351/Q sky130_fd_sc_hd__dfxtp_1_354/CLK
+ sky130_fd_sc_hd__and2_0_315/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1659 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_362 sky130_fd_sc_hd__a221o_1_0/B1 sky130_fd_sc_hd__dfxtp_1_29/CLK
+ sky130_fd_sc_hd__ha_2_3/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_373 sky130_fd_sc_hd__dfxtp_1_373/Q sky130_fd_sc_hd__dfxtp_1_375/CLK
+ sky130_fd_sc_hd__nor2b_1_110/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_384 sky130_fd_sc_hd__dfxtp_1_384/Q sky130_fd_sc_hd__dfxtp_1_392/CLK
+ sky130_fd_sc_hd__nor2b_1_99/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_4 sky130_fd_sc_hd__nand2_1_4/Y sky130_fd_sc_hd__nand2_1_7/B
+ sky130_fd_sc_hd__or2_0_82/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_395 sky130_fd_sc_hd__dfxtp_1_395/Q sky130_fd_sc_hd__dfxtp_1_395/CLK
+ sky130_fd_sc_hd__nor2b_1_89/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_201 sky130_fd_sc_hd__nor2_2_13/A sky130_fd_sc_hd__or2_0_30/B
+ sky130_fd_sc_hd__fa_2_201/A sky130_fd_sc_hd__fa_2_201/B sky130_fd_sc_hd__fa_2_201/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_212 sky130_fd_sc_hd__fa_2_208/B sky130_fd_sc_hd__fa_2_215/CIN
+ sky130_fd_sc_hd__fa_2_212/A sky130_fd_sc_hd__fa_2_212/B sky130_fd_sc_hd__fa_2_212/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_223 sky130_fd_sc_hd__fa_2_219/CIN sky130_fd_sc_hd__fa_2_228/A
+ sky130_fd_sc_hd__fa_2_223/A sky130_fd_sc_hd__fa_2_223/B sky130_fd_sc_hd__fa_2_227/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_234 sky130_fd_sc_hd__or2_0_34/A sky130_fd_sc_hd__nor2_2_15/B
+ sky130_fd_sc_hd__fa_2_234/A sky130_fd_sc_hd__fa_2_234/B sky130_fd_sc_hd__fa_2_234/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_245 sky130_fd_sc_hd__or2_0_35/A sky130_fd_sc_hd__nor2_2_14/B
+ sky130_fd_sc_hd__fa_2_245/A sky130_fd_sc_hd__fa_2_245/B sky130_fd_sc_hd__fa_2_245/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_256 sky130_fd_sc_hd__fa_2_254/CIN sky130_fd_sc_hd__fa_2_259/A
+ sky130_fd_sc_hd__fa_2_256/A sky130_fd_sc_hd__fa_2_256/B sky130_fd_sc_hd__xor2_1_375/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_267 sky130_fd_sc_hd__fa_2_265/B sky130_fd_sc_hd__fa_2_268/A
+ sky130_fd_sc_hd__fa_2_267/A sky130_fd_sc_hd__fa_2_267/B sky130_fd_sc_hd__fa_2_267/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_278 sky130_fd_sc_hd__nor2_1_155/A sky130_fd_sc_hd__or2_0_43/B
+ sky130_fd_sc_hd__fa_2_278/A sky130_fd_sc_hd__fa_2_278/B sky130_fd_sc_hd__fa_2_278/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_289 sky130_fd_sc_hd__xor3_1_27/B sky130_fd_sc_hd__fa_2_290/CIN
+ sky130_fd_sc_hd__fa_2_289/A sky130_fd_sc_hd__fa_2_289/B sky130_fd_sc_hd__xor2_1_437/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_5 vccd1 vssd1 sky130_fd_sc_hd__and2_0_5/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_5/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__fa_2_70 sky130_fd_sc_hd__fa_2_66/B sky130_fd_sc_hd__fa_2_73/CIN
+ sky130_fd_sc_hd__fa_2_70/A sky130_fd_sc_hd__fa_2_70/B sky130_fd_sc_hd__fa_2_70/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_81 sky130_fd_sc_hd__fa_2_77/CIN sky130_fd_sc_hd__fa_2_86/A
+ sky130_fd_sc_hd__fa_2_81/A sky130_fd_sc_hd__fa_2_81/B sky130_fd_sc_hd__fa_2_85/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_92 sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__nor2_1_69/B
+ sky130_fd_sc_hd__fa_2_92/A sky130_fd_sc_hd__fa_2_92/B sky130_fd_sc_hd__fa_2_92/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a21oi_1_20 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_49/Y
+ sky130_fd_sc_hd__a21oi_1_20/Y sky130_fd_sc_hd__dfxtp_1_77/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_31 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_60/Y
+ sky130_fd_sc_hd__a21oi_1_31/Y sky130_fd_sc_hd__dfxtp_1_66/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_42 sky130_fd_sc_hd__a21oi_1_45/A1 sky130_fd_sc_hd__o21ai_1_221/Y
+ sky130_fd_sc_hd__a21oi_1_42/Y sky130_fd_sc_hd__nor2_1_54/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_206 sky130_fd_sc_hd__buf_6_58/X sky130_fd_sc_hd__buf_12_296/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_53 sky130_fd_sc_hd__xnor2_1_41/B sky130_fd_sc_hd__o21ai_1_335/Y
+ sky130_fd_sc_hd__xor2_1_146/A sky130_fd_sc_hd__nor2_1_79/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_217 sky130_fd_sc_hd__buf_6_67/X sky130_fd_sc_hd__buf_12_357/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_64 sky130_fd_sc_hd__or2_0_23/X sky130_fd_sc_hd__a21oi_1_64/B1
+ sky130_fd_sc_hd__a21oi_1_64/Y sky130_fd_sc_hd__a21oi_1_66/B1 vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_228 sky130_fd_sc_hd__buf_6_85/X sky130_fd_sc_hd__buf_12_411/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_75 sky130_fd_sc_hd__a21oi_1_80/A1 sky130_fd_sc_hd__o21ai_1_436/Y
+ sky130_fd_sc_hd__a21oi_1_75/Y sky130_fd_sc_hd__nor2_1_112/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_239 sky130_fd_sc_hd__buf_6_55/X sky130_fd_sc_hd__buf_12_428/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_86 sky130_fd_sc_hd__a21oi_1_89/A1 sky130_fd_sc_hd__o21ai_1_562/Y
+ sky130_fd_sc_hd__a21oi_1_86/Y sky130_fd_sc_hd__nor2_1_134/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_97 sky130_fd_sc_hd__xnor2_1_119/B sky130_fd_sc_hd__nand2_1_464/Y
+ sky130_fd_sc_hd__xnor2_1_63/A sky130_fd_sc_hd__nor2_1_156/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_1_109 sky130_fd_sc_hd__inv_2_54/Y sky130_fd_sc_hd__inv_4_7/Y
+ sky130_fd_sc_hd__dfxtp_1_177/Q sky130_fd_sc_hd__dfxtp_1_145/Q sky130_fd_sc_hd__o21ai_1_15/B1
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor3_1_1 sky130_fd_sc_hd__or4_1_1/X sky130_fd_sc_hd__nor3_1_1/Y
+ sky130_fd_sc_hd__ha_2_8/A sky130_fd_sc_hd__ha_2_6/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__clkinv_1_406 sky130_fd_sc_hd__and3_4_0/A sky130_fd_sc_hd__xor2_1_212/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_417 sky130_fd_sc_hd__o21ai_1_421/A2 sky130_fd_sc_hd__xnor2_1_70/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_428 sky130_fd_sc_hd__nor2_1_113/B sky130_fd_sc_hd__nor2_1_115/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_439 sky130_fd_sc_hd__nor2_1_119/B sky130_fd_sc_hd__nand2_1_376/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_60 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_71 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_82 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_93 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_60 vccd1 vssd1 sky130_fd_sc_hd__buf_6_60/X sky130_fd_sc_hd__buf_8_75/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_71 vccd1 vssd1 sky130_fd_sc_hd__buf_6_71/X sky130_fd_sc_hd__buf_8_13/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_82 vccd1 vssd1 sky130_fd_sc_hd__buf_6_82/X sky130_fd_sc_hd__buf_6_82/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_93 vccd1 vssd1 sky130_fd_sc_hd__buf_6_93/X wbs_dat_i[5] vssd1
+ vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_40 sky130_fd_sc_hd__buf_2_193/A vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_51 sky130_fd_sc_hd__buf_2_189/A vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_62 sky130_fd_sc_hd__dfxtp_1_12/Q vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a222oi_1_6 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_347/Q sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__o211ai_1_22/Y sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__a222oi_1_6/Y sky130_fd_sc_hd__dfxtp_1_298/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_402 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_413 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_424 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_435 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_446 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_330 sky130_fd_sc_hd__nand2_1_330/Y sky130_fd_sc_hd__nor2_4_13/Y
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_457 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_341 sky130_fd_sc_hd__nor2_1_108/A sky130_fd_sc_hd__or2_0_38/X
+ sky130_fd_sc_hd__nand2_1_341/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_468 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_940 sky130_fd_sc_hd__clkinv_1_941/A sky130_fd_sc_hd__buf_8_79/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_352 sky130_fd_sc_hd__nand2_1_352/Y sky130_fd_sc_hd__nor2_1_113/Y
+ sky130_fd_sc_hd__nand2_1_374/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_479 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_951 sky130_fd_sc_hd__clkbuf_1_52/A sky130_fd_sc_hd__clkinv_4_20/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_363 sky130_fd_sc_hd__nand2_1_363/Y sky130_fd_sc_hd__nor2_1_118/Y
+ sky130_fd_sc_hd__nand2_1_374/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_962 sky130_fd_sc_hd__inv_8_1/A sky130_fd_sc_hd__clkinv_1_962/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_374 sky130_fd_sc_hd__nand2_1_374/Y sky130_fd_sc_hd__or2_0_41/X
+ sky130_fd_sc_hd__nand2_1_374/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_973 sky130_fd_sc_hd__clkinv_1_973/Y sky130_fd_sc_hd__clkinv_4_23/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_385 sky130_fd_sc_hd__nand2_1_385/Y sky130_fd_sc_hd__or2_0_47/X
+ sky130_fd_sc_hd__nor2_1_126/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_984 sky130_fd_sc_hd__clkinv_1_984/Y sky130_fd_sc_hd__clkinv_4_28/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_396 sky130_fd_sc_hd__xnor2_1_92/A sky130_fd_sc_hd__nand2_1_397/Y
+ sky130_fd_sc_hd__or2_0_45/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_995 sky130_fd_sc_hd__clkinv_1_996/A sky130_fd_sc_hd__inv_4_6/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1401 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1412 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1423 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1434 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1445 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1456 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1467 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_170 sky130_fd_sc_hd__dfxtp_1_170/Q sky130_fd_sc_hd__dfxtp_1_170/CLK
+ sky130_fd_sc_hd__and2_0_157/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1478 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_181 sky130_fd_sc_hd__dfxtp_1_181/Q sky130_fd_sc_hd__clkinv_4_2/Y
+ sky130_fd_sc_hd__and2_0_213/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_909 vssd1 vccd1 sky130_fd_sc_hd__nor2_2_1/B sky130_fd_sc_hd__a31oi_1_0/Y
+ sky130_fd_sc_hd__a31oi_1_2/Y sky130_fd_sc_hd__o21ai_1_909/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1489 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_192 sky130_fd_sc_hd__xor2_1_637/A sky130_fd_sc_hd__dfxtp_4_3/CLK
+ sky130_fd_sc_hd__and2_0_33/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_2_18 vccd1 vssd1 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__buf_2_18/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_29 vccd1 vssd1 sky130_fd_sc_hd__buf_2_29/X sky130_fd_sc_hd__buf_8_0/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_980 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_991 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o211ai_1_12 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_51/B1
+ sky130_fd_sc_hd__a22oi_1_6/A2 sky130_fd_sc_hd__a22oi_1_56/Y sky130_fd_sc_hd__a22oi_1_57/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_23 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_40/B1
+ sky130_fd_sc_hd__o211ai_1_23/Y sky130_fd_sc_hd__a22oi_1_78/Y sky130_fd_sc_hd__a22oi_1_79/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_34 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o21ai_1_4/A2
+ sky130_fd_sc_hd__fa_2_310/B sky130_fd_sc_hd__nand2_1_54/Y sky130_fd_sc_hd__a21oi_1_5/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_45 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o22ai_1_18/B1
+ sky130_fd_sc_hd__fa_2_379/B sky130_fd_sc_hd__nand2_1_65/Y sky130_fd_sc_hd__a21oi_1_16/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_56 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o22ai_1_7/B1
+ sky130_fd_sc_hd__fa_2_408/A sky130_fd_sc_hd__nand2_1_76/Y sky130_fd_sc_hd__a21oi_1_27/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__clkinv_1_203 sky130_fd_sc_hd__nor2_1_18/A sky130_fd_sc_hd__dfxtp_1_141/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_214 sky130_fd_sc_hd__o22ai_1_53/B1 sky130_fd_sc_hd__dfxtp_1_169/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_225 sky130_fd_sc_hd__o22ai_1_7/B1 sky130_fd_sc_hd__dfxtp_1_102/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_236 sky130_fd_sc_hd__nor2_1_7/A sky130_fd_sc_hd__dfxtp_1_130/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_247 sky130_fd_sc_hd__o21ai_1_57/A2 sky130_fd_sc_hd__xnor2_1_141/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_258 sky130_fd_sc_hd__o21ai_1_121/A2 sky130_fd_sc_hd__xor2_1_602/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_269 sky130_fd_sc_hd__nor2_1_37/A sky130_fd_sc_hd__nor2_1_40/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_2_3 sky130_fd_sc_hd__buf_2_16/A sky130_fd_sc_hd__o21ai_2_3/Y
+ sky130_fd_sc_hd__o21ai_2_3/A2 sky130_fd_sc_hd__o21ai_2_4/A2 vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__o21ai_2
Xsky130_fd_sc_hd__xor3_1_9 sky130_fd_sc_hd__xor3_1_9/X sky130_fd_sc_hd__xor3_1_9/C
+ sky130_fd_sc_hd__xor3_1_9/B sky130_fd_sc_hd__xor3_1_9/A vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__xor3_1
Xsky130_fd_sc_hd__and3_4_16 sky130_fd_sc_hd__nor2_2_19/B sky130_fd_sc_hd__nor2b_2_3/A
+ sky130_fd_sc_hd__nor2_2_19/A sky130_fd_sc_hd__and3_4_16/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__a21oi_1_100 sky130_fd_sc_hd__nand2_1_483/Y sky130_fd_sc_hd__nand2_1_472/Y
+ sky130_fd_sc_hd__a21oi_1_100/Y sky130_fd_sc_hd__nor2_1_158/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_111 sky130_fd_sc_hd__clkinv_1_549/Y sky130_fd_sc_hd__o21ai_1_681/Y
+ sky130_fd_sc_hd__a21oi_1_111/Y sky130_fd_sc_hd__nor2_1_170/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_122 sky130_fd_sc_hd__clkinv_1_580/Y sky130_fd_sc_hd__nand2_1_593/Y
+ sky130_fd_sc_hd__a21oi_1_122/Y sky130_fd_sc_hd__nor2_1_192/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_133 sky130_fd_sc_hd__xnor2_1_181/B sky130_fd_sc_hd__clkinv_1_602/Y
+ sky130_fd_sc_hd__xnor2_1_128/A sky130_fd_sc_hd__nand2_1_644/A vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_144 sky130_fd_sc_hd__xnor2_1_194/B sky130_fd_sc_hd__clkinv_1_637/Y
+ sky130_fd_sc_hd__xor2_1_645/A sky130_fd_sc_hd__or2_0_78/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_155 sky130_fd_sc_hd__xnor2_1_208/B sky130_fd_sc_hd__clkinv_1_669/Y
+ sky130_fd_sc_hd__xor2_1_655/A sky130_fd_sc_hd__or2_0_89/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_166 sky130_fd_sc_hd__nor2_1_250/Y sky130_fd_sc_hd__o21ai_1_888/Y
+ sky130_fd_sc_hd__a21oi_1_166/Y sky130_fd_sc_hd__o21ai_1_889/Y vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_177 sky130_fd_sc_hd__xnor2_1_298/B sky130_fd_sc_hd__clkinv_1_822/Y
+ sky130_fd_sc_hd__xor2_1_683/A sky130_fd_sc_hd__or2_0_107/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_188 sky130_fd_sc_hd__nand2_1_854/Y sky130_fd_sc_hd__nor2_1_273/A
+ sky130_fd_sc_hd__nor2_1_273/B sky130_fd_sc_hd__nor2b_1_121/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_199 la_data_out[52] sky130_fd_sc_hd__xor2_1_696/X sky130_fd_sc_hd__a21oi_1_199/Y
+ sky130_fd_sc_hd__nand2_1_861/B vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_107 sky130_fd_sc_hd__buf_8_107/A sky130_fd_sc_hd__buf_8_107/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_118 sky130_fd_sc_hd__buf_8_118/A sky130_fd_sc_hd__buf_6_50/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_129 sky130_fd_sc_hd__buf_8_129/A sky130_fd_sc_hd__buf_8_129/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_12_570 sky130_fd_sc_hd__buf_12_570/A sky130_fd_sc_hd__buf_12_570/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_581 sky130_fd_sc_hd__buf_12_581/A sky130_fd_sc_hd__buf_12_581/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_210 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_592 sky130_fd_sc_hd__buf_12_592/A sky130_fd_sc_hd__buf_12_592/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_221 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_232 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_243 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_254 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_265 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_300 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_300/B sky130_fd_sc_hd__xnor2_1_300/Y
+ sky130_fd_sc_hd__xnor2_1_300/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__decap_12_276 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_311 vssd1 vccd1 sky130_fd_sc_hd__ha_2_59/SUM sky130_fd_sc_hd__xnor2_1_311/Y
+ la_data_out[55] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_160 sky130_fd_sc_hd__nand2_1_160/Y sky130_fd_sc_hd__nor2_4_9/Y
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_287 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_171 sky130_fd_sc_hd__xnor2_1_7/A sky130_fd_sc_hd__nand2_1_172/Y
+ sky130_fd_sc_hd__or2_0_9/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_298 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_770 sky130_fd_sc_hd__or2_0_112/A sky130_fd_sc_hd__clkinv_1_770/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_182 sky130_fd_sc_hd__xnor2_1_11/A sky130_fd_sc_hd__nand2_1_183/Y
+ sky130_fd_sc_hd__or2_0_12/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_781 sky130_fd_sc_hd__and2_0_326/A sky130_fd_sc_hd__clkinv_1_781/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_193 sky130_fd_sc_hd__xnor2_1_16/A sky130_fd_sc_hd__nand2_1_194/Y
+ sky130_fd_sc_hd__or2_0_15/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_792 sky130_fd_sc_hd__and2_0_315/A sky130_fd_sc_hd__clkinv_1_792/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1220 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1231 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1242 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1253 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1264 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1275 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_706 vssd1 vccd1 sky130_fd_sc_hd__inv_2_48/Y sky130_fd_sc_hd__nand2b_1_20/Y
+ sky130_fd_sc_hd__o21ai_1_706/B1 sky130_fd_sc_hd__xor2_1_485/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1286 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_717 vssd1 vccd1 sky130_fd_sc_hd__inv_2_46/Y sky130_fd_sc_hd__nand2b_1_20/Y
+ sky130_fd_sc_hd__o21ai_1_717/B1 sky130_fd_sc_hd__xor2_1_494/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1297 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_728 vssd1 vccd1 sky130_fd_sc_hd__inv_2_45/Y sky130_fd_sc_hd__nand2b_1_16/Y
+ sky130_fd_sc_hd__o21ai_1_728/B1 sky130_fd_sc_hd__xor2_1_505/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_739 vssd1 vccd1 sky130_fd_sc_hd__inv_2_43/Y sky130_fd_sc_hd__nand2b_1_16/Y
+ sky130_fd_sc_hd__o21ai_1_739/B1 sky130_fd_sc_hd__xor2_1_515/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_13 sky130_fd_sc_hd__fa_2_75/A sky130_fd_sc_hd__fa_2_7/A sky130_fd_sc_hd__xor2_1_13/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__and3_1_0 vssd1 vccd1 sky130_fd_sc_hd__and3_1_0/X sky130_fd_sc_hd__and3_1_0/B
+ sky130_fd_sc_hd__and3_1_0/A sky130_fd_sc_hd__and3_1_0/C vssd1 vccd1 sky130_fd_sc_hd__and3_1
Xsky130_fd_sc_hd__xor2_1_24 sky130_fd_sc_hd__fa_2_56/A sky130_fd_sc_hd__fa_2_9/A sky130_fd_sc_hd__xor2_1_24/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_35 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__xor2_1_35/X
+ sky130_fd_sc_hd__xor2_1_35/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_46 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__xor2_1_46/X
+ sky130_fd_sc_hd__xor2_1_46/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_57 sky130_fd_sc_hd__xor2_1_6/B sky130_fd_sc_hd__xor2_1_57/X
+ sky130_fd_sc_hd__xor2_1_57/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_68 sky130_fd_sc_hd__fa_2_75/A sky130_fd_sc_hd__fa_2_49/B
+ sky130_fd_sc_hd__xor2_1_68/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_79 sky130_fd_sc_hd__xor2_1_9/B sky130_fd_sc_hd__fa_2_57/A
+ sky130_fd_sc_hd__xor2_1_79/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2b_1_7 sky130_fd_sc_hd__nand2b_1_7/Y sky130_fd_sc_hd__nor2_2_7/A
+ sky130_fd_sc_hd__nor2_2_7/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__xor2_1_500 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__fa_2_336/A
+ sky130_fd_sc_hd__xor2_1_500/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_511 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__fa_2_344/B
+ sky130_fd_sc_hd__xor2_1_511/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a21o_2_3 sky130_fd_sc_hd__a21o_2_3/X sky130_fd_sc_hd__a21o_2_3/B1
+ wbs_adr_i[7] sky130_fd_sc_hd__a21o_2_3/A2 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__xor2_1_522 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__fa_2_350/A
+ sky130_fd_sc_hd__xor2_1_522/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_533 sky130_fd_sc_hd__xor2_1_548/B sky130_fd_sc_hd__fa_2_361/B
+ sky130_fd_sc_hd__xor2_1_533/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_544 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__xor2_1_544/X
+ sky130_fd_sc_hd__xor2_1_544/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_555 sky130_fd_sc_hd__fa_2_389/A sky130_fd_sc_hd__fa_2_376/B
+ sky130_fd_sc_hd__xor2_1_555/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_566 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__xor2_1_566/X
+ sky130_fd_sc_hd__xor2_1_566/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_577 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__xor2_1_577/X
+ sky130_fd_sc_hd__xor2_1_577/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_588 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__xor2_1_588/X
+ sky130_fd_sc_hd__xor2_1_588/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_599 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__xor2_1_599/X
+ sky130_fd_sc_hd__xor2_1_599/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a222oi_1_608 vccd1 vssd1 sky130_fd_sc_hd__nor2_1_273/Y sky130_fd_sc_hd__o31ai_1_1/A1
+ sky130_fd_sc_hd__a21o_2_0/X sky130_fd_sc_hd__nand3_1_5/B sky130_fd_sc_hd__nand2_1_853/Y
+ sky130_fd_sc_hd__o21ai_1_913/A1 sky130_fd_sc_hd__nor2_1_271/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__ha_2_40 vssd1 vccd1 sky130_fd_sc_hd__or4_1_3/C sky130_fd_sc_hd__xor2_1_692/A
+ sky130_fd_sc_hd__ha_2_40/SUM sky130_fd_sc_hd__ha_2_40/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__and2b_4_2 sky130_fd_sc_hd__and3_4_3/B sky130_fd_sc_hd__and2b_4_2/X
+ sky130_fd_sc_hd__and3_4_3/C vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__and2b_4
Xsky130_fd_sc_hd__ha_2_51 vssd1 vccd1 sky130_fd_sc_hd__ha_2_51/A sky130_fd_sc_hd__ha_2_53/B
+ sky130_fd_sc_hd__ha_2_51/SUM sky130_fd_sc_hd__ha_2_51/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_3 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_3/X sky130_fd_sc_hd__or2_0_52/B
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkinv_1_3 la_data_out[124] sky130_fd_sc_hd__clkinv_1_3/A vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_160 sky130_fd_sc_hd__buf_8_0/X sky130_fd_sc_hd__nor2_1_160/Y
+ sky130_fd_sc_hd__buf_6_2/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_171 sky130_fd_sc_hd__nor2_1_171/B sky130_fd_sc_hd__nor2_1_171/Y
+ sky130_fd_sc_hd__nor2_1_171/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_182 sky130_fd_sc_hd__nor2_1_182/B sky130_fd_sc_hd__nor2_1_182/Y
+ sky130_fd_sc_hd__nor2_1_182/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_193 sky130_fd_sc_hd__nor2_2_10/B sky130_fd_sc_hd__nor2_1_193/Y
+ sky130_fd_sc_hd__buf_6_4/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_80 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__nor2_4_3/Y
+ sky130_fd_sc_hd__nand2_1_58/B sky130_fd_sc_hd__dfxtp_1_151/Q sky130_fd_sc_hd__a22oi_1_80/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_91 sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__dfxtp_1_124/Q sky130_fd_sc_hd__dfxtp_1_92/Q sky130_fd_sc_hd__a22oi_1_91/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__and2_0_18 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_4_3/D sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__buf_2_14/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_29 vccd1 vssd1 sky130_fd_sc_hd__and2_0_29/X sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__buf_8_0/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_8_17 sky130_fd_sc_hd__inv_2_76/Y sky130_fd_sc_hd__buf_8_17/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xnor2_1_130 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_134/A sky130_fd_sc_hd__nor2b_1_13/A
+ sky130_fd_sc_hd__nor2_1_167/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__buf_8_28 sky130_fd_sc_hd__inv_2_70/Y sky130_fd_sc_hd__buf_8_28/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xnor2_1_141 vssd1 vccd1 sky130_fd_sc_hd__o21ai_2_13/Y sky130_fd_sc_hd__xnor2_1_141/Y
+ sky130_fd_sc_hd__xnor2_1_141/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__buf_8_39 sky130_fd_sc_hd__inv_2_92/Y sky130_fd_sc_hd__buf_8_39/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xnor2_1_152 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_152/B sky130_fd_sc_hd__xnor2_1_152/Y
+ sky130_fd_sc_hd__xnor2_1_152/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_163 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_163/B sky130_fd_sc_hd__inv_2_50/A
+ sky130_fd_sc_hd__xnor2_1_163/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_174 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_174/B sky130_fd_sc_hd__inv_2_44/A
+ sky130_fd_sc_hd__xnor2_1_174/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_185 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_185/B sky130_fd_sc_hd__xnor2_1_185/Y
+ sky130_fd_sc_hd__xnor2_1_185/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_196 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_196/B sky130_fd_sc_hd__and2_0_261/A
+ sky130_fd_sc_hd__xnor2_1_196/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_4_80 wbs_dat_i[26] sky130_fd_sc_hd__inv_2_94/A vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_91 wbs_dat_i[3] sky130_fd_sc_hd__inv_2_107/A vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_1050 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1061 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1072 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_503 vssd1 vccd1 sky130_fd_sc_hd__buf_2_7/X sky130_fd_sc_hd__nand2b_1_13/Y
+ sky130_fd_sc_hd__o21ai_1_503/B1 sky130_fd_sc_hd__xor2_1_303/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1083 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_514 vssd1 vccd1 sky130_fd_sc_hd__inv_2_41/Y sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_514/B1 sky130_fd_sc_hd__xor2_1_314/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1094 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_525 vssd1 vccd1 sky130_fd_sc_hd__inv_2_34/Y sky130_fd_sc_hd__nand2b_1_9/Y
+ sky130_fd_sc_hd__o21ai_1_525/B1 sky130_fd_sc_hd__xor2_1_324/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_536 vssd1 vccd1 sky130_fd_sc_hd__buf_2_8/X sky130_fd_sc_hd__nand2b_1_9/Y
+ sky130_fd_sc_hd__o21ai_1_536/B1 sky130_fd_sc_hd__xor2_1_334/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_547 vssd1 vccd1 sky130_fd_sc_hd__inv_2_35/Y sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_547/B1 sky130_fd_sc_hd__xor2_1_345/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_558 vssd1 vccd1 sky130_fd_sc_hd__inv_2_33/Y sky130_fd_sc_hd__nand2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_558/B1 sky130_fd_sc_hd__xor2_1_356/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_569 vssd1 vccd1 sky130_fd_sc_hd__buf_2_9/X sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_569/B1 sky130_fd_sc_hd__xor2_1_366/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_330 sky130_fd_sc_hd__xor2_1_330/B sky130_fd_sc_hd__xor2_1_330/X
+ sky130_fd_sc_hd__xor2_1_330/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_341 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__xor2_1_341/X
+ sky130_fd_sc_hd__xor2_1_341/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_352 sky130_fd_sc_hd__fa_2_262/A sky130_fd_sc_hd__fa_2_242/A
+ sky130_fd_sc_hd__xor2_1_352/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_363 sky130_fd_sc_hd__dfxtp_2_5/Q sky130_fd_sc_hd__fa_2_251/A
+ sky130_fd_sc_hd__xor2_1_363/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_374 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__fa_2_257/B
+ sky130_fd_sc_hd__xor2_1_374/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_385 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__xor2_1_385/X
+ sky130_fd_sc_hd__xor2_1_385/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_396 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__nor2_4_12/B
+ sky130_fd_sc_hd__xor2_1_396/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_301 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_302/A sky130_fd_sc_hd__buf_8_18/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_312 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_312/X sky130_fd_sc_hd__clkinv_1_877/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_323 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_323/X sky130_fd_sc_hd__clkinv_1_873/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_334 vssd1 vccd1 la_data_out[38] sky130_fd_sc_hd__nor2b_2_0/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_405 vccd1 vssd1 sky130_fd_sc_hd__and3_4_19/X sky130_fd_sc_hd__or2_0_58/B
+ sky130_fd_sc_hd__or2_0_58/A sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__or2_0_9/B
+ sky130_fd_sc_hd__o21ai_1_671/B1 sky130_fd_sc_hd__and2b_4_9/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_345 vssd1 vccd1 sky130_fd_sc_hd__inv_4_5/A sky130_fd_sc_hd__a222oi_1_11/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_416 vccd1 vssd1 sky130_fd_sc_hd__and3_4_26/X sky130_fd_sc_hd__buf_2_21/X
+ sky130_fd_sc_hd__nor2_1_87/A sky130_fd_sc_hd__nor2_2_31/Y sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__o21ai_1_687/B1 sky130_fd_sc_hd__nor2b_1_12/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_356 vssd1 vccd1 sky130_fd_sc_hd__clkinv_2_0/A sky130_fd_sc_hd__a222oi_1_0/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_427 vccd1 vssd1 sky130_fd_sc_hd__and3_4_20/X sky130_fd_sc_hd__buf_6_4/X
+ sky130_fd_sc_hd__buf_6_0/X sky130_fd_sc_hd__nor2_4_16/Y sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__o21ai_1_701/B1 sky130_fd_sc_hd__and2b_4_11/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_438 vccd1 vssd1 sky130_fd_sc_hd__and3_4_21/X sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__buf_4_3/X sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__o21ai_1_715/B1 sky130_fd_sc_hd__and2b_4_12/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_449 vccd1 vssd1 sky130_fd_sc_hd__and3_4_20/X sky130_fd_sc_hd__nor2_1_85/B
+ sky130_fd_sc_hd__nor2_2_10/B sky130_fd_sc_hd__nor2_4_16/Y sky130_fd_sc_hd__buf_6_4/X
+ sky130_fd_sc_hd__o21ai_1_729/B1 sky130_fd_sc_hd__and2b_4_11/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__dfxtp_1_60 sky130_fd_sc_hd__nand2_1_52/B sky130_fd_sc_hd__dfxtp_1_62/CLK
+ sky130_fd_sc_hd__and2_0_6/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_71 sky130_fd_sc_hd__dfxtp_1_71/Q sky130_fd_sc_hd__dfxtp_1_72/CLK
+ sky130_fd_sc_hd__dfxtp_1_71/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_82 sky130_fd_sc_hd__dfxtp_1_82/Q sky130_fd_sc_hd__dfxtp_1_85/CLK
+ sky130_fd_sc_hd__dfxtp_1_82/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_93 sky130_fd_sc_hd__dfxtp_1_93/Q sky130_fd_sc_hd__dfxtp_1_94/CLK
+ sky130_fd_sc_hd__and2_0_14/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_310 vccd1 vssd1 sky130_fd_sc_hd__and2_0_310/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_310/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_321 vccd1 vssd1 sky130_fd_sc_hd__and2_0_321/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_321/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_332 vccd1 vssd1 sky130_fd_sc_hd__and2_0_332/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_332/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_343 vccd1 vssd1 sky130_fd_sc_hd__and2_0_343/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__clkbuf_4_9/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_354 vccd1 vssd1 sky130_fd_sc_hd__and2_0_354/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__and2_0_354/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_365 vccd1 vssd1 sky130_fd_sc_hd__and2_0_365/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_56/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_376 vccd1 vssd1 sky130_fd_sc_hd__and2_0_376/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_57/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_387 vccd1 vssd1 sky130_fd_sc_hd__and2_0_387/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_74/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_398 vccd1 vssd1 sky130_fd_sc_hd__and2_0_398/X sky130_fd_sc_hd__and2_0_401/B
+ sky130_fd_sc_hd__and2_0_398/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__conb_1_7 sky130_fd_sc_hd__conb_1_7/LO sky130_fd_sc_hd__conb_1_7/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__inv_2_110 sky130_fd_sc_hd__inv_4_10/Y sky130_fd_sc_hd__inv_2_113/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__or2_0_1 sky130_fd_sc_hd__or2_0_1/A sky130_fd_sc_hd__or2_0_1/X sky130_fd_sc_hd__or2_0_1/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__inv_2_121 sky130_fd_sc_hd__inv_2_121/A sky130_fd_sc_hd__inv_2_121/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_132 sky130_fd_sc_hd__inv_2_132/A sky130_fd_sc_hd__inv_2_132/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_143 sky130_fd_sc_hd__inv_2_143/A sky130_fd_sc_hd__buf_12_4/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_154 sky130_fd_sc_hd__inv_2_155/A sky130_fd_sc_hd__inv_2_154/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_165 sky130_fd_sc_hd__inv_2_166/A sky130_fd_sc_hd__inv_2_165/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_176 sky130_fd_sc_hd__inv_2_176/A sky130_fd_sc_hd__inv_2_177/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_187 sky130_fd_sc_hd__inv_2_187/A sky130_fd_sc_hd__inv_2_187/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_198 sky130_fd_sc_hd__inv_2_95/A sky130_fd_sc_hd__inv_2_198/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__o22ai_1_106 sky130_fd_sc_hd__nor2b_1_20/A sky130_fd_sc_hd__xnor2_1_255/Y
+ sky130_fd_sc_hd__fa_2_427/CIN sky130_fd_sc_hd__xnor2_1_267/Y sky130_fd_sc_hd__o22ai_1_78/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_117 sky130_fd_sc_hd__xnor2_2_6/Y sky130_fd_sc_hd__xnor2_1_263/Y
+ sky130_fd_sc_hd__fa_2_449/B sky130_fd_sc_hd__xnor2_1_269/Y sky130_fd_sc_hd__o22ai_1_98/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_128 sky130_fd_sc_hd__xnor2_2_5/Y sky130_fd_sc_hd__xnor2_1_276/Y
+ sky130_fd_sc_hd__fa_2_458/B sky130_fd_sc_hd__xnor2_1_281/Y sky130_fd_sc_hd__o22ai_1_95/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_139 sky130_fd_sc_hd__nand2_1_849/Y sky130_fd_sc_hd__a31o_1_0/X
+ sky130_fd_sc_hd__and2_0_399/A sky130_fd_sc_hd__nor2_1_277/B sky130_fd_sc_hd__o31ai_1_1/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_2_17 sky130_fd_sc_hd__buf_2_23/X sky130_fd_sc_hd__nor2_2_17/Y
+ sky130_fd_sc_hd__buf_4_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__nor2_2_28 sky130_fd_sc_hd__nor2_2_29/Y sky130_fd_sc_hd__nor2_2_28/Y
+ sky130_fd_sc_hd__nor2_2_28/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__o211ai_1_7 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_7/A2
+ sky130_fd_sc_hd__o211ai_1_7/Y sky130_fd_sc_hd__a22oi_1_46/Y sky130_fd_sc_hd__a22oi_1_47/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__a211o_1_0 vssd1 vccd1 sky130_fd_sc_hd__or2_0_51/B sky130_fd_sc_hd__dfxtp_1_63/Q
+ sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_0/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__o21ai_1_300 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_2/X sky130_fd_sc_hd__nor2_1_67/B
+ sky130_fd_sc_hd__o21ai_1_300/B1 sky130_fd_sc_hd__xnor2_1_30/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_311 vssd1 vccd1 sky130_fd_sc_hd__inv_2_26/Y sky130_fd_sc_hd__nand2b_1_6/Y
+ sky130_fd_sc_hd__nand2_1_156/Y sky130_fd_sc_hd__xor2_1_130/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_322 vssd1 vccd1 sky130_fd_sc_hd__nand2_4_4/Y sky130_fd_sc_hd__nand2b_1_7/Y
+ sky130_fd_sc_hd__a22oi_1_196/Y sky130_fd_sc_hd__xor2_1_142/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_333 vssd1 vccd1 sky130_fd_sc_hd__buf_2_1/X sky130_fd_sc_hd__nand2b_2_0/Y
+ sky130_fd_sc_hd__o21ai_1_333/B1 sky130_fd_sc_hd__xor2_1_152/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_344 vssd1 vccd1 sky130_fd_sc_hd__inv_2_11/Y sky130_fd_sc_hd__nor2_1_74/B
+ sky130_fd_sc_hd__a21oi_1_57/Y sky130_fd_sc_hd__xnor2_1_42/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_355 vssd1 vccd1 sky130_fd_sc_hd__inv_2_9/Y sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__o21ai_1_355/B1 sky130_fd_sc_hd__xor2_1_172/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_366 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_94/Y sky130_fd_sc_hd__nand2_1_286/Y
+ sky130_fd_sc_hd__nand2_1_280/Y sky130_fd_sc_hd__o21ai_1_366/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_377 vssd1 vccd1 sky130_fd_sc_hd__buf_2_5/X sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__o21ai_1_377/B1 sky130_fd_sc_hd__xor2_1_192/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_388 vssd1 vccd1 sky130_fd_sc_hd__nand2_4_4/Y sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__a22oi_1_201/Y sky130_fd_sc_hd__xor2_1_203/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_399 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_330/A sky130_fd_sc_hd__nor2_2_15/Y
+ sky130_fd_sc_hd__nand2_1_399/Y sky130_fd_sc_hd__xnor2_1_91/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_809 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_704 sky130_fd_sc_hd__xor2_1_650/B sky130_fd_sc_hd__nand2_1_705/Y
+ sky130_fd_sc_hd__nand2_1_704/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_715 sky130_fd_sc_hd__o22ai_1_96/B2 sky130_fd_sc_hd__xnor2_2_4/Y
+ sky130_fd_sc_hd__xor2_1_667/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_13 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_13/A1 sky130_fd_sc_hd__buf_2_70/X
+ sky130_fd_sc_hd__mux2_8_1/S sky130_fd_sc_hd__fa_2_415/A vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_726 sky130_fd_sc_hd__nand2_1_726/Y sky130_fd_sc_hd__nor2_1_235/A
+ sky130_fd_sc_hd__xor2_1_660/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_24 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_24/A1 sky130_fd_sc_hd__buf_4_22/X
+ sky130_fd_sc_hd__mux2_8_1/S sky130_fd_sc_hd__mux2_2_24/X vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_737 sky130_fd_sc_hd__xor2_1_655/B sky130_fd_sc_hd__nand2_1_738/Y
+ sky130_fd_sc_hd__or2_0_90/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_35 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_35/A1 sky130_fd_sc_hd__buf_2_89/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__mux2_2_35/X vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_748 sky130_fd_sc_hd__nand2_1_748/Y sky130_fd_sc_hd__nor2_1_240/A
+ sky130_fd_sc_hd__nor2_1_240/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_46 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_46/A1 sky130_fd_sc_hd__buf_2_150/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__mux2_2_46/X vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_759 sky130_fd_sc_hd__xnor2_1_214/A sky130_fd_sc_hd__nand2_1_775/Y
+ sky130_fd_sc_hd__nand2_1_759/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__conb_1_110 sky130_fd_sc_hd__conb_1_110/LO sky130_fd_sc_hd__conb_1_110/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_121 sky130_fd_sc_hd__conb_1_121/LO sky130_fd_sc_hd__conb_1_121/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_132 sky130_fd_sc_hd__conb_1_132/LO sky130_fd_sc_hd__conb_1_132/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_143 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__conb_1_143/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__dfxtp_1_500 la_data_out[35] sky130_fd_sc_hd__dfxtp_1_509/CLK sky130_fd_sc_hd__and2_0_400/X
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_160 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__xor2_1_160/X
+ sky130_fd_sc_hd__xor2_1_160/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1808 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_511 la_data_out[34] sky130_fd_sc_hd__dfxtp_1_520/CLK sky130_fd_sc_hd__and2_0_344/X
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_171 sky130_fd_sc_hd__xor2_1_171/B sky130_fd_sc_hd__xor2_1_171/X
+ sky130_fd_sc_hd__xor2_1_171/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1819 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_522 wbs_dat_o[1] sky130_fd_sc_hd__dfxtp_1_532/CLK sky130_fd_sc_hd__nor2b_1_156/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_182 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__xor2_1_182/X
+ sky130_fd_sc_hd__xor2_1_182/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_533 wbs_dat_o[12] sky130_fd_sc_hd__dfxtp_1_533/CLK sky130_fd_sc_hd__nor2b_1_145/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_193 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__fa_2_136/B
+ sky130_fd_sc_hd__xor2_1_193/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_544 wbs_dat_o[23] sky130_fd_sc_hd__dfxtp_1_544/CLK sky130_fd_sc_hd__nor2b_1_134/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_120 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_120/X sky130_fd_sc_hd__inv_4_5/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_131 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_131/X sky130_fd_sc_hd__buf_2_135/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_202 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__nor2_2_5/A
+ sky130_fd_sc_hd__nor2_2_5/B sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__nor2_2_4/B
+ sky130_fd_sc_hd__o21ai_1_373/B1 sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_142 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_142/X sky130_fd_sc_hd__clkinv_1_862/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_213 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__or2_0_52/B
+ sky130_fd_sc_hd__or2_0_53/A sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__buf_2_32/X
+ sky130_fd_sc_hd__o21ai_1_392/B1 sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_153 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_28/A1 sky130_fd_sc_hd__clkbuf_1_153/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_0 sky130_fd_sc_hd__dfxtp_1_0/Q sky130_fd_sc_hd__dfxtp_1_0/CLK
+ sky130_fd_sc_hd__nor2b_1_0/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a222oi_1_224 vccd1 vssd1 sky130_fd_sc_hd__and3_4_16/X sky130_fd_sc_hd__and2_0_49/A
+ sky130_fd_sc_hd__and2_0_45/A sky130_fd_sc_hd__nor2_2_19/Y sky130_fd_sc_hd__and2_0_87/A
+ sky130_fd_sc_hd__o21ai_1_415/B1 sky130_fd_sc_hd__nor2b_2_3/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_164 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_255/A sky130_fd_sc_hd__clkbuf_1_60/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_235 vccd1 vssd1 sky130_fd_sc_hd__and3_1_1/X sky130_fd_sc_hd__or2_0_52/B
+ sky130_fd_sc_hd__or2_0_53/A sky130_fd_sc_hd__nor2_1_117/Y sky130_fd_sc_hd__buf_2_32/X
+ sky130_fd_sc_hd__o21ai_1_429/B1 sky130_fd_sc_hd__nor2b_1_8/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_175 vssd1 vccd1 sky130_fd_sc_hd__a22o_1_26/B2 sky130_fd_sc_hd__clkbuf_1_175/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_246 vccd1 vssd1 sky130_fd_sc_hd__and3_4_9/X sky130_fd_sc_hd__or2_0_42/B
+ sky130_fd_sc_hd__or2_0_39/B sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__or2_0_58/A
+ sky130_fd_sc_hd__o21ai_1_442/B1 sky130_fd_sc_hd__and2b_4_5/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_186 vssd1 vccd1 sky130_fd_sc_hd__buf_12_59/A sky130_fd_sc_hd__clkinv_1_948/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_257 vccd1 vssd1 sky130_fd_sc_hd__and3_4_13/X sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__buf_2_32/X sky130_fd_sc_hd__nor2_1_121/Y sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__o21ai_1_458/B1 sky130_fd_sc_hd__nor2b_1_9/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_197 vssd1 vccd1 sky130_fd_sc_hd__buf_8_58/A sky130_fd_sc_hd__clkbuf_1_197/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_405 sky130_fd_sc_hd__nor2_1_203/A sky130_fd_sc_hd__nor2_1_206/B
+ sky130_fd_sc_hd__fa_2_405/A sky130_fd_sc_hd__fa_2_405/B sky130_fd_sc_hd__fa_2_405/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_268 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__or2_0_66/A sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__or2_0_60/B
+ sky130_fd_sc_hd__o21ai_1_470/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_416 sky130_fd_sc_hd__fa_2_415/CIN sky130_fd_sc_hd__fa_2_416/SUM
+ sky130_fd_sc_hd__fa_2_416/A sky130_fd_sc_hd__fa_2_416/B sky130_fd_sc_hd__fa_2_416/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a222oi_1_279 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__buf_4_4/X sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__o21ai_1_485/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_427 sky130_fd_sc_hd__fa_2_421/B sky130_fd_sc_hd__fa_2_422/A
+ sky130_fd_sc_hd__fa_2_427/A sky130_fd_sc_hd__fa_2_427/B sky130_fd_sc_hd__fa_2_427/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_438 sky130_fd_sc_hd__or2_0_94/A sky130_fd_sc_hd__or2_0_93/B
+ sky130_fd_sc_hd__fa_2_438/A sky130_fd_sc_hd__fa_2_438/B sky130_fd_sc_hd__fa_2_441/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_449 sky130_fd_sc_hd__fah_1_18/A sky130_fd_sc_hd__fa_2_421/A
+ sky130_fd_sc_hd__fa_2_449/A sky130_fd_sc_hd__fa_2_449/B sky130_fd_sc_hd__fa_2_449/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_4_10 sky130_fd_sc_hd__inv_4_10/Y sky130_fd_sc_hd__inv_4_10/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__inv_4_21 sky130_fd_sc_hd__inv_4_21/Y wbs_dat_i[6] vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__and2_0_140 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_38/D sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_140/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_151 vccd1 vssd1 sky130_fd_sc_hd__and2_0_151/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_151/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_162 vccd1 vssd1 sky130_fd_sc_hd__and2_0_162/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_162/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_70 io_out[31] sky130_fd_sc_hd__conb_1_72/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_173 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_47/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_173/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_81 io_out[20] sky130_fd_sc_hd__conb_1_61/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_184 vccd1 vssd1 sky130_fd_sc_hd__and2_0_184/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_184/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_92 io_out[9] sky130_fd_sc_hd__conb_1_50/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_195 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_49/D sky130_fd_sc_hd__o21ai_2_0/B1
+ sky130_fd_sc_hd__o21ai_1_86/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__sdlclkp_1_1 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_8_4/Y
+ sky130_fd_sc_hd__clkinv_2_9/A sky130_fd_sc_hd__o21ai_2_3/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__sdlclkp_1
Xsky130_fd_sc_hd__o21ai_1_130 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_133/A2 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_132/Y sky130_fd_sc_hd__and2_0_140/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_141 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_141/A2 sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__a22oi_1_181/Y sky130_fd_sc_hd__and2_0_127/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_152 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_153/A2 sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__a22oi_1_186/Y sky130_fd_sc_hd__and2_0_112/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_163 vssd1 vccd1 sky130_fd_sc_hd__a21oi_2_4/Y sky130_fd_sc_hd__nor2_1_65/Y
+ sky130_fd_sc_hd__nand2_1_218/Y sky130_fd_sc_hd__xnor2_1_23/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_174 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_207/A2 sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__a222oi_1_55/Y sky130_fd_sc_hd__xor2_1_7/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_185 vssd1 vccd1 sky130_fd_sc_hd__inv_2_24/Y sky130_fd_sc_hd__nand2b_1_1/Y
+ sky130_fd_sc_hd__a222oi_1_64/Y sky130_fd_sc_hd__xor2_1_16/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_196 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_261/A2 sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__a222oi_1_72/Y sky130_fd_sc_hd__xor2_1_25/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_19 vccd1 vssd1 sky130_fd_sc_hd__nand2_1_135/A sky130_fd_sc_hd__nor2_4_7/Y
+ sky130_fd_sc_hd__xnor2_1_179/Y sky130_fd_sc_hd__xnor2_1_54/Y sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__a222oi_1_19/Y sky130_fd_sc_hd__buf_2_17/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_606 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_617 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_501 sky130_fd_sc_hd__nand2_1_501/Y sky130_fd_sc_hd__nor2_4_15/Y
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_628 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_512 sky130_fd_sc_hd__nand2_1_512/Y sky130_fd_sc_hd__or2_1_9/A
+ sky130_fd_sc_hd__or2_1_9/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_639 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_523 sky130_fd_sc_hd__nand2_1_523/Y sky130_fd_sc_hd__or2_1_8/A
+ sky130_fd_sc_hd__or2_1_8/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_534 sky130_fd_sc_hd__nand2_1_534/Y sky130_fd_sc_hd__or2_1_7/A
+ sky130_fd_sc_hd__or2_1_7/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_545 sky130_fd_sc_hd__nand2_1_545/Y sky130_fd_sc_hd__or2_1_6/A
+ sky130_fd_sc_hd__or2_1_6/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_556 sky130_fd_sc_hd__nand2_1_556/Y sky130_fd_sc_hd__or2_1_5/A
+ sky130_fd_sc_hd__or2_1_5/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_567 sky130_fd_sc_hd__nand2_1_567/Y sky130_fd_sc_hd__or2_0_63/X
+ sky130_fd_sc_hd__nor2_1_184/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_3 sky130_fd_sc_hd__and3_1_0/C sky130_fd_sc_hd__nor2b_1_3/Y
+ sky130_fd_sc_hd__and3_1_0/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nand2_1_578 sky130_fd_sc_hd__nand2_1_578/Y sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__nor2_1_73/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_589 sky130_fd_sc_hd__xnor2_1_163/A sky130_fd_sc_hd__nand2_1_590/Y
+ sky130_fd_sc_hd__nand2_1_589/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_1103 sky130_fd_sc_hd__clkinv_4_46/A sky130_fd_sc_hd__a22o_1_23/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1114 sky130_fd_sc_hd__clkinv_4_57/A sky130_fd_sc_hd__a22o_1_34/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1125 sky130_fd_sc_hd__clkinv_4_68/A sky130_fd_sc_hd__a22o_1_45/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1136 sky130_fd_sc_hd__and2_4_0/B sky130_fd_sc_hd__clkinv_1_846/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1147 sky130_fd_sc_hd__buf_2_42/A sky130_fd_sc_hd__inv_4_19/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1605 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1616 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1627 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_330 sky130_fd_sc_hd__dfxtp_1_330/Q sky130_fd_sc_hd__dfxtp_1_343/CLK
+ sky130_fd_sc_hd__and2_0_319/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1638 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_341 sky130_fd_sc_hd__dfxtp_1_341/Q sky130_fd_sc_hd__dfxtp_1_343/CLK
+ sky130_fd_sc_hd__and2_0_329/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1649 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_352 sky130_fd_sc_hd__dfxtp_1_352/Q sky130_fd_sc_hd__dfxtp_1_354/CLK
+ sky130_fd_sc_hd__and2_0_314/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_363 sky130_fd_sc_hd__dfxtp_1_363/Q sky130_fd_sc_hd__dfxtp_1_29/CLK
+ sky130_fd_sc_hd__or4_1_1/C vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_374 sky130_fd_sc_hd__dfxtp_1_374/Q sky130_fd_sc_hd__dfxtp_1_375/CLK
+ sky130_fd_sc_hd__nor2b_1_109/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_385 sky130_fd_sc_hd__dfxtp_1_385/Q sky130_fd_sc_hd__dfxtp_1_395/CLK
+ sky130_fd_sc_hd__nor2b_1_98/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_5 sky130_fd_sc_hd__nand2_2_0/A sky130_fd_sc_hd__nand2_1_7/B
+ sky130_fd_sc_hd__or2_0_84/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_396 sky130_fd_sc_hd__dfxtp_1_396/Q sky130_fd_sc_hd__dfxtp_1_423/CLK
+ sky130_fd_sc_hd__nor2b_1_119/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_202 sky130_fd_sc_hd__fa_2_197/CIN sky130_fd_sc_hd__fa_2_208/A
+ sky130_fd_sc_hd__fa_2_202/A sky130_fd_sc_hd__fa_2_202/B sky130_fd_sc_hd__fa_2_202/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_213 sky130_fd_sc_hd__fa_2_202/CIN sky130_fd_sc_hd__fa_2_213/SUM
+ sky130_fd_sc_hd__fa_2_213/A sky130_fd_sc_hd__fa_2_213/B sky130_fd_sc_hd__xor2_1_310/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_224 sky130_fd_sc_hd__fa_2_220/CIN sky130_fd_sc_hd__fa_2_227/B
+ sky130_fd_sc_hd__fa_2_224/A sky130_fd_sc_hd__fa_2_224/B sky130_fd_sc_hd__xor2_1_327/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_235 sky130_fd_sc_hd__fa_2_231/CIN sky130_fd_sc_hd__fa_2_240/A
+ sky130_fd_sc_hd__fa_2_235/A sky130_fd_sc_hd__fa_2_235/B sky130_fd_sc_hd__xor2_1_341/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_246 sky130_fd_sc_hd__fa_2_244/B sky130_fd_sc_hd__fa_2_247/A
+ sky130_fd_sc_hd__fa_2_246/A sky130_fd_sc_hd__fa_2_246/B sky130_fd_sc_hd__fa_2_246/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_257 sky130_fd_sc_hd__fa_2_255/B sky130_fd_sc_hd__fa_2_259/CIN
+ sky130_fd_sc_hd__fa_2_257/A sky130_fd_sc_hd__fa_2_257/B sky130_fd_sc_hd__xor2_1_373/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_268 sky130_fd_sc_hd__fa_2_266/B sky130_fd_sc_hd__fa_2_269/CIN
+ sky130_fd_sc_hd__fa_2_268/A sky130_fd_sc_hd__fa_2_268/B sky130_fd_sc_hd__xor2_1_390/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_279 sky130_fd_sc_hd__fa_2_278/CIN sky130_fd_sc_hd__or2_0_49/B
+ sky130_fd_sc_hd__fa_2_279/A sky130_fd_sc_hd__fa_2_279/B sky130_fd_sc_hd__xor2_1_412/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_6 vccd1 vssd1 sky130_fd_sc_hd__and2_0_6/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_6/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__fa_2_60 sky130_fd_sc_hd__fa_2_55/CIN sky130_fd_sc_hd__fa_2_66/A
+ sky130_fd_sc_hd__fa_2_60/A sky130_fd_sc_hd__fa_2_60/B sky130_fd_sc_hd__fa_2_60/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_71 sky130_fd_sc_hd__fa_2_60/CIN sky130_fd_sc_hd__fa_2_71/SUM
+ sky130_fd_sc_hd__fa_2_71/A sky130_fd_sc_hd__fa_2_71/B sky130_fd_sc_hd__xor2_1_97/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_82 sky130_fd_sc_hd__fa_2_78/CIN sky130_fd_sc_hd__fa_2_85/B
+ sky130_fd_sc_hd__fa_2_82/A sky130_fd_sc_hd__fa_2_82/B sky130_fd_sc_hd__fa_2_82/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_93 sky130_fd_sc_hd__fa_2_89/CIN sky130_fd_sc_hd__fa_2_98/A
+ sky130_fd_sc_hd__fa_2_93/A sky130_fd_sc_hd__fa_2_93/B sky130_fd_sc_hd__fa_2_93/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a21oi_1_10 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_39/Y
+ sky130_fd_sc_hd__a21oi_1_10/Y sky130_fd_sc_hd__dfxtp_1_94/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_21 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_50/Y
+ sky130_fd_sc_hd__a21oi_1_21/Y sky130_fd_sc_hd__dfxtp_1_76/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_32 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_61/Y
+ sky130_fd_sc_hd__a21oi_1_32/Y sky130_fd_sc_hd__dfxtp_1_63/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_43 sky130_fd_sc_hd__a21oi_1_45/A1 sky130_fd_sc_hd__o21ai_1_239/Y
+ sky130_fd_sc_hd__a21oi_1_43/Y sky130_fd_sc_hd__nor2_1_57/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_207 sky130_fd_sc_hd__buf_6_69/X sky130_fd_sc_hd__buf_12_207/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_54 sky130_fd_sc_hd__a21oi_1_54/A1 sky130_fd_sc_hd__a21oi_1_54/B1
+ sky130_fd_sc_hd__a21oi_1_54/Y sky130_fd_sc_hd__nand2_1_263/A vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_218 sky130_fd_sc_hd__buf_6_36/X sky130_fd_sc_hd__buf_12_286/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_65 sky130_fd_sc_hd__nand2_1_312/Y sky130_fd_sc_hd__nand2_1_301/Y
+ sky130_fd_sc_hd__a21oi_1_65/Y sky130_fd_sc_hd__nor2_1_100/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_229 sky130_fd_sc_hd__buf_6_63/X sky130_fd_sc_hd__buf_12_337/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_76 sky130_fd_sc_hd__a21oi_1_80/A1 sky130_fd_sc_hd__o21ai_1_444/Y
+ sky130_fd_sc_hd__a21oi_1_76/Y sky130_fd_sc_hd__nor2_1_113/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_87 sky130_fd_sc_hd__a21oi_1_89/A1 sky130_fd_sc_hd__nand2_1_421/Y
+ sky130_fd_sc_hd__a21oi_1_87/Y sky130_fd_sc_hd__nor2_1_136/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_98 sky130_fd_sc_hd__xnor2_1_119/B sky130_fd_sc_hd__a21oi_1_98/B1
+ sky130_fd_sc_hd__xnor2_1_65/A sky130_fd_sc_hd__nand2_1_473/A vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__inv_1_0 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__inv_1_0/A vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__nor3_1_2 sky130_fd_sc_hd__or4_1_3/X sky130_fd_sc_hd__nor3_1_2/Y
+ sky130_fd_sc_hd__ha_2_42/A sky130_fd_sc_hd__ha_2_43/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__clkinv_1_407 sky130_fd_sc_hd__or2b_2_0/A sky130_fd_sc_hd__dfxtp_1_247/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_418 sky130_fd_sc_hd__nor2_1_106/A sky130_fd_sc_hd__nand2_1_349/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_429 sky130_fd_sc_hd__nand2_1_355/A sky130_fd_sc_hd__nor2_2_11/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_50 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_61 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_72 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_83 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_94 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_50 vccd1 vssd1 sky130_fd_sc_hd__buf_6_50/X sky130_fd_sc_hd__buf_6_50/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_61 vccd1 vssd1 sky130_fd_sc_hd__buf_6_61/X sky130_fd_sc_hd__buf_8_2/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_72 vccd1 vssd1 sky130_fd_sc_hd__buf_6_72/X sky130_fd_sc_hd__buf_8_29/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_83 vccd1 vssd1 sky130_fd_sc_hd__buf_6_83/X sky130_fd_sc_hd__buf_6_83/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_94 vccd1 vssd1 la_data_out[77] sky130_fd_sc_hd__or2_0_83/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_30 sky130_fd_sc_hd__clkinv_4_67/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_41 sky130_fd_sc_hd__buf_2_193/A vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_52 sky130_fd_sc_hd__buf_2_189/A vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_63 sky130_fd_sc_hd__dfxtp_1_12/Q vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a222oi_1_7 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_348/Q sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__o211ai_1_23/Y sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__a222oi_1_7/Y sky130_fd_sc_hd__dfxtp_1_299/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_403 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_414 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_425 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_436 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_320 sky130_fd_sc_hd__xnor2_1_62/A sky130_fd_sc_hd__nand2_1_321/Y
+ sky130_fd_sc_hd__or2_0_24/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_447 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_331 sky130_fd_sc_hd__nand2_1_331/Y sky130_fd_sc_hd__nor2_4_11/Y
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_458 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_930 sky130_fd_sc_hd__buf_8_18/A sky130_fd_sc_hd__inv_2_120/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_342 sky130_fd_sc_hd__xnor2_1_70/A sky130_fd_sc_hd__nand2_1_343/Y
+ sky130_fd_sc_hd__or2_0_36/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_469 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_941 sky130_fd_sc_hd__buf_8_29/A sky130_fd_sc_hd__clkinv_1_941/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_353 sky130_fd_sc_hd__xnor2_1_74/A sky130_fd_sc_hd__nand2_1_354/Y
+ sky130_fd_sc_hd__or2_0_39/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_952 sky130_fd_sc_hd__inv_2_148/A sky130_fd_sc_hd__buf_8_2/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_364 sky130_fd_sc_hd__xnor2_1_79/A sky130_fd_sc_hd__nand2_1_365/Y
+ sky130_fd_sc_hd__or2_0_42/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_963 sky130_fd_sc_hd__clkinv_4_21/A sky130_fd_sc_hd__nand2_1_846/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_375 sky130_fd_sc_hd__xnor2_1_83/A sky130_fd_sc_hd__nand2_1_376/Y
+ sky130_fd_sc_hd__or2_0_40/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_974 sky130_fd_sc_hd__buf_2_131/A sky130_fd_sc_hd__clkinv_4_93/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_386 sky130_fd_sc_hd__xnor2_1_87/A sky130_fd_sc_hd__nand2_1_387/Y
+ sky130_fd_sc_hd__or2_0_46/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_985 sky130_fd_sc_hd__clkinv_1_985/Y sky130_fd_sc_hd__clkinv_4_29/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_397 sky130_fd_sc_hd__nand2_1_397/Y sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__buf_4_4/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_996 sky130_fd_sc_hd__clkinv_1_996/Y sky130_fd_sc_hd__clkinv_1_996/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1402 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1413 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1424 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1435 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1446 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1457 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_160 sky130_fd_sc_hd__dfxtp_1_160/Q sky130_fd_sc_hd__dfxtp_1_176/CLK
+ sky130_fd_sc_hd__and2_0_108/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1468 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_171 sky130_fd_sc_hd__dfxtp_1_171/Q sky130_fd_sc_hd__dfxtp_1_177/CLK
+ sky130_fd_sc_hd__and2_0_162/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1479 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_182 sky130_fd_sc_hd__dfxtp_1_182/Q sky130_fd_sc_hd__clkinv_4_2/Y
+ sky130_fd_sc_hd__and2_0_217/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_193 sky130_fd_sc_hd__xnor2_1_186/A sky130_fd_sc_hd__dfxtp_4_3/CLK
+ sky130_fd_sc_hd__and2_0_35/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_2_19 vccd1 vssd1 sky130_fd_sc_hd__buf_2_19/X sky130_fd_sc_hd__buf_2_4/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_970 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_981 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_992 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o211ai_1_13 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_50/B1
+ sky130_fd_sc_hd__a22oi_1_4/A2 sky130_fd_sc_hd__a22oi_1_58/Y sky130_fd_sc_hd__a22oi_1_59/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_24 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_38/B1
+ sky130_fd_sc_hd__o211ai_1_24/Y sky130_fd_sc_hd__a22oi_1_80/Y sky130_fd_sc_hd__a22oi_1_81/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_35 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o21ai_1_5/A2
+ sky130_fd_sc_hd__ha_2_2/B sky130_fd_sc_hd__nand2_1_55/Y sky130_fd_sc_hd__a21oi_1_6/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_46 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o22ai_1_17/B1
+ sky130_fd_sc_hd__fa_2_382/A sky130_fd_sc_hd__nand2_1_66/Y sky130_fd_sc_hd__a21oi_1_17/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_57 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o22ai_1_6/B1
+ sky130_fd_sc_hd__fa_2_410/B sky130_fd_sc_hd__nand2_1_77/Y sky130_fd_sc_hd__a21oi_1_28/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__clkinv_1_204 sky130_fd_sc_hd__o22ai_1_14/B1 sky130_fd_sc_hd__dfxtp_1_109/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_215 sky130_fd_sc_hd__nor2_1_14/A sky130_fd_sc_hd__dfxtp_1_137/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_226 sky130_fd_sc_hd__o22ai_1_6/A2 sky130_fd_sc_hd__dfxtp_1_165/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_237 sky130_fd_sc_hd__o22ai_1_3/B1 sky130_fd_sc_hd__dfxtp_1_98/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_248 sky130_fd_sc_hd__o21ai_1_81/A2 sky130_fd_sc_hd__xnor2_1_154/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_259 sky130_fd_sc_hd__o21ai_1_125/A2 sky130_fd_sc_hd__xnor2_1_175/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_2_4 sky130_fd_sc_hd__buf_2_16/A sky130_fd_sc_hd__o21ai_2_4/Y
+ sky130_fd_sc_hd__o21ai_2_4/A2 sky130_fd_sc_hd__a21oi_1_2/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__o21ai_2
Xsky130_fd_sc_hd__and3_4_17 sky130_fd_sc_hd__nor2_2_20/B sky130_fd_sc_hd__nor2b_2_4/A
+ sky130_fd_sc_hd__nor2_2_20/A sky130_fd_sc_hd__and3_4_17/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__a21oi_1_101 sky130_fd_sc_hd__xnor2_1_120/B sky130_fd_sc_hd__a21oi_1_99/A2
+ sky130_fd_sc_hd__xor2_1_411/A sky130_fd_sc_hd__or2_0_50/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_112 sky130_fd_sc_hd__clkinv_1_549/Y sky130_fd_sc_hd__o21ai_1_693/Y
+ sky130_fd_sc_hd__a21oi_1_112/Y sky130_fd_sc_hd__nor2_1_172/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_123 sky130_fd_sc_hd__xnor2_1_166/B sky130_fd_sc_hd__o21ai_1_633/Y
+ sky130_fd_sc_hd__xor2_1_572/A sky130_fd_sc_hd__nor2_2_28/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_134 sky130_fd_sc_hd__or2_0_69/X sky130_fd_sc_hd__clkinv_1_603/Y
+ sky130_fd_sc_hd__a21oi_1_134/Y sky130_fd_sc_hd__clkinv_1_606/Y vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_145 sky130_fd_sc_hd__xnor2_1_195/B sky130_fd_sc_hd__clkinv_1_639/Y
+ sky130_fd_sc_hd__xor2_1_646/A sky130_fd_sc_hd__or2_0_79/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_156 sky130_fd_sc_hd__xnor2_1_209/B sky130_fd_sc_hd__clkinv_1_671/Y
+ sky130_fd_sc_hd__a21oi_1_156/Y sky130_fd_sc_hd__or2_0_88/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_167 sky130_fd_sc_hd__xnor2_1_217/B sky130_fd_sc_hd__clkinv_1_696/Y
+ sky130_fd_sc_hd__xor2_1_665/B sky130_fd_sc_hd__or2_0_96/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_178 sky130_fd_sc_hd__xnor2_1_299/B sky130_fd_sc_hd__clkinv_1_824/Y
+ sky130_fd_sc_hd__xor2_1_684/A sky130_fd_sc_hd__or2_0_108/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_189 sky130_fd_sc_hd__a21o_2_0/A2 sky130_fd_sc_hd__maj3_1_0/X
+ sky130_fd_sc_hd__a21oi_1_189/Y sky130_fd_sc_hd__o211ai_1_64/Y vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_108 sky130_fd_sc_hd__buf_8_108/A sky130_fd_sc_hd__buf_6_57/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_119 sky130_fd_sc_hd__inv_2_113/Y sky130_fd_sc_hd__buf_8_159/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_12_560 sky130_fd_sc_hd__buf_12_560/A sky130_fd_sc_hd__buf_12_560/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_571 sky130_fd_sc_hd__buf_12_571/A sky130_fd_sc_hd__buf_12_571/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_200 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_582 sky130_fd_sc_hd__buf_12_582/A sky130_fd_sc_hd__buf_12_582/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_211 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_593 sky130_fd_sc_hd__buf_12_593/A sky130_fd_sc_hd__buf_12_593/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_222 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_233 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_244 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_255 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_266 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_301 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_301/B sky130_fd_sc_hd__xnor2_1_301/Y
+ sky130_fd_sc_hd__xnor2_1_301/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_150 sky130_fd_sc_hd__nor2_4_6/A sky130_fd_sc_hd__ha_2_9/B
+ sky130_fd_sc_hd__ha_2_9/SUM vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_277 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_161 sky130_fd_sc_hd__nand2_1_161/Y sky130_fd_sc_hd__nor2_4_8/Y
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_288 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_760 sky130_fd_sc_hd__fa_2_483/A sky130_fd_sc_hd__clkinv_1_760/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_172 sky130_fd_sc_hd__nand2_1_172/Y sky130_fd_sc_hd__or2_0_9/A
+ sky130_fd_sc_hd__or2_0_9/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_299 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_771 sky130_fd_sc_hd__ha_2_18/B sky130_fd_sc_hd__clkinv_1_771/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_183 sky130_fd_sc_hd__nand2_1_183/Y sky130_fd_sc_hd__or2_0_58/A
+ sky130_fd_sc_hd__or2_0_58/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_782 sky130_fd_sc_hd__and2_0_325/A sky130_fd_sc_hd__clkinv_1_782/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_194 sky130_fd_sc_hd__nand2_1_194/Y sky130_fd_sc_hd__or2_0_61/A
+ sky130_fd_sc_hd__or2_0_42/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_793 sky130_fd_sc_hd__and2_0_314/A sky130_fd_sc_hd__clkinv_1_793/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1210 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1221 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1232 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1243 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1254 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1265 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1276 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_707 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_733/A2 sky130_fd_sc_hd__nand2b_2_8/Y
+ sky130_fd_sc_hd__o21ai_1_707/B1 sky130_fd_sc_hd__xor2_1_486/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1287 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_718 vssd1 vccd1 sky130_fd_sc_hd__nand2_2_13/Y sky130_fd_sc_hd__nand2b_1_19/Y
+ sky130_fd_sc_hd__a22oi_1_215/Y sky130_fd_sc_hd__xor2_1_495/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1298 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_729 vssd1 vccd1 sky130_fd_sc_hd__inv_2_51/Y sky130_fd_sc_hd__nand2b_2_6/Y
+ sky130_fd_sc_hd__o21ai_1_729/B1 sky130_fd_sc_hd__xor2_1_506/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_14 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__fa_2_8/A
+ sky130_fd_sc_hd__xor2_1_14/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__and3_1_1 vssd1 vccd1 sky130_fd_sc_hd__and3_1_1/X sky130_fd_sc_hd__and3_1_1/B
+ sky130_fd_sc_hd__and3_1_1/A sky130_fd_sc_hd__and3_1_1/C vssd1 vccd1 sky130_fd_sc_hd__and3_1
Xsky130_fd_sc_hd__xor2_1_25 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__fa_2_10/B
+ sky130_fd_sc_hd__xor2_1_25/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_36 sky130_fd_sc_hd__fa_2_75/A sky130_fd_sc_hd__xor2_1_36/X
+ sky130_fd_sc_hd__xor2_1_36/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_47 sky130_fd_sc_hd__fa_2_56/A sky130_fd_sc_hd__fa_2_30/B
+ sky130_fd_sc_hd__xor2_1_47/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_58 sky130_fd_sc_hd__fa_2_56/A sky130_fd_sc_hd__xor2_1_58/X
+ sky130_fd_sc_hd__xor2_1_58/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_69 sky130_fd_sc_hd__fa_2_56/A sky130_fd_sc_hd__fa_2_45/B
+ sky130_fd_sc_hd__xor2_1_69/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2b_1_8 sky130_fd_sc_hd__nand2b_1_8/Y sky130_fd_sc_hd__nor2_2_19/A
+ sky130_fd_sc_hd__nor2_2_19/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__xor2_1_501 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__xor2_1_501/X
+ sky130_fd_sc_hd__xor2_1_501/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a21o_2_4 sky130_fd_sc_hd__a21o_2_4/X sky130_fd_sc_hd__a21o_2_4/B1
+ wbs_adr_i[9] sky130_fd_sc_hd__a21o_2_4/A2 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__xor2_1_512 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__xor2_1_512/X
+ sky130_fd_sc_hd__xor2_1_512/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_523 sky130_fd_sc_hd__fah_1_14/A sky130_fd_sc_hd__xor2_1_523/X
+ sky130_fd_sc_hd__xor2_1_523/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_534 sky130_fd_sc_hd__fah_1_14/A sky130_fd_sc_hd__fa_2_361/A
+ sky130_fd_sc_hd__xor2_1_534/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_545 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__fa_2_370/B
+ sky130_fd_sc_hd__xor2_1_545/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_556 sky130_fd_sc_hd__fa_2_379/A sky130_fd_sc_hd__xor2_1_556/X
+ sky130_fd_sc_hd__xor2_1_556/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_567 sky130_fd_sc_hd__fah_1_14/A sky130_fd_sc_hd__fa_2_384/B
+ sky130_fd_sc_hd__xor2_1_567/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_578 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__fa_2_388/B
+ sky130_fd_sc_hd__xor2_1_578/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_589 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__fa_2_396/B
+ sky130_fd_sc_hd__xor2_1_589/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__ha_2_30 vssd1 vccd1 sky130_fd_sc_hd__ha_2_30/A sky130_fd_sc_hd__ha_2_29/B
+ sky130_fd_sc_hd__ha_2_30/SUM sky130_fd_sc_hd__ha_2_30/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_41 vssd1 vccd1 sky130_fd_sc_hd__or4_1_3/A sky130_fd_sc_hd__ha_2_40/B
+ sky130_fd_sc_hd__ha_2_41/SUM sky130_fd_sc_hd__ha_2_41/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__and2b_4_3 sky130_fd_sc_hd__nor2_2_9/A sky130_fd_sc_hd__and2b_4_3/X
+ sky130_fd_sc_hd__and3_4_1/C vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__and2b_4
Xsky130_fd_sc_hd__ha_2_52 vssd1 vccd1 sky130_fd_sc_hd__ha_2_52/A sky130_fd_sc_hd__ha_2_51/B
+ sky130_fd_sc_hd__ha_2_52/SUM sky130_fd_sc_hd__ha_2_52/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_4 vssd1 vccd1 sky130_fd_sc_hd__fa_2_250/A sky130_fd_sc_hd__xor2_1_362/B
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__nor2_1_150 sky130_fd_sc_hd__buf_2_19/X sky130_fd_sc_hd__nor2_1_150/Y
+ sky130_fd_sc_hd__buf_6_5/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_1_4 la_data_out[123] sky130_fd_sc_hd__clkinv_1_4/A vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_161 sky130_fd_sc_hd__inv_6_0/Y sky130_fd_sc_hd__nor2_1_161/Y
+ sky130_fd_sc_hd__buf_8_0/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_172 sky130_fd_sc_hd__nor2_1_175/B sky130_fd_sc_hd__nor2_1_172/Y
+ sky130_fd_sc_hd__nor2_1_172/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_183 sky130_fd_sc_hd__and3_4_24/A sky130_fd_sc_hd__nor2_1_183/Y
+ sky130_fd_sc_hd__and3_4_24/C vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_194 sky130_fd_sc_hd__nor2_2_10/B sky130_fd_sc_hd__nor2_1_194/Y
+ sky130_fd_sc_hd__nor2_1_85/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_70 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__nor2_4_3/Y
+ sky130_fd_sc_hd__nand2_1_64/B sky130_fd_sc_hd__dfxtp_1_146/Q sky130_fd_sc_hd__a22oi_1_70/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_81 sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__dfxtp_1_119/Q sky130_fd_sc_hd__dfxtp_1_87/Q sky130_fd_sc_hd__a22oi_1_81/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_92 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__nor2_4_3/Y
+ sky130_fd_sc_hd__nand2_1_55/B sky130_fd_sc_hd__dfxtp_1_157/Q sky130_fd_sc_hd__a22oi_1_92/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__and2_0_19 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_4_2/D sky130_fd_sc_hd__and2_0_99/B
+ sky130_fd_sc_hd__buf_2_32/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_12_390 sky130_fd_sc_hd__buf_12_390/A sky130_fd_sc_hd__buf_12_471/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xnor2_1_120 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_120/B sky130_fd_sc_hd__xnor2_1_120/Y
+ sky130_fd_sc_hd__xnor2_1_120/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__buf_8_18 sky130_fd_sc_hd__buf_8_18/A sky130_fd_sc_hd__buf_8_18/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xnor2_1_131 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_131/B sky130_fd_sc_hd__xnor2_1_131/Y
+ sky130_fd_sc_hd__xnor2_1_131/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__buf_8_29 sky130_fd_sc_hd__buf_8_29/A sky130_fd_sc_hd__buf_8_29/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xnor2_1_142 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_142/B sky130_fd_sc_hd__xnor2_1_142/Y
+ sky130_fd_sc_hd__xnor2_1_142/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_590 sky130_fd_sc_hd__nand2_1_615/A sky130_fd_sc_hd__nor2_1_202/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_153 vssd1 vccd1 sky130_fd_sc_hd__fa_2_379/A sky130_fd_sc_hd__and3_4_24/C
+ sky130_fd_sc_hd__xnor2_1_153/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_164 vssd1 vccd1 sky130_fd_sc_hd__fah_1_14/A sky130_fd_sc_hd__nor2_2_31/A
+ sky130_fd_sc_hd__xnor2_1_164/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_175 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_175/B sky130_fd_sc_hd__xnor2_1_175/Y
+ sky130_fd_sc_hd__xnor2_1_175/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_186 vssd1 vccd1 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__nor2_4_18/A
+ sky130_fd_sc_hd__xnor2_1_186/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_197 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_197/B sky130_fd_sc_hd__and2_0_259/A
+ sky130_fd_sc_hd__xnor2_1_197/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_4_70 sky130_fd_sc_hd__clkinv_4_70/A sky130_fd_sc_hd__clkinv_4_70/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_81 wbs_dat_i[25] sky130_fd_sc_hd__clkinv_4_81/Y vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_92 sky130_fd_sc_hd__nand2_1_13/Y sky130_fd_sc_hd__inv_2_153/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_1040 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1051 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1062 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__or2_0_52/B sky130_fd_sc_hd__inv_4_8/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__decap_12_1073 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_504 vssd1 vccd1 sky130_fd_sc_hd__inv_2_29/Y sky130_fd_sc_hd__nand2b_1_14/Y
+ sky130_fd_sc_hd__o21ai_1_504/B1 sky130_fd_sc_hd__xor2_1_304/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1084 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_515 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_7/X sky130_fd_sc_hd__o21ai_1_515/A1
+ sky130_fd_sc_hd__o21ai_1_515/B1 sky130_fd_sc_hd__xnor2_1_89/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1095 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_526 vssd1 vccd1 sky130_fd_sc_hd__inv_2_30/Y sky130_fd_sc_hd__nand2b_2_3/Y
+ sky130_fd_sc_hd__o21ai_1_526/B1 sky130_fd_sc_hd__xor2_1_325/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_537 vssd1 vccd1 sky130_fd_sc_hd__inv_2_28/Y sky130_fd_sc_hd__nand2b_1_8/Y
+ sky130_fd_sc_hd__o21ai_1_537/B1 sky130_fd_sc_hd__xor2_1_335/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_548 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_0/Y sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_548/B1 sky130_fd_sc_hd__xor2_1_347/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_559 vssd1 vccd1 sky130_fd_sc_hd__inv_2_31/Y sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_559/B1 sky130_fd_sc_hd__xor2_1_357/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_320 sky130_fd_sc_hd__fa_2_250/A sky130_fd_sc_hd__fa_2_221/B
+ sky130_fd_sc_hd__xor2_1_320/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_331 sky130_fd_sc_hd__dfxtp_2_5/Q sky130_fd_sc_hd__xor2_1_331/X
+ sky130_fd_sc_hd__xor2_1_331/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_342 sky130_fd_sc_hd__fa_2_250/A sky130_fd_sc_hd__fa_2_236/B
+ sky130_fd_sc_hd__xor2_1_342/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_353 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__xor2_1_353/X
+ sky130_fd_sc_hd__xor2_1_353/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_364 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__xor2_1_364/X
+ sky130_fd_sc_hd__xor2_1_364/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_375 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__xor2_1_375/X
+ sky130_fd_sc_hd__xor2_1_375/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_386 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__xor2_1_386/X
+ sky130_fd_sc_hd__xor2_1_386/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_397 sky130_fd_sc_hd__fa_2_281/A sky130_fd_sc_hd__fa_2_272/B
+ sky130_fd_sc_hd__xor2_1_397/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_302 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_302/X sky130_fd_sc_hd__clkbuf_1_302/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_313 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_313/X sky130_fd_sc_hd__clkinv_1_913/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_324 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_324/X sky130_fd_sc_hd__clkinv_1_981/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_335 vssd1 vccd1 sky130_fd_sc_hd__a22o_1_67/A2 sky130_fd_sc_hd__clkbuf_4_9/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_406 vccd1 vssd1 sky130_fd_sc_hd__and3_4_18/X sky130_fd_sc_hd__buf_6_4/X
+ sky130_fd_sc_hd__buf_6_0/X sky130_fd_sc_hd__nor2_2_32/Y sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__o21ai_1_674/B1 sky130_fd_sc_hd__nor2b_2_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_346 vssd1 vccd1 sky130_fd_sc_hd__inv_4_4/A sky130_fd_sc_hd__a222oi_1_10/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_417 vccd1 vssd1 sky130_fd_sc_hd__and3_4_25/X sky130_fd_sc_hd__buf_2_15/X
+ sky130_fd_sc_hd__buf_2_4/A sky130_fd_sc_hd__nor2_1_186/Y sky130_fd_sc_hd__buf_2_20/X
+ sky130_fd_sc_hd__o21ai_1_688/B1 sky130_fd_sc_hd__nor2b_1_17/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_357 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_4/B sky130_fd_sc_hd__or2_0_82/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_428 vccd1 vssd1 sky130_fd_sc_hd__and3_4_25/X sky130_fd_sc_hd__buf_2_24/X
+ sky130_fd_sc_hd__buf_2_27/X sky130_fd_sc_hd__nor2_1_186/Y sky130_fd_sc_hd__buf_2_15/X
+ sky130_fd_sc_hd__o21ai_1_702/B1 sky130_fd_sc_hd__nor2b_1_17/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_439 vccd1 vssd1 sky130_fd_sc_hd__and3_4_25/X sky130_fd_sc_hd__buf_2_26/X
+ sky130_fd_sc_hd__buf_2_24/X sky130_fd_sc_hd__nor2_1_186/Y sky130_fd_sc_hd__buf_2_27/X
+ sky130_fd_sc_hd__o21ai_1_716/B1 sky130_fd_sc_hd__nor2b_1_17/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__dfxtp_1_50 sky130_fd_sc_hd__nand2_1_64/B sky130_fd_sc_hd__dfxtp_1_51/CLK
+ sky130_fd_sc_hd__dfxtp_1_50/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_61 sky130_fd_sc_hd__nand2_1_55/B sky130_fd_sc_hd__dfxtp_1_62/CLK
+ sky130_fd_sc_hd__and2_0_13/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_72 sky130_fd_sc_hd__dfxtp_1_72/Q sky130_fd_sc_hd__dfxtp_1_72/CLK
+ sky130_fd_sc_hd__dfxtp_1_72/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_83 sky130_fd_sc_hd__dfxtp_1_83/Q sky130_fd_sc_hd__dfxtp_1_85/CLK
+ sky130_fd_sc_hd__dfxtp_1_83/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_94 sky130_fd_sc_hd__dfxtp_1_94/Q sky130_fd_sc_hd__dfxtp_1_94/CLK
+ sky130_fd_sc_hd__and2_0_3/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_300 vccd1 vssd1 sky130_fd_sc_hd__and2_0_300/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_21/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_311 vccd1 vssd1 sky130_fd_sc_hd__and2_0_311/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_311/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_322 vccd1 vssd1 sky130_fd_sc_hd__and2_0_322/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_322/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_333 vccd1 vssd1 sky130_fd_sc_hd__and2_0_333/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_333/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_344 vccd1 vssd1 sky130_fd_sc_hd__and2_0_344/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__buf_2_50/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_355 vccd1 vssd1 sky130_fd_sc_hd__and2_0_355/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__buf_2_48/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_366 vccd1 vssd1 sky130_fd_sc_hd__and2_0_366/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_71/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_377 vccd1 vssd1 sky130_fd_sc_hd__and2_0_377/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_67/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_388 vccd1 vssd1 sky130_fd_sc_hd__and2_0_388/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_72/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_399 vccd1 vssd1 sky130_fd_sc_hd__and2_0_399/X sky130_fd_sc_hd__and2_0_401/B
+ sky130_fd_sc_hd__and2_0_399/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__conb_1_8 sky130_fd_sc_hd__conb_1_8/LO sky130_fd_sc_hd__conb_1_8/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__inv_2_100 sky130_fd_sc_hd__inv_4_19/Y sky130_fd_sc_hd__inv_2_100/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_111 sky130_fd_sc_hd__inv_2_111/A sky130_fd_sc_hd__buf_12_7/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__or2_0_2 sky130_fd_sc_hd__or2_0_2/A sky130_fd_sc_hd__or2_0_2/X sky130_fd_sc_hd__or2_0_2/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__inv_2_122 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__inv_2_123/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_133 sky130_fd_sc_hd__inv_2_134/A sky130_fd_sc_hd__buf_8_41/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_144 sky130_fd_sc_hd__inv_2_144/A sky130_fd_sc_hd__inv_2_144/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_155 sky130_fd_sc_hd__inv_2_155/A sky130_fd_sc_hd__inv_2_155/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_166 sky130_fd_sc_hd__inv_2_166/A sky130_fd_sc_hd__buf_8_62/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_177 sky130_fd_sc_hd__inv_2_177/A sky130_fd_sc_hd__inv_2_177/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_188 sky130_fd_sc_hd__inv_2_188/A sky130_fd_sc_hd__inv_2_188/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_199 wbs_dat_i[9] sky130_fd_sc_hd__inv_2_199/Y vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__o22ai_1_107 sky130_fd_sc_hd__xnor2_2_6/Y sky130_fd_sc_hd__xnor2_1_256/Y
+ sky130_fd_sc_hd__fa_2_427/B sky130_fd_sc_hd__xnor2_1_263/Y sky130_fd_sc_hd__o22ai_1_98/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_118 sky130_fd_sc_hd__xnor2_1_273/Y sky130_fd_sc_hd__xnor2_1_264/Y
+ sky130_fd_sc_hd__fa_2_449/A sky130_fd_sc_hd__nor2b_1_19/A sky130_fd_sc_hd__o22ai_1_66/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_129 sky130_fd_sc_hd__xnor2_1_287/Y sky130_fd_sc_hd__xnor2_1_277/Y
+ sky130_fd_sc_hd__fa_2_458/A sky130_fd_sc_hd__nor2b_1_25/A sky130_fd_sc_hd__nand2_1_717/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_2_18 sky130_fd_sc_hd__buf_2_31/X sky130_fd_sc_hd__nor2_2_18/Y
+ sky130_fd_sc_hd__buf_2_19/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__nor2_2_29 sky130_fd_sc_hd__nor2_2_29/B sky130_fd_sc_hd__nor2_2_29/Y
+ sky130_fd_sc_hd__nor2_2_29/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__o211ai_1_8 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_8/A2
+ sky130_fd_sc_hd__o211ai_1_8/Y sky130_fd_sc_hd__a22oi_1_48/Y sky130_fd_sc_hd__a22oi_1_49/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__a211o_1_1 vssd1 vccd1 sky130_fd_sc_hd__a211o_1_1/X sky130_fd_sc_hd__dfxtp_1_64/Q
+ sky130_fd_sc_hd__nor2_1_5/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_1/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__o21ai_1_301 vssd1 vccd1 sky130_fd_sc_hd__buf_2_5/X sky130_fd_sc_hd__nand2b_1_1/Y
+ sky130_fd_sc_hd__o21ai_1_301/B1 sky130_fd_sc_hd__xor2_1_121/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_312 vssd1 vccd1 sky130_fd_sc_hd__inv_2_21/Y sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__o21ai_1_312/B1 sky130_fd_sc_hd__xor2_1_132/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_323 vssd1 vccd1 sky130_fd_sc_hd__inv_2_12/Y sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__o21ai_1_323/B1 sky130_fd_sc_hd__xor2_1_143/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_334 vssd1 vccd1 sky130_fd_sc_hd__inv_2_19/Y sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__o21ai_1_334/B1 sky130_fd_sc_hd__xor2_1_153/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_345 vssd1 vccd1 sky130_fd_sc_hd__buf_2_5/X sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__o21ai_1_345/B1 sky130_fd_sc_hd__xor2_1_162/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_356 vssd1 vccd1 sky130_fd_sc_hd__inv_2_11/Y sky130_fd_sc_hd__o21ai_1_356/A1
+ sky130_fd_sc_hd__o21ai_1_356/B1 sky130_fd_sc_hd__xnor2_1_47/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_367 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_187/B sky130_fd_sc_hd__nor2_1_97/Y
+ sky130_fd_sc_hd__nand2_1_286/Y sky130_fd_sc_hd__xnor2_1_50/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_378 vssd1 vccd1 sky130_fd_sc_hd__inv_2_15/Y sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__o21ai_1_378/B1 sky130_fd_sc_hd__xor2_1_193/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_389 vssd1 vccd1 sky130_fd_sc_hd__buf_2_3/X sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__o21ai_1_389/B1 sky130_fd_sc_hd__xor2_1_204/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nand2_1_705 sky130_fd_sc_hd__nand2_1_705/Y sky130_fd_sc_hd__buf_4_41/X
+ sky130_fd_sc_hd__xnor2_2_4/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_716 sky130_fd_sc_hd__o22ai_1_95/B2 sky130_fd_sc_hd__xnor2_2_5/Y
+ sky130_fd_sc_hd__xor2_1_669/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_14 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_14/A1 sky130_fd_sc_hd__buf_2_75/X
+ sky130_fd_sc_hd__mux2_8_0/S sky130_fd_sc_hd__or2_0_73/B vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_727 sky130_fd_sc_hd__nand2_1_727/Y sky130_fd_sc_hd__or2_0_86/X
+ sky130_fd_sc_hd__or2_0_87/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_25 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_25/A1 sky130_fd_sc_hd__buf_4_20/X
+ sky130_fd_sc_hd__mux2_8_1/S sky130_fd_sc_hd__or2_0_79/B vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_738 sky130_fd_sc_hd__nand2_1_738/Y sky130_fd_sc_hd__or2_0_90/A
+ sky130_fd_sc_hd__or2_0_90/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_36 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_36/A1 sky130_fd_sc_hd__buf_2_153/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__or2_1_11/A vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_749 sky130_fd_sc_hd__xnor2_1_211/B sky130_fd_sc_hd__nand2_1_750/Y
+ sky130_fd_sc_hd__or2_0_92/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_47 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_47/A1 sky130_fd_sc_hd__buf_2_149/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__mux2_2_47/X vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__conb_1_100 sky130_fd_sc_hd__conb_1_100/LO sky130_fd_sc_hd__conb_1_100/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_111 sky130_fd_sc_hd__conb_1_111/LO sky130_fd_sc_hd__conb_1_111/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_122 sky130_fd_sc_hd__conb_1_122/LO sky130_fd_sc_hd__conb_1_122/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_133 sky130_fd_sc_hd__conb_1_133/LO sky130_fd_sc_hd__clkinv_1_9/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_144 sky130_fd_sc_hd__conb_1_144/LO sky130_fd_sc_hd__conb_1_144/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__xor2_1_150 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__fa_2_111/A
+ sky130_fd_sc_hd__xor2_1_150/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_501 sky130_fd_sc_hd__ha_2_46/A sky130_fd_sc_hd__dfxtp_1_509/CLK
+ sky130_fd_sc_hd__and2_0_396/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_161 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__fa_2_117/B
+ sky130_fd_sc_hd__xor2_1_161/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1809 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_512 sky130_fd_sc_hd__xnor2_1_309/A sky130_fd_sc_hd__dfxtp_1_520/CLK
+ sky130_fd_sc_hd__and2_0_352/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_172 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__xor2_1_172/X
+ sky130_fd_sc_hd__xor2_1_172/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_523 wbs_dat_o[2] sky130_fd_sc_hd__dfxtp_1_533/CLK sky130_fd_sc_hd__nor2b_1_155/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_183 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__nor2_2_9/B
+ sky130_fd_sc_hd__xor2_1_183/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_534 wbs_dat_o[13] sky130_fd_sc_hd__dfxtp_1_538/CLK sky130_fd_sc_hd__nor2b_1_144/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_194 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__fa_2_135/B
+ sky130_fd_sc_hd__xor2_1_194/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_545 wbs_dat_o[24] sky130_fd_sc_hd__dfxtp_1_552/CLK sky130_fd_sc_hd__nor2b_1_133/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_110 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_110/X sky130_fd_sc_hd__clkbuf_1_110/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_121 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_121/X sky130_fd_sc_hd__inv_4_4/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_132 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_132/X sky130_fd_sc_hd__clkinv_2_0/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_203 vccd1 vssd1 sky130_fd_sc_hd__and3_4_2/X sky130_fd_sc_hd__or2_0_52/B
+ sky130_fd_sc_hd__or2_0_53/A sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__buf_2_32/X
+ sky130_fd_sc_hd__o21ai_1_375/B1 sky130_fd_sc_hd__and2b_4_4/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_143 vssd1 vccd1 sky130_fd_sc_hd__buf_8_16/A la_data_out[40]
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_214 vccd1 vssd1 sky130_fd_sc_hd__and3_4_10/X sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__buf_4_5/X sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__o21ai_1_402/B1 sky130_fd_sc_hd__and2b_4_7/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_154 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_11/A1 sky130_fd_sc_hd__clkbuf_1_154/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_1 sky130_fd_sc_hd__dfxtp_1_1/Q sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__dfxtp_1_1/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a222oi_1_225 vccd1 vssd1 sky130_fd_sc_hd__and3_4_13/X sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__buf_4_7/X sky130_fd_sc_hd__nor2_1_121/Y sky130_fd_sc_hd__nor2_2_5/A
+ sky130_fd_sc_hd__o21ai_1_416/B1 sky130_fd_sc_hd__nor2b_1_9/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_165 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_165/X sky130_fd_sc_hd__buf_2_184/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_236 vccd1 vssd1 sky130_fd_sc_hd__and3_4_13/X sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__buf_6_2/X sky130_fd_sc_hd__nor2_1_121/Y sky130_fd_sc_hd__buf_4_7/X
+ sky130_fd_sc_hd__o21ai_1_430/B1 sky130_fd_sc_hd__nor2b_1_9/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_176 vssd1 vccd1 sky130_fd_sc_hd__a22o_1_28/B2 sky130_fd_sc_hd__clkbuf_1_176/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_247 vccd1 vssd1 sky130_fd_sc_hd__and3_4_10/X sky130_fd_sc_hd__nor2_1_73/B
+ sky130_fd_sc_hd__buf_4_3/X sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__o21ai_1_445/B1 sky130_fd_sc_hd__and2b_4_7/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_187 vssd1 vccd1 sky130_fd_sc_hd__buf_8_50/A sky130_fd_sc_hd__conb_1_147/HI
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_258 vccd1 vssd1 sky130_fd_sc_hd__and3_4_16/X sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__buf_6_1/X sky130_fd_sc_hd__nor2_2_19/Y sky130_fd_sc_hd__and2_0_38/A
+ sky130_fd_sc_hd__o21ai_1_460/B1 sky130_fd_sc_hd__nor2b_2_3/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_198 vssd1 vccd1 sky130_fd_sc_hd__buf_8_134/A sky130_fd_sc_hd__buf_8_44/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_406 sky130_fd_sc_hd__fa_2_404/CIN sky130_fd_sc_hd__fa_2_407/B
+ sky130_fd_sc_hd__fa_2_406/A sky130_fd_sc_hd__fa_2_406/B sky130_fd_sc_hd__xor2_1_614/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o21ai_1_890 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_248/Y sky130_fd_sc_hd__xor2_1_666/B
+ sky130_fd_sc_hd__nand2_1_784/Y sky130_fd_sc_hd__xnor2_1_217/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_269 vccd1 vssd1 sky130_fd_sc_hd__and3_4_11/X sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__buf_4_2/X sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__o21ai_1_471/B1 sky130_fd_sc_hd__and2b_4_8/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__fa_2_417 sky130_fd_sc_hd__fa_2_416/CIN sky130_fd_sc_hd__fa_2_417/SUM
+ sky130_fd_sc_hd__fa_2_417/A sky130_fd_sc_hd__fa_2_417/B sky130_fd_sc_hd__fa_2_417/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_428 sky130_fd_sc_hd__fa_2_424/B sky130_fd_sc_hd__fa_2_430/CIN
+ sky130_fd_sc_hd__fa_2_428/A sky130_fd_sc_hd__fa_2_428/B sky130_fd_sc_hd__fa_2_428/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_439 sky130_fd_sc_hd__or2_0_93/A sky130_fd_sc_hd__nor2_1_251/B
+ sky130_fd_sc_hd__fa_2_439/A sky130_fd_sc_hd__fa_2_439/B sky130_fd_sc_hd__fa_2_442/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_4_11 sky130_fd_sc_hd__inv_4_11/Y sky130_fd_sc_hd__inv_4_11/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__and2_0_130 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_36/D sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_130/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_141 vccd1 vssd1 sky130_fd_sc_hd__and2_0_141/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_141/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_152 vccd1 vssd1 sky130_fd_sc_hd__and2_0_152/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_152/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_60 la_data_out[3] sky130_fd_sc_hd__conb_1_82/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_163 vccd1 vssd1 sky130_fd_sc_hd__and2_0_163/X sky130_fd_sc_hd__o21ai_2_0/B1
+ sky130_fd_sc_hd__and2_0_163/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_71 io_out[30] sky130_fd_sc_hd__conb_1_71/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_174 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_79/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_174/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_82 io_out[19] sky130_fd_sc_hd__conb_1_60/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_185 vccd1 vssd1 sky130_fd_sc_hd__and2_0_185/X sky130_fd_sc_hd__o21ai_2_0/B1
+ sky130_fd_sc_hd__and2_0_185/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_93 io_out[8] sky130_fd_sc_hd__conb_1_49/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_196 vccd1 vssd1 sky130_fd_sc_hd__and2_0_196/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_196/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__sdlclkp_1_2 sky130_fd_sc_hd__conb_1_143/LO sky130_fd_sc_hd__clkinv_8_4/Y
+ sky130_fd_sc_hd__clkinv_2_10/A sky130_fd_sc_hd__o21ai_2_4/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__sdlclkp_1
Xsky130_fd_sc_hd__o21ai_1_120 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_121/A2 sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__a22oi_1_170/Y sky130_fd_sc_hd__and2_0_153/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_131 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_133/A2 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_133/Y sky130_fd_sc_hd__and2_0_139/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_142 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_145/A2 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_138/Y sky130_fd_sc_hd__and2_0_125/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_153 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_153/A2 sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__a22oi_1_187/Y sky130_fd_sc_hd__and2_0_111/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_164 vssd1 vccd1 sky130_fd_sc_hd__a21oi_2_6/Y sky130_fd_sc_hd__nor2_2_3/Y
+ sky130_fd_sc_hd__nand2_1_237/Y sky130_fd_sc_hd__xnor2_1_32/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_175 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_241/A2 sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__a222oi_1_56/Y sky130_fd_sc_hd__xor2_1_8/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_186 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_186/A2 sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__a222oi_1_65/Y sky130_fd_sc_hd__xor2_1_17/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_197 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_237/A2 sky130_fd_sc_hd__nand2b_2_2/Y
+ sky130_fd_sc_hd__a222oi_1_73/Y sky130_fd_sc_hd__xor2_1_26/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_607 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_618 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_502 sky130_fd_sc_hd__nand2_1_502/Y sky130_fd_sc_hd__nor2_4_18/Y
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_629 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_513 sky130_fd_sc_hd__nand2_1_513/Y sky130_fd_sc_hd__nor2_1_166/Y
+ sky130_fd_sc_hd__nand2_1_546/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_524 sky130_fd_sc_hd__nand2_1_524/Y sky130_fd_sc_hd__nor2_1_170/Y
+ sky130_fd_sc_hd__nand2_1_546/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_535 sky130_fd_sc_hd__nand2_1_535/Y sky130_fd_sc_hd__nor2_1_175/Y
+ sky130_fd_sc_hd__nand2_1_546/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_546 sky130_fd_sc_hd__nand2_1_546/Y sky130_fd_sc_hd__or2_0_59/X
+ sky130_fd_sc_hd__nand2_1_546/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_557 sky130_fd_sc_hd__nand2_1_557/Y sky130_fd_sc_hd__or2_0_65/X
+ sky130_fd_sc_hd__nor2_1_182/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_568 sky130_fd_sc_hd__xnor2_1_155/A sky130_fd_sc_hd__nand2_1_569/Y
+ sky130_fd_sc_hd__or2_0_64/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_4 sky130_fd_sc_hd__and3_4_4/C sky130_fd_sc_hd__nor2b_1_4/Y
+ sky130_fd_sc_hd__and3_4_4/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nand2_1_579 sky130_fd_sc_hd__xor2_1_559/B sky130_fd_sc_hd__o21ai_2_15/B1
+ sky130_fd_sc_hd__nand2_1_579/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_1104 sky130_fd_sc_hd__clkinv_4_47/A sky130_fd_sc_hd__a22o_1_24/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1115 sky130_fd_sc_hd__clkinv_4_58/A sky130_fd_sc_hd__a22o_1_35/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1126 sky130_fd_sc_hd__clkinv_4_69/A sky130_fd_sc_hd__a22o_1_46/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1137 sky130_fd_sc_hd__buf_6_92/A sky130_fd_sc_hd__clkinv_4_81/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1148 sky130_fd_sc_hd__buf_2_44/A sky130_fd_sc_hd__inv_4_20/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1606 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1617 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_320 sky130_fd_sc_hd__or2_0_86/A sky130_fd_sc_hd__dfxtp_1_323/CLK
+ sky130_fd_sc_hd__and2_0_297/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1628 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_331 sky130_fd_sc_hd__dfxtp_1_331/Q sky130_fd_sc_hd__dfxtp_1_343/CLK
+ sky130_fd_sc_hd__and2_0_325/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1639 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_342 sky130_fd_sc_hd__dfxtp_1_342/Q sky130_fd_sc_hd__dfxtp_1_354/CLK
+ sky130_fd_sc_hd__and2_0_323/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_353 sky130_fd_sc_hd__dfxtp_1_353/Q sky130_fd_sc_hd__dfxtp_1_354/CLK
+ sky130_fd_sc_hd__and2_0_304/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_364 sky130_fd_sc_hd__dfxtp_1_364/Q sky130_fd_sc_hd__dfxtp_1_380/CLK
+ sky130_fd_sc_hd__nor2b_1_119/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_375 sky130_fd_sc_hd__dfxtp_1_375/Q sky130_fd_sc_hd__dfxtp_1_375/CLK
+ sky130_fd_sc_hd__nor2b_1_108/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_386 sky130_fd_sc_hd__dfxtp_1_386/Q sky130_fd_sc_hd__dfxtp_1_395/CLK
+ sky130_fd_sc_hd__nor2b_1_97/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_6 sky130_fd_sc_hd__nand2_1_6/Y sky130_fd_sc_hd__nand2_1_7/B
+ sky130_fd_sc_hd__or2_1_10/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_397 sky130_fd_sc_hd__dfxtp_1_397/Q sky130_fd_sc_hd__dfxtp_1_423/CLK
+ sky130_fd_sc_hd__nor2b_1_118/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_203 sky130_fd_sc_hd__fa_2_196/CIN sky130_fd_sc_hd__fa_2_202/A
+ sky130_fd_sc_hd__fa_2_203/A sky130_fd_sc_hd__fa_2_203/B sky130_fd_sc_hd__xor2_1_302/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_214 sky130_fd_sc_hd__fa_2_206/B sky130_fd_sc_hd__fa_2_211/A
+ sky130_fd_sc_hd__fa_2_214/A sky130_fd_sc_hd__fa_2_214/B sky130_fd_sc_hd__fa_2_214/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_225 sky130_fd_sc_hd__fa_2_219/A sky130_fd_sc_hd__fa_2_226/A
+ sky130_fd_sc_hd__fa_2_225/A sky130_fd_sc_hd__fa_2_225/B sky130_fd_sc_hd__xor2_1_323/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_236 sky130_fd_sc_hd__fa_2_230/A sky130_fd_sc_hd__fa_2_235/B
+ sky130_fd_sc_hd__fa_2_236/A sky130_fd_sc_hd__fa_2_236/B sky130_fd_sc_hd__fa_2_236/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_247 sky130_fd_sc_hd__fa_2_243/A sky130_fd_sc_hd__fah_1_4/B
+ sky130_fd_sc_hd__fa_2_247/A sky130_fd_sc_hd__fa_2_247/B sky130_fd_sc_hd__xor2_1_353/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_258 sky130_fd_sc_hd__fa_2_253/B sky130_fd_sc_hd__fa_2_256/A
+ sky130_fd_sc_hd__fa_2_258/A sky130_fd_sc_hd__fa_2_258/B sky130_fd_sc_hd__fa_2_258/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_269 sky130_fd_sc_hd__nor2_1_147/A sky130_fd_sc_hd__nor2_1_149/B
+ sky130_fd_sc_hd__fa_2_269/A sky130_fd_sc_hd__fa_2_269/B sky130_fd_sc_hd__fa_2_269/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_7 vccd1 vssd1 sky130_fd_sc_hd__and2_0_7/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_7/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__fa_2_50 sky130_fd_sc_hd__fa_2_42/A sky130_fd_sc_hd__fa_2_44/A sky130_fd_sc_hd__fa_2_50/A
+ sky130_fd_sc_hd__fa_2_50/B sky130_fd_sc_hd__xor2_1_71/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_61 sky130_fd_sc_hd__fa_2_54/CIN sky130_fd_sc_hd__fa_2_60/A
+ sky130_fd_sc_hd__fa_2_61/A sky130_fd_sc_hd__fa_2_61/B sky130_fd_sc_hd__xor2_1_89/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_72 sky130_fd_sc_hd__fa_2_64/B sky130_fd_sc_hd__fa_2_69/A sky130_fd_sc_hd__fa_2_72/A
+ sky130_fd_sc_hd__fa_2_72/B sky130_fd_sc_hd__fa_2_72/CIN vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_83 sky130_fd_sc_hd__fa_2_77/A sky130_fd_sc_hd__fa_2_84/A sky130_fd_sc_hd__fa_2_83/A
+ sky130_fd_sc_hd__fa_2_83/B sky130_fd_sc_hd__fa_2_83/CIN vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_94 sky130_fd_sc_hd__fa_2_88/A sky130_fd_sc_hd__fa_2_93/B sky130_fd_sc_hd__fa_2_94/A
+ sky130_fd_sc_hd__fa_2_94/B sky130_fd_sc_hd__fa_2_94/CIN vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a21oi_1_11 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_40/Y
+ sky130_fd_sc_hd__a21oi_1_11/Y sky130_fd_sc_hd__dfxtp_1_86/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_22 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_51/Y
+ sky130_fd_sc_hd__a21oi_1_22/Y sky130_fd_sc_hd__dfxtp_1_75/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_33 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_62/Y
+ sky130_fd_sc_hd__a21oi_1_33/Y sky130_fd_sc_hd__dfxtp_1_64/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_44 sky130_fd_sc_hd__a21oi_1_45/A1 sky130_fd_sc_hd__a21oi_1_44/B1
+ sky130_fd_sc_hd__a21oi_1_44/Y sky130_fd_sc_hd__nand2_1_197/B vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_208 sky130_fd_sc_hd__buf_6_65/X sky130_fd_sc_hd__buf_12_345/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_55 sky130_fd_sc_hd__xnor2_1_41/B sky130_fd_sc_hd__a21oi_1_55/B1
+ sky130_fd_sc_hd__xor2_1_154/A sky130_fd_sc_hd__nand2_1_259/A vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_219 sky130_fd_sc_hd__buf_4_28/X sky130_fd_sc_hd__buf_12_436/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_66 sky130_fd_sc_hd__xnor2_1_57/B sky130_fd_sc_hd__a21oi_1_66/B1
+ sky130_fd_sc_hd__xor2_1_199/A sky130_fd_sc_hd__or2_0_22/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_77 sky130_fd_sc_hd__a21oi_1_80/A1 sky130_fd_sc_hd__o21ai_1_456/Y
+ sky130_fd_sc_hd__a21oi_1_77/Y sky130_fd_sc_hd__nor2_1_115/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_88 sky130_fd_sc_hd__xnor2_1_104/B sky130_fd_sc_hd__o21ai_1_570/Y
+ sky130_fd_sc_hd__xor2_1_359/A sky130_fd_sc_hd__nor2_1_138/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_99 sky130_fd_sc_hd__or2_0_49/X sky130_fd_sc_hd__a21oi_1_99/B1
+ sky130_fd_sc_hd__a21oi_1_99/Y sky130_fd_sc_hd__a21oi_1_99/A2 vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__nor3_1_3 sky130_fd_sc_hd__nor3_1_3/C sky130_fd_sc_hd__nor3_1_3/Y
+ sky130_fd_sc_hd__nor3_1_3/A sky130_fd_sc_hd__nor3_1_3/B vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__clkinv_1_408 sky130_fd_sc_hd__nand2_1_277/A sky130_fd_sc_hd__nor2_1_92/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_419 sky130_fd_sc_hd__a21oi_1_74/A1 sky130_fd_sc_hd__nor2_1_111/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__bufinv_16_0 sky130_fd_sc_hd__bufinv_16_0/A sky130_fd_sc_hd__buf_12_484/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__bufinv_16
Xsky130_fd_sc_hd__decap_12_40 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_51 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_62 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_73 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_84 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_95 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_40 vccd1 vssd1 sky130_fd_sc_hd__buf_6_40/X sky130_fd_sc_hd__buf_8_76/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_51 vccd1 vssd1 sky130_fd_sc_hd__buf_6_51/X sky130_fd_sc_hd__buf_8_78/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_62 vccd1 vssd1 sky130_fd_sc_hd__buf_6_62/X sky130_fd_sc_hd__buf_8_82/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_73 vccd1 vssd1 sky130_fd_sc_hd__buf_6_73/X sky130_fd_sc_hd__buf_6_73/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_84 vccd1 vssd1 sky130_fd_sc_hd__buf_6_84/X sky130_fd_sc_hd__buf_6_84/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_20 sky130_fd_sc_hd__clkinv_4_62/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_31 sky130_fd_sc_hd__clkinv_4_76/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_42 sky130_fd_sc_hd__buf_2_193/A vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_53 sky130_fd_sc_hd__buf_2_192/A vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_64 sky130_fd_sc_hd__dfxtp_1_17/D vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a222oi_1_8 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_349/Q sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__o211ai_1_24/Y sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__a222oi_1_8/Y sky130_fd_sc_hd__dfxtp_1_300/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_404 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_415 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_426 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_310 sky130_fd_sc_hd__xnor2_1_3/B sky130_fd_sc_hd__nand2_1_311/Y
+ sky130_fd_sc_hd__nand2_1_310/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_437 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_321 sky130_fd_sc_hd__nand2_1_321/Y sky130_fd_sc_hd__or2_0_24/A
+ sky130_fd_sc_hd__or2_0_24/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_448 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_920 sky130_fd_sc_hd__clkinv_4_14/A sky130_fd_sc_hd__dfxtp_1_553/D
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_332 sky130_fd_sc_hd__nand2_1_332/Y sky130_fd_sc_hd__nor2_4_14/Y
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_459 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_931 sky130_fd_sc_hd__inv_2_121/A sky130_fd_sc_hd__clkinv_1_931/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_343 sky130_fd_sc_hd__nand2_1_343/Y sky130_fd_sc_hd__or2_0_9/A
+ sky130_fd_sc_hd__or2_0_9/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_942 sky130_fd_sc_hd__buf_2_156/A sky130_fd_sc_hd__inv_2_134/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_354 sky130_fd_sc_hd__nand2_1_354/Y sky130_fd_sc_hd__or2_0_58/A
+ sky130_fd_sc_hd__or2_0_39/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_953 sky130_fd_sc_hd__clkinv_1_954/A sky130_fd_sc_hd__nand2b_2_10/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_365 sky130_fd_sc_hd__nand2_1_365/Y sky130_fd_sc_hd__or2_0_61/A
+ sky130_fd_sc_hd__or2_0_42/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_964 sky130_fd_sc_hd__clkinv_1_964/Y sky130_fd_sc_hd__inv_2_152/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_376 sky130_fd_sc_hd__nand2_1_376/Y sky130_fd_sc_hd__or2_0_60/A
+ sky130_fd_sc_hd__or2_0_60/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_975 sky130_fd_sc_hd__clkinv_1_975/Y sky130_fd_sc_hd__clkinv_4_93/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_387 sky130_fd_sc_hd__nand2_1_387/Y sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__buf_4_5/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_986 sky130_fd_sc_hd__clkinv_1_986/Y sky130_fd_sc_hd__clkinv_4_29/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_398 sky130_fd_sc_hd__xor2_1_330/B sky130_fd_sc_hd__nand2_1_399/Y
+ sky130_fd_sc_hd__nand2_1_398/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_997 sky130_fd_sc_hd__clkinv_1_998/A sky130_fd_sc_hd__inv_4_5/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1403 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1414 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1425 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1436 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1447 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_150 sky130_fd_sc_hd__dfxtp_1_150/Q sky130_fd_sc_hd__dfxtp_1_152/CLK
+ sky130_fd_sc_hd__and2_0_221/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1458 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_161 sky130_fd_sc_hd__dfxtp_1_161/Q sky130_fd_sc_hd__dfxtp_1_176/CLK
+ sky130_fd_sc_hd__and2_0_111/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1469 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_172 sky130_fd_sc_hd__dfxtp_1_172/Q sky130_fd_sc_hd__dfxtp_1_177/CLK
+ sky130_fd_sc_hd__and2_0_166/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_183 sky130_fd_sc_hd__dfxtp_1_183/Q sky130_fd_sc_hd__clkinv_4_2/Y
+ sky130_fd_sc_hd__and2_0_222/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_194 sky130_fd_sc_hd__xor2_1_631/A sky130_fd_sc_hd__dfxtp_2_1/CLK
+ sky130_fd_sc_hd__and2_0_21/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_960 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_971 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_982 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_993 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o211ai_1_14 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_49/B1
+ sky130_fd_sc_hd__a22oi_1_2/A2 sky130_fd_sc_hd__a22oi_1_60/Y sky130_fd_sc_hd__a22oi_1_61/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_25 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_37/B1
+ sky130_fd_sc_hd__o211ai_1_25/Y sky130_fd_sc_hd__a22oi_1_82/Y sky130_fd_sc_hd__a22oi_1_83/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_36 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o21ai_1_6/A2
+ sky130_fd_sc_hd__fa_2_319/A sky130_fd_sc_hd__nand2_1_56/Y sky130_fd_sc_hd__a21oi_1_7/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_47 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o22ai_1_16/B1
+ sky130_fd_sc_hd__fa_2_383/A sky130_fd_sc_hd__nand2_1_67/Y sky130_fd_sc_hd__a21oi_1_18/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_58 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o22ai_1_5/B1
+ sky130_fd_sc_hd__fa_2_412/A sky130_fd_sc_hd__nand2_1_78/Y sky130_fd_sc_hd__a21oi_1_29/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__clkinv_1_205 sky130_fd_sc_hd__o22ai_1_50/B1 sky130_fd_sc_hd__dfxtp_1_172/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_216 sky130_fd_sc_hd__o22ai_1_10/B1 sky130_fd_sc_hd__dfxtp_1_105/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_227 sky130_fd_sc_hd__nor2_1_10/A sky130_fd_sc_hd__dfxtp_1_133/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_238 sky130_fd_sc_hd__o22ai_1_0/A2 sky130_fd_sc_hd__dfxtp_1_159/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_249 sky130_fd_sc_hd__o21ai_1_85/A2 sky130_fd_sc_hd__xor2_1_543/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_2_5 sky130_fd_sc_hd__o21ai_2_5/B1 sky130_fd_sc_hd__o21ai_2_5/Y
+ sky130_fd_sc_hd__xor2_1_42/A sky130_fd_sc_hd__nor2_1_52/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__o21ai_2
Xsky130_fd_sc_hd__and3_4_18 sky130_fd_sc_hd__nor2_2_32/B sky130_fd_sc_hd__nor2b_2_5/A
+ sky130_fd_sc_hd__nor2_2_32/A sky130_fd_sc_hd__and3_4_18/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__a21oi_1_102 sky130_fd_sc_hd__xnor2_1_123/A sky130_fd_sc_hd__clkinv_1_503/Y
+ sky130_fd_sc_hd__a21oi_1_102/Y sky130_fd_sc_hd__or2_0_48/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_113 sky130_fd_sc_hd__clkinv_1_549/Y sky130_fd_sc_hd__o21ai_1_711/Y
+ sky130_fd_sc_hd__a21oi_1_113/Y sky130_fd_sc_hd__nor2_1_175/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_124 sky130_fd_sc_hd__clkinv_1_580/Y sky130_fd_sc_hd__clkinv_1_579/Y
+ sky130_fd_sc_hd__a21oi_1_124/Y sky130_fd_sc_hd__nand2_1_605/A vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_135 sky130_fd_sc_hd__xnor2_1_182/B sky130_fd_sc_hd__clkinv_1_606/Y
+ sky130_fd_sc_hd__xor2_1_624/A sky130_fd_sc_hd__or2_0_68/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_146 sky130_fd_sc_hd__xnor2_1_196/B sky130_fd_sc_hd__clkinv_1_641/Y
+ sky130_fd_sc_hd__xor2_1_647/A sky130_fd_sc_hd__or2_0_80/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_157 sky130_fd_sc_hd__xnor2_1_210/A sky130_fd_sc_hd__clkinv_1_673/Y
+ sky130_fd_sc_hd__xor2_1_656/A sky130_fd_sc_hd__or2_0_91/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_168 sky130_fd_sc_hd__or2_0_97/X sky130_fd_sc_hd__clkinv_1_697/Y
+ sky130_fd_sc_hd__xor2_1_666/B sky130_fd_sc_hd__xnor2_1_218/A vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_179 sky130_fd_sc_hd__xnor2_1_300/B sky130_fd_sc_hd__clkinv_1_826/Y
+ sky130_fd_sc_hd__xor2_1_685/A sky130_fd_sc_hd__or2_0_109/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_109 sky130_fd_sc_hd__buf_8_109/A sky130_fd_sc_hd__buf_8_109/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_12_550 sky130_fd_sc_hd__buf_12_550/A sky130_fd_sc_hd__buf_12_550/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_561 sky130_fd_sc_hd__buf_12_561/A sky130_fd_sc_hd__buf_12_561/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_572 sky130_fd_sc_hd__buf_12_572/A sky130_fd_sc_hd__buf_12_572/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_201 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_583 sky130_fd_sc_hd__buf_12_583/A sky130_fd_sc_hd__buf_12_583/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_212 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_594 sky130_fd_sc_hd__buf_12_594/A sky130_fd_sc_hd__buf_12_594/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_223 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_234 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_245 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_256 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_140 sky130_fd_sc_hd__nand2_1_140/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__xnor2_1_123/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_267 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xnor2_1_302 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_302/B sky130_fd_sc_hd__xnor2_1_302/Y
+ sky130_fd_sc_hd__xnor2_1_302/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_151 sky130_fd_sc_hd__nor2_4_7/A sky130_fd_sc_hd__nor2_1_40/A
+ sky130_fd_sc_hd__ha_2_9/SUM vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_278 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_750 sky130_fd_sc_hd__fa_2_473/A sky130_fd_sc_hd__clkinv_1_750/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_162 sky130_fd_sc_hd__nand2_1_162/Y sky130_fd_sc_hd__nor2_4_10/Y
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_289 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_761 sky130_fd_sc_hd__fa_2_484/A sky130_fd_sc_hd__clkinv_1_761/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_173 sky130_fd_sc_hd__xor2_1_21/B sky130_fd_sc_hd__nand2_1_174/Y
+ sky130_fd_sc_hd__nand2_1_173/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_772 sky130_fd_sc_hd__xor2_1_675/B sky130_fd_sc_hd__clkinv_1_772/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_184 sky130_fd_sc_hd__xor2_1_42/B sky130_fd_sc_hd__o21ai_2_5/B1
+ sky130_fd_sc_hd__nand2_1_184/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_783 sky130_fd_sc_hd__and2_0_324/A sky130_fd_sc_hd__clkinv_1_783/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_195 sky130_fd_sc_hd__xor2_1_63/B sky130_fd_sc_hd__o21ai_2_6/B1
+ sky130_fd_sc_hd__nand2_1_195/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_794 sky130_fd_sc_hd__and2_0_313/A sky130_fd_sc_hd__clkinv_1_794/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1200 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_0 sky130_fd_sc_hd__xor2_1_0/B sky130_fd_sc_hd__xor2_2_0/A
+ sky130_fd_sc_hd__xor3_1_0/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1211 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1222 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1233 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1244 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1255 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1266 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1277 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_708 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_767/A2 sky130_fd_sc_hd__nand2b_2_7/Y
+ sky130_fd_sc_hd__o21ai_1_708/B1 sky130_fd_sc_hd__xor2_1_487/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1288 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_719 vssd1 vccd1 sky130_fd_sc_hd__inv_2_47/Y sky130_fd_sc_hd__nand2b_1_16/Y
+ sky130_fd_sc_hd__o21ai_1_719/B1 sky130_fd_sc_hd__xor2_1_496/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1299 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_15 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__fa_2_2/CIN
+ sky130_fd_sc_hd__xor2_1_15/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__and3_1_2 vssd1 vccd1 sky130_fd_sc_hd__and3_1_2/X sky130_fd_sc_hd__and3_1_2/B
+ sky130_fd_sc_hd__and3_1_2/A sky130_fd_sc_hd__and3_1_2/C vssd1 vccd1 sky130_fd_sc_hd__and3_1
Xsky130_fd_sc_hd__xor2_1_26 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__fa_2_10/A
+ sky130_fd_sc_hd__xor2_1_26/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_37 sky130_fd_sc_hd__fa_2_56/A sky130_fd_sc_hd__fa_2_22/B
+ sky130_fd_sc_hd__xor2_1_37/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_48 sky130_fd_sc_hd__fa_2_28/A sky130_fd_sc_hd__xor2_1_48/X
+ sky130_fd_sc_hd__xor2_1_48/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_59 sky130_fd_sc_hd__fa_2_75/A sky130_fd_sc_hd__fa_2_39/A
+ sky130_fd_sc_hd__xor2_1_59/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_790 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2b_1_9 sky130_fd_sc_hd__nand2b_1_9/Y sky130_fd_sc_hd__nor2_2_20/A
+ sky130_fd_sc_hd__nor2_2_20/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__xor2_1_502 sky130_fd_sc_hd__fa_2_357/A sky130_fd_sc_hd__fa_2_340/B
+ sky130_fd_sc_hd__xor2_1_502/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_513 sky130_fd_sc_hd__xor2_1_548/B sky130_fd_sc_hd__fa_2_347/B
+ sky130_fd_sc_hd__xor2_1_513/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_524 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__fa_2_353/B
+ sky130_fd_sc_hd__xor2_1_524/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_535 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__fa_2_356/A
+ sky130_fd_sc_hd__xor2_1_535/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_546 sky130_fd_sc_hd__or2_0_70/A sky130_fd_sc_hd__xor2_1_546/X
+ sky130_fd_sc_hd__xor2_1_546/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_557 sky130_fd_sc_hd__fa_2_379/A sky130_fd_sc_hd__and3_4_25/A
+ sky130_fd_sc_hd__xor2_1_557/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_568 sky130_fd_sc_hd__fa_2_389/A sky130_fd_sc_hd__fa_2_383/B
+ sky130_fd_sc_hd__xor2_1_568/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_579 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__fa_2_388/A
+ sky130_fd_sc_hd__xor2_1_579/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__ha_2_20 vssd1 vccd1 la_data_out[63] sky130_fd_sc_hd__ha_2_19/B sky130_fd_sc_hd__ha_2_20/SUM
+ sky130_fd_sc_hd__ha_2_20/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_31 vssd1 vccd1 la_data_out[41] sky130_fd_sc_hd__ha_2_30/B sky130_fd_sc_hd__ha_2_31/SUM
+ sky130_fd_sc_hd__ha_2_31/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_42 vssd1 vccd1 sky130_fd_sc_hd__ha_2_42/A sky130_fd_sc_hd__ha_2_41/B
+ sky130_fd_sc_hd__ha_2_42/SUM sky130_fd_sc_hd__ha_2_42/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__and2b_4_4 sky130_fd_sc_hd__nor2_4_9/A sky130_fd_sc_hd__and2b_4_4/X
+ sky130_fd_sc_hd__and3_4_2/C vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__and2b_4
Xsky130_fd_sc_hd__ha_2_53 vssd1 vccd1 sky130_fd_sc_hd__ha_2_53/A sky130_fd_sc_hd__ha_2_53/COUT
+ sky130_fd_sc_hd__ha_2_53/SUM sky130_fd_sc_hd__ha_2_53/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_5 vssd1 vccd1 sky130_fd_sc_hd__fa_2_262/A sky130_fd_sc_hd__xor2_1_383/B
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__nor2_1_140 sky130_fd_sc_hd__nor2_2_10/B sky130_fd_sc_hd__nor2_1_140/Y
+ sky130_fd_sc_hd__nor2_1_85/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_151 sky130_fd_sc_hd__nor2_1_152/Y sky130_fd_sc_hd__nor2_1_151/Y
+ sky130_fd_sc_hd__nor2_1_154/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_1_5 la_data_out[122] sky130_fd_sc_hd__clkinv_1_5/A vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_162 sky130_fd_sc_hd__xor2_1_420/X sky130_fd_sc_hd__nor2_1_162/Y
+ sky130_fd_sc_hd__a211o_1_2/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_173 sky130_fd_sc_hd__or2_0_61/B sky130_fd_sc_hd__nor2_1_173/Y
+ sky130_fd_sc_hd__or2_0_58/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_184 sky130_fd_sc_hd__nor2_1_187/Y sky130_fd_sc_hd__nor2_1_184/Y
+ sky130_fd_sc_hd__nor2_1_185/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_60 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__clkbuf_1_25/X
+ sky130_fd_sc_hd__nand2_1_69/B sky130_fd_sc_hd__dfxtp_1_141/Q sky130_fd_sc_hd__a22oi_1_60/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_71 sky130_fd_sc_hd__clkbuf_1_24/X sky130_fd_sc_hd__clkbuf_1_23/X
+ sky130_fd_sc_hd__dfxtp_1_114/Q sky130_fd_sc_hd__dfxtp_1_82/Q sky130_fd_sc_hd__a22oi_1_71/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_195 sky130_fd_sc_hd__nor2_2_30/Y sky130_fd_sc_hd__nor2_1_195/Y
+ sky130_fd_sc_hd__nor2_1_200/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_82 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__nor2_4_3/Y
+ sky130_fd_sc_hd__nand2_1_57/B sky130_fd_sc_hd__dfxtp_1_152/Q sky130_fd_sc_hd__a22oi_1_82/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_93 sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__dfxtp_1_125/Q sky130_fd_sc_hd__dfxtp_1_93/Q sky130_fd_sc_hd__a22oi_1_93/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_380 sky130_fd_sc_hd__buf_12_380/A sky130_fd_sc_hd__buf_12_577/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_391 sky130_fd_sc_hd__buf_12_391/A sky130_fd_sc_hd__buf_12_477/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xnor2_1_110 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_110/B sky130_fd_sc_hd__inv_2_30/A
+ sky130_fd_sc_hd__xnor2_1_110/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_121 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_121/B sky130_fd_sc_hd__inv_2_28/A
+ sky130_fd_sc_hd__xnor2_1_121/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__buf_8_19 sky130_fd_sc_hd__inv_2_73/Y sky130_fd_sc_hd__buf_8_19/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xnor2_1_132 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_132/B sky130_fd_sc_hd__buf_2_22/A
+ sky130_fd_sc_hd__xnor2_1_132/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_580 sky130_fd_sc_hd__clkinv_1_580/Y sky130_fd_sc_hd__a21oi_1_127/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_143 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_143/B sky130_fd_sc_hd__xnor2_1_143/Y
+ sky130_fd_sc_hd__xnor2_1_143/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_591 sky130_fd_sc_hd__xor2_1_597/A sky130_fd_sc_hd__o21ai_1_828/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_154 vssd1 vccd1 sky130_fd_sc_hd__o21ai_2_14/Y sky130_fd_sc_hd__xnor2_1_154/Y
+ sky130_fd_sc_hd__xnor2_1_154/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_165 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_165/B sky130_fd_sc_hd__inv_2_51/A
+ sky130_fd_sc_hd__xnor2_1_165/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_176 vssd1 vccd1 sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__nor2_4_16/A
+ sky130_fd_sc_hd__xnor2_1_176/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_187 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_636/X sky130_fd_sc_hd__xnor2_1_187/Y
+ sky130_fd_sc_hd__xnor2_1_187/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_198 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_198/B sky130_fd_sc_hd__and2_0_257/A
+ sky130_fd_sc_hd__xnor2_1_198/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_4_60 sky130_fd_sc_hd__clkinv_4_60/A sky130_fd_sc_hd__clkinv_4_60/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_71 sky130_fd_sc_hd__clkinv_4_71/A sky130_fd_sc_hd__clkinv_4_71/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_82 wbs_dat_i[24] sky130_fd_sc_hd__inv_2_95/A vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_93 sky130_fd_sc_hd__nand2_1_15/Y sky130_fd_sc_hd__clkinv_4_93/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_1030 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1041 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1052 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1063 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_1/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__decap_12_1074 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_505 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_505/A2 sky130_fd_sc_hd__or2b_2_1/X
+ sky130_fd_sc_hd__o21ai_1_505/B1 sky130_fd_sc_hd__xor2_1_305/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1085 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_516 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_535/B1 sky130_fd_sc_hd__nor2_1_126/A
+ sky130_fd_sc_hd__nor2_1_125/Y sky130_fd_sc_hd__o21ai_1_516/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1096 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_527 vssd1 vccd1 sky130_fd_sc_hd__inv_2_38/Y sky130_fd_sc_hd__nand2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_527/B1 sky130_fd_sc_hd__xor2_1_326/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_538 vssd1 vccd1 sky130_fd_sc_hd__nand2_2_12/Y sky130_fd_sc_hd__nand2b_1_14/Y
+ sky130_fd_sc_hd__a22oi_1_206/Y sky130_fd_sc_hd__xor2_1_336/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_549 vssd1 vccd1 sky130_fd_sc_hd__a21oi_1_92/Y sky130_fd_sc_hd__nor2_1_132/A
+ sky130_fd_sc_hd__a21oi_1_84/Y sky130_fd_sc_hd__o21ai_1_549/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_310 sky130_fd_sc_hd__fa_2_262/A sky130_fd_sc_hd__xor2_1_310/X
+ sky130_fd_sc_hd__xor2_1_310/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_321 sky130_fd_sc_hd__fa_2_262/A sky130_fd_sc_hd__fa_2_221/A
+ sky130_fd_sc_hd__xor2_1_321/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_332 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__fa_2_230/B
+ sky130_fd_sc_hd__xor2_1_332/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_343 sky130_fd_sc_hd__fa_2_239/A sky130_fd_sc_hd__xor2_1_343/X
+ sky130_fd_sc_hd__xor2_1_343/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_354 sky130_fd_sc_hd__fa_2_262/A sky130_fd_sc_hd__fa_2_247/B
+ sky130_fd_sc_hd__xor2_1_354/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_365 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__fa_2_249/B
+ sky130_fd_sc_hd__xor2_1_365/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_376 sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__fa_2_256/B
+ sky130_fd_sc_hd__xor2_1_376/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_387 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__fa_2_264/A
+ sky130_fd_sc_hd__xor2_1_387/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_398 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__fa_2_272/A
+ sky130_fd_sc_hd__xor2_1_398/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_303 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_303/X sky130_fd_sc_hd__buf_12_78/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_314 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_76/A sky130_fd_sc_hd__clkbuf_1_314/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_325 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_325/X sky130_fd_sc_hd__buf_8_21/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_336 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1_0/B_N sky130_fd_sc_hd__nor3b_1_1/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_407 vccd1 vssd1 sky130_fd_sc_hd__and3_4_24/X sky130_fd_sc_hd__buf_4_0/X
+ sky130_fd_sc_hd__buf_2_23/X sky130_fd_sc_hd__nor2_1_183/Y sky130_fd_sc_hd__buf_2_31/X
+ sky130_fd_sc_hd__o21ai_1_675/B1 sky130_fd_sc_hd__nor2b_1_16/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_347 vssd1 vccd1 sky130_fd_sc_hd__inv_4_3/A sky130_fd_sc_hd__a222oi_1_9/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_418 vccd1 vssd1 sky130_fd_sc_hd__and3_4_22/X sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__or2_0_60/B sky130_fd_sc_hd__nor2_4_18/Y sky130_fd_sc_hd__or2_0_60/A
+ sky130_fd_sc_hd__o21ai_1_689/B1 sky130_fd_sc_hd__and2b_4_10/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_358 vssd1 vccd1 sky130_fd_sc_hd__xnor2_2_5/B sky130_fd_sc_hd__or2_0_81/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_429 vccd1 vssd1 sky130_fd_sc_hd__and3_4_18/X sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__nor2_1_85/B sky130_fd_sc_hd__nor2_2_32/Y sky130_fd_sc_hd__nor2_2_10/B
+ sky130_fd_sc_hd__o21ai_1_703/B1 sky130_fd_sc_hd__nor2b_2_5/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__dfxtp_1_40 sky130_fd_sc_hd__nand2_1_74/B sky130_fd_sc_hd__dfxtp_1_45/CLK
+ sky130_fd_sc_hd__dfxtp_1_40/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_51 sky130_fd_sc_hd__nand2_1_63/B sky130_fd_sc_hd__dfxtp_1_51/CLK
+ sky130_fd_sc_hd__dfxtp_1_51/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_62 sky130_fd_sc_hd__nand2_1_59/B sky130_fd_sc_hd__dfxtp_1_62/CLK
+ sky130_fd_sc_hd__and2_0_2/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_73 sky130_fd_sc_hd__dfxtp_1_73/Q sky130_fd_sc_hd__dfxtp_1_81/CLK
+ sky130_fd_sc_hd__dfxtp_1_73/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_84 sky130_fd_sc_hd__dfxtp_1_84/Q sky130_fd_sc_hd__dfxtp_1_89/CLK
+ sky130_fd_sc_hd__dfxtp_1_84/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_95 sky130_fd_sc_hd__dfxtp_1_95/Q sky130_fd_sc_hd__dfxtp_1_97/CLK
+ sky130_fd_sc_hd__dfxtp_1_95/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_301 vccd1 vssd1 sky130_fd_sc_hd__a22o_1_6/B1 sky130_fd_sc_hd__and2_0_301/B
+ sky130_fd_sc_hd__or2_0_85/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_312 vccd1 vssd1 sky130_fd_sc_hd__and2_0_312/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_312/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_323 vccd1 vssd1 sky130_fd_sc_hd__and2_0_323/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_323/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_334 vccd1 vssd1 sky130_fd_sc_hd__and2_0_334/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_334/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_345 vccd1 vssd1 sky130_fd_sc_hd__and2_0_345/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__buf_2_40/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_356 vccd1 vssd1 sky130_fd_sc_hd__and2_0_356/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__and2_0_356/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_367 vccd1 vssd1 sky130_fd_sc_hd__and2_0_367/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_70/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_378 vccd1 vssd1 sky130_fd_sc_hd__and2_0_378/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_59/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_389 vccd1 vssd1 sky130_fd_sc_hd__and2_0_389/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_76/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__conb_1_9 sky130_fd_sc_hd__conb_1_9/LO sky130_fd_sc_hd__conb_1_9/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__inv_2_101 sky130_fd_sc_hd__inv_4_20/Y sky130_fd_sc_hd__inv_2_101/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_112 sky130_fd_sc_hd__inv_2_112/A sky130_fd_sc_hd__inv_2_112/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__or2_0_3 sky130_fd_sc_hd__or2_0_3/A sky130_fd_sc_hd__or2_0_3/X sky130_fd_sc_hd__or2_0_3/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__inv_2_123 sky130_fd_sc_hd__inv_2_123/A sky130_fd_sc_hd__buf_8_30/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_134 sky130_fd_sc_hd__inv_2_134/A sky130_fd_sc_hd__buf_8_46/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_145 sky130_fd_sc_hd__inv_2_145/A sky130_fd_sc_hd__inv_2_145/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_156 sky130_fd_sc_hd__inv_2_156/A sky130_fd_sc_hd__inv_2_156/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_167 sky130_fd_sc_hd__inv_2_167/A sky130_fd_sc_hd__buf_8_63/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_178 sky130_fd_sc_hd__inv_2_178/A sky130_fd_sc_hd__inv_2_178/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_189 sky130_fd_sc_hd__buf_6_24/A sky130_fd_sc_hd__inv_2_189/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__o22ai_1_108 sky130_fd_sc_hd__xnor2_2_5/Y sky130_fd_sc_hd__xnor2_1_257/Y
+ sky130_fd_sc_hd__fa_2_427/A sky130_fd_sc_hd__xnor2_1_265/Y sky130_fd_sc_hd__o22ai_1_95/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_119 sky130_fd_sc_hd__xnor2_2_5/Y sky130_fd_sc_hd__xnor2_1_265/Y
+ sky130_fd_sc_hd__fa_2_450/CIN sky130_fd_sc_hd__xnor2_1_266/Y sky130_fd_sc_hd__o22ai_1_95/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_2_19 sky130_fd_sc_hd__nor2_2_19/B sky130_fd_sc_hd__nor2_2_19/Y
+ sky130_fd_sc_hd__nor2_2_19/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__o211ai_1_9 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_9/A2
+ sky130_fd_sc_hd__o211ai_1_9/Y sky130_fd_sc_hd__a22oi_1_50/Y sky130_fd_sc_hd__a22oi_1_51/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__a211o_1_2 vssd1 vccd1 sky130_fd_sc_hd__a211o_1_2/X sky130_fd_sc_hd__dfxtp_1_65/Q
+ sky130_fd_sc_hd__nor2_1_6/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_2/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__o21ai_1_302 vssd1 vccd1 sky130_fd_sc_hd__inv_2_15/Y sky130_fd_sc_hd__nand2b_1_7/Y
+ sky130_fd_sc_hd__o21ai_1_302/B1 sky130_fd_sc_hd__xor2_1_122/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_313 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_0/Y sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__o21ai_1_313/B1 sky130_fd_sc_hd__xor2_1_134/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_324 vssd1 vccd1 sky130_fd_sc_hd__inv_2_17/Y sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__o21ai_1_324/B1 sky130_fd_sc_hd__xor2_1_144/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_335 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_80/Y sky130_fd_sc_hd__nand2_1_260/Y
+ sky130_fd_sc_hd__nand2_1_255/Y sky130_fd_sc_hd__o21ai_1_335/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_346 vssd1 vccd1 sky130_fd_sc_hd__inv_2_15/Y sky130_fd_sc_hd__nand2b_2_0/Y
+ sky130_fd_sc_hd__o21ai_1_346/B1 sky130_fd_sc_hd__xor2_1_163/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_357 vssd1 vccd1 sky130_fd_sc_hd__buf_2_2/X sky130_fd_sc_hd__nand2b_2_0/Y
+ sky130_fd_sc_hd__o21ai_1_357/B1 sky130_fd_sc_hd__xor2_1_173/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_368 vssd1 vccd1 sky130_fd_sc_hd__buf_2_3/X sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__o21ai_1_368/B1 sky130_fd_sc_hd__xor2_1_181/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_379 vssd1 vccd1 sky130_fd_sc_hd__nand2_4_4/Y sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__a22oi_1_199/Y sky130_fd_sc_hd__xor2_1_194/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nand2_1_706 sky130_fd_sc_hd__xnor2_1_199/A sky130_fd_sc_hd__nand2_1_707/Y
+ sky130_fd_sc_hd__or2_0_82/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_717 sky130_fd_sc_hd__nand2_1_717/Y sky130_fd_sc_hd__nor2b_1_25/A
+ sky130_fd_sc_hd__xor2_1_672/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_15 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_15/A1 sky130_fd_sc_hd__buf_2_76/X
+ sky130_fd_sc_hd__mux2_8_0/S sky130_fd_sc_hd__mux2_2_15/X vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_728 sky130_fd_sc_hd__xor2_1_653/B sky130_fd_sc_hd__nand2_1_729/Y
+ sky130_fd_sc_hd__or2_0_87/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_26 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_26/A1 sky130_fd_sc_hd__buf_2_154/X
+ sky130_fd_sc_hd__mux2_8_0/S sky130_fd_sc_hd__or2_1_11/B vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_739 sky130_fd_sc_hd__xnor2_1_208/A sky130_fd_sc_hd__nand2_1_740/Y
+ sky130_fd_sc_hd__or2_0_89/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_37 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_37/A1 sky130_fd_sc_hd__buf_2_96/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__mux2_2_37/X vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_48 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_48/A1 sky130_fd_sc_hd__buf_4_15/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__mux2_2_48/X vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__conb_1_101 sky130_fd_sc_hd__conb_1_101/LO sky130_fd_sc_hd__conb_1_101/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_112 sky130_fd_sc_hd__conb_1_112/LO sky130_fd_sc_hd__conb_1_112/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_123 sky130_fd_sc_hd__conb_1_123/LO sky130_fd_sc_hd__conb_1_123/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_134 sky130_fd_sc_hd__conb_1_134/LO sky130_fd_sc_hd__clkinv_1_8/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_145 sky130_fd_sc_hd__conb_1_145/LO sky130_fd_sc_hd__conb_1_145/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__xor2_1_140 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__xor2_1_140/X
+ sky130_fd_sc_hd__xor2_1_140/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_151 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__xor2_1_151/X
+ sky130_fd_sc_hd__xor2_1_151/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_502 sky130_fd_sc_hd__ha_2_45/A sky130_fd_sc_hd__dfxtp_1_509/CLK
+ sky130_fd_sc_hd__and2_0_395/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_162 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__xor2_1_162/X
+ sky130_fd_sc_hd__xor2_1_162/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_513 sky130_fd_sc_hd__ha_2_56/B sky130_fd_sc_hd__dfxtp_1_515/CLK
+ sky130_fd_sc_hd__and2_0_350/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_173 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__xor2_1_173/X
+ sky130_fd_sc_hd__xor2_1_173/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_524 wbs_dat_o[3] sky130_fd_sc_hd__dfxtp_1_532/CLK sky130_fd_sc_hd__nor2b_1_154/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_184 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__fa_2_132/B
+ sky130_fd_sc_hd__xor2_1_184/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_535 wbs_dat_o[14] sky130_fd_sc_hd__dfxtp_1_538/CLK sky130_fd_sc_hd__nor2b_1_143/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_195 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__fa_2_138/B
+ sky130_fd_sc_hd__xor2_1_195/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_546 wbs_dat_o[25] sky130_fd_sc_hd__dfxtp_1_552/CLK sky130_fd_sc_hd__nor2b_1_132/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_100 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_42/A1 sky130_fd_sc_hd__clkbuf_1_100/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_111 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_111/X sky130_fd_sc_hd__clkbuf_1_225/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_122 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_122/X sky130_fd_sc_hd__inv_4_3/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_133 vssd1 vccd1 sky130_fd_sc_hd__buf_12_61/A sky130_fd_sc_hd__buf_8_2/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_204 vccd1 vssd1 sky130_fd_sc_hd__and3_4_3/X sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__buf_4_6/X sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__buf_4_1/X
+ sky130_fd_sc_hd__o21ai_1_376/B1 sky130_fd_sc_hd__and2b_4_2/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_144 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_26/A1 sky130_fd_sc_hd__clkbuf_1_144/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_215 vccd1 vssd1 sky130_fd_sc_hd__and3_4_13/X sky130_fd_sc_hd__buf_4_7/X
+ sky130_fd_sc_hd__nor2_2_5/A sky130_fd_sc_hd__nor2_1_121/Y sky130_fd_sc_hd__nor2_2_5/B
+ sky130_fd_sc_hd__o21ai_1_403/B1 sky130_fd_sc_hd__nor2b_1_9/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_155 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_46/A1 sky130_fd_sc_hd__clkbuf_1_155/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_2 sky130_fd_sc_hd__dfxtp_1_2/Q sky130_fd_sc_hd__dfxtp_1_2/CLK
+ sky130_fd_sc_hd__dfxtp_1_2/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a222oi_1_226 vccd1 vssd1 sky130_fd_sc_hd__and3_4_14/X sky130_fd_sc_hd__buf_2_23/X
+ sky130_fd_sc_hd__buf_2_31/X sky130_fd_sc_hd__nor2_1_127/Y sky130_fd_sc_hd__buf_2_19/X
+ sky130_fd_sc_hd__o21ai_1_417/B1 sky130_fd_sc_hd__nor2b_1_10/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_166 vssd1 vccd1 sky130_fd_sc_hd__buf_8_23/A sky130_fd_sc_hd__inv_2_86/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_237 vccd1 vssd1 sky130_fd_sc_hd__and3_4_11/X sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__or2_0_66/A sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__or2_0_60/B
+ sky130_fd_sc_hd__o21ai_1_431/B1 sky130_fd_sc_hd__and2b_4_8/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_177 vssd1 vccd1 sky130_fd_sc_hd__a22o_1_27/B2 sky130_fd_sc_hd__clkbuf_1_177/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_248 vccd1 vssd1 sky130_fd_sc_hd__and3_4_14/X sky130_fd_sc_hd__buf_4_7/X
+ sky130_fd_sc_hd__buf_4_0/X sky130_fd_sc_hd__nor2_1_127/Y sky130_fd_sc_hd__buf_2_23/X
+ sky130_fd_sc_hd__o21ai_1_446/B1 sky130_fd_sc_hd__nor2b_1_10/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_188 vssd1 vccd1 sky130_fd_sc_hd__buf_12_21/A sky130_fd_sc_hd__buf_12_49/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o21ai_1_880 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_657/A sky130_fd_sc_hd__nor2_1_240/Y
+ sky130_fd_sc_hd__nand2_1_748/Y sky130_fd_sc_hd__xnor2_1_210/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_259 vccd1 vssd1 sky130_fd_sc_hd__and3_4_17/X sky130_fd_sc_hd__and2_0_49/A
+ sky130_fd_sc_hd__and2_0_45/A sky130_fd_sc_hd__nor2_2_20/Y sky130_fd_sc_hd__and2_0_87/A
+ sky130_fd_sc_hd__o21ai_1_461/B1 sky130_fd_sc_hd__nor2b_2_4/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_199 vssd1 vccd1 sky130_fd_sc_hd__buf_12_36/A sky130_fd_sc_hd__clkbuf_1_47/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_407 sky130_fd_sc_hd__nor2_1_206/A sky130_fd_sc_hd__nor2_1_209/B
+ sky130_fd_sc_hd__fa_2_407/A sky130_fd_sc_hd__fa_2_407/B sky130_fd_sc_hd__xor2_1_613/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o21ai_1_891 vssd1 vccd1 sky130_fd_sc_hd__inv_2_68/A sky130_fd_sc_hd__nand4_1_0/Y
+ sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__o21ai_1_891/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_418 sky130_fd_sc_hd__fa_2_417/CIN sky130_fd_sc_hd__fa_2_418/SUM
+ sky130_fd_sc_hd__fa_2_418/A sky130_fd_sc_hd__mux2_2_9/X sky130_fd_sc_hd__fa_2_418/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_429 sky130_fd_sc_hd__fa_2_421/CIN sky130_fd_sc_hd__fa_2_424/A
+ sky130_fd_sc_hd__fa_2_429/A sky130_fd_sc_hd__fa_2_429/B sky130_fd_sc_hd__fa_2_448/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_4_12 sky130_fd_sc_hd__inv_8_2/A sky130_fd_sc_hd__inv_4_12/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__and2_0_120 vccd1 vssd1 sky130_fd_sc_hd__and2_0_120/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_120/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_8_0 sky130_fd_sc_hd__nand2_8_0/A sky130_fd_sc_hd__nand2_8_0/B
+ sky130_fd_sc_hd__nor2_1_73/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_8
Xsky130_fd_sc_hd__and2_0_131 vccd1 vssd1 sky130_fd_sc_hd__and2_0_131/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_131/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_142 vccd1 vssd1 sky130_fd_sc_hd__and2_0_142/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_142/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_50 la_data_out[13] sky130_fd_sc_hd__conb_1_92/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_153 vccd1 vssd1 sky130_fd_sc_hd__and2_0_153/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_153/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_61 la_data_out[2] sky130_fd_sc_hd__conb_1_81/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_164 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_43/D sky130_fd_sc_hd__o21ai_2_0/B1
+ sky130_fd_sc_hd__and2_0_164/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_72 io_out[29] sky130_fd_sc_hd__conb_1_70/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_175 vccd1 vssd1 sky130_fd_sc_hd__and2_0_175/X sky130_fd_sc_hd__o21ai_2_0/B1
+ sky130_fd_sc_hd__and2_0_175/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_83 io_out[18] sky130_fd_sc_hd__conb_1_59/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_186 vccd1 vssd1 sky130_fd_sc_hd__and2_0_186/X sky130_fd_sc_hd__o21ai_2_0/B1
+ sky130_fd_sc_hd__and2_0_186/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_94 io_out[7] sky130_fd_sc_hd__conb_1_48/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_197 vccd1 vssd1 sky130_fd_sc_hd__and2_0_197/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_85/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__sdlclkp_1_3 sky130_fd_sc_hd__conb_1_145/LO sky130_fd_sc_hd__clkinv_8_7/Y
+ sky130_fd_sc_hd__clkinv_2_13/A sky130_fd_sc_hd__o21ai_1_891/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_1
Xsky130_fd_sc_hd__o21ai_1_110 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_113/A2 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_122/Y sky130_fd_sc_hd__and2_0_165/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_121 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_121/A2 sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__a22oi_1_171/Y sky130_fd_sc_hd__and2_0_152/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_132 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_133/A2 sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__a22oi_1_176/Y sky130_fd_sc_hd__and2_0_138/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_143 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_145/A2 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_139/Y sky130_fd_sc_hd__and2_0_124/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_154 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_157/A2 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_144/Y sky130_fd_sc_hd__and2_0_110/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_165 vssd1 vccd1 sky130_fd_sc_hd__inv_2_13/Y sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__o21ai_1_165/B1 sky130_fd_sc_hd__xor2_1_157/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_176 vssd1 vccd1 sky130_fd_sc_hd__inv_2_23/Y sky130_fd_sc_hd__nand2b_1_1/Y
+ sky130_fd_sc_hd__a222oi_1_57/Y sky130_fd_sc_hd__xor2_1_9/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_187 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_2/X sky130_fd_sc_hd__nand2_1_169/Y
+ sky130_fd_sc_hd__a21oi_1_38/Y sky130_fd_sc_hd__xnor2_1_7/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_198 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_295/A2 sky130_fd_sc_hd__nand2b_2_0/Y
+ sky130_fd_sc_hd__a222oi_1_74/Y sky130_fd_sc_hd__xor2_1_27/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_608 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_619 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_503 sky130_fd_sc_hd__nand2_1_503/Y sky130_fd_sc_hd__nand2_2_13/B
+ sky130_fd_sc_hd__nand2_1_657/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_514 sky130_fd_sc_hd__nor2_1_166/A sky130_fd_sc_hd__or2_0_57/X
+ sky130_fd_sc_hd__nand2_1_514/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_525 sky130_fd_sc_hd__xnor2_1_137/A sky130_fd_sc_hd__nand2_1_526/Y
+ sky130_fd_sc_hd__or2_0_58/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_536 sky130_fd_sc_hd__xnor2_1_142/A sky130_fd_sc_hd__nand2_1_537/Y
+ sky130_fd_sc_hd__or2_0_61/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_547 sky130_fd_sc_hd__xnor2_1_146/A sky130_fd_sc_hd__nand2_1_548/Y
+ sky130_fd_sc_hd__or2_0_60/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_558 sky130_fd_sc_hd__xnor2_1_150/A sky130_fd_sc_hd__nand2_1_559/Y
+ sky130_fd_sc_hd__or2_0_66/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_569 sky130_fd_sc_hd__nand2_1_569/Y sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__buf_4_4/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_5 sky130_fd_sc_hd__and3_4_5/C sky130_fd_sc_hd__nor2b_1_5/Y
+ sky130_fd_sc_hd__and3_4_5/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1105 sky130_fd_sc_hd__clkinv_4_48/A sky130_fd_sc_hd__a22o_1_25/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1116 sky130_fd_sc_hd__clkinv_4_59/A sky130_fd_sc_hd__a22o_1_36/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1127 sky130_fd_sc_hd__clkinv_4_70/A sky130_fd_sc_hd__a22o_1_47/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1138 sky130_fd_sc_hd__buf_4_38/A sky130_fd_sc_hd__clkinv_4_83/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1149 sky130_fd_sc_hd__and2_0_352/A sky130_fd_sc_hd__clkinv_4_88/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1607 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_310 sky130_fd_sc_hd__nor2_1_241/A sky130_fd_sc_hd__dfxtp_1_323/CLK
+ sky130_fd_sc_hd__and2_0_287/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1618 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_321 sky130_fd_sc_hd__or2_0_87/A sky130_fd_sc_hd__dfxtp_1_323/CLK
+ sky130_fd_sc_hd__and2_0_298/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1629 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_332 sky130_fd_sc_hd__dfxtp_1_332/Q sky130_fd_sc_hd__dfxtp_1_339/CLK
+ sky130_fd_sc_hd__and2_0_333/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_343 sky130_fd_sc_hd__dfxtp_1_343/Q sky130_fd_sc_hd__dfxtp_1_343/CLK
+ sky130_fd_sc_hd__and2_0_328/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_354 sky130_fd_sc_hd__dfxtp_1_354/Q sky130_fd_sc_hd__dfxtp_1_354/CLK
+ sky130_fd_sc_hd__and2_0_303/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_365 sky130_fd_sc_hd__dfxtp_1_365/Q sky130_fd_sc_hd__dfxtp_1_375/CLK
+ sky130_fd_sc_hd__nor2b_1_118/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_376 sky130_fd_sc_hd__dfxtp_1_376/Q sky130_fd_sc_hd__dfxtp_1_380/CLK
+ sky130_fd_sc_hd__nor2b_1_107/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_387 sky130_fd_sc_hd__dfxtp_1_387/Q sky130_fd_sc_hd__dfxtp_1_395/CLK
+ sky130_fd_sc_hd__nor2b_1_96/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_7 sky130_fd_sc_hd__nand2_8_4/A sky130_fd_sc_hd__nand2_1_7/B
+ sky130_fd_sc_hd__or2_0_80/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_398 sky130_fd_sc_hd__dfxtp_1_398/Q sky130_fd_sc_hd__clkinv_4_8/Y
+ sky130_fd_sc_hd__nor2b_1_117/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_204 sky130_fd_sc_hd__fa_2_197/A sky130_fd_sc_hd__fa_2_205/A
+ sky130_fd_sc_hd__fa_2_204/A sky130_fd_sc_hd__fa_2_204/B sky130_fd_sc_hd__xor2_1_297/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_215 sky130_fd_sc_hd__nor2_2_12/A sky130_fd_sc_hd__or2_0_33/B
+ sky130_fd_sc_hd__fa_2_215/A sky130_fd_sc_hd__fa_2_215/B sky130_fd_sc_hd__fa_2_215/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_226 sky130_fd_sc_hd__fa_2_222/B sky130_fd_sc_hd__fa_2_228/CIN
+ sky130_fd_sc_hd__fa_2_226/A sky130_fd_sc_hd__fa_2_226/B sky130_fd_sc_hd__fa_2_226/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_237 sky130_fd_sc_hd__fa_2_231/A sky130_fd_sc_hd__fa_2_238/B
+ sky130_fd_sc_hd__fa_2_237/A sky130_fd_sc_hd__fa_2_237/B sky130_fd_sc_hd__xor2_1_338/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_248 sky130_fd_sc_hd__fa_2_245/A sky130_fd_sc_hd__fah_1_3/A
+ sky130_fd_sc_hd__fa_2_248/A sky130_fd_sc_hd__fa_2_248/B sky130_fd_sc_hd__xor2_1_357/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_259 sky130_fd_sc_hd__nor2_1_139/A sky130_fd_sc_hd__nor2_1_142/B
+ sky130_fd_sc_hd__fa_2_259/A sky130_fd_sc_hd__fa_2_259/B sky130_fd_sc_hd__fa_2_259/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_40 sky130_fd_sc_hd__fa_2_33/A sky130_fd_sc_hd__fa_2_41/B sky130_fd_sc_hd__fa_2_40/A
+ sky130_fd_sc_hd__fa_2_40/B sky130_fd_sc_hd__fa_2_40/CIN vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_8 vccd1 vssd1 sky130_fd_sc_hd__and2_0_8/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_8/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__fa_2_51 sky130_fd_sc_hd__or2_0_2/A sky130_fd_sc_hd__nor2_1_58/B
+ sky130_fd_sc_hd__fa_2_51/A sky130_fd_sc_hd__fa_2_51/B sky130_fd_sc_hd__fa_2_51/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_62 sky130_fd_sc_hd__fa_2_55/A sky130_fd_sc_hd__fa_2_63/A sky130_fd_sc_hd__fa_2_62/A
+ sky130_fd_sc_hd__fa_2_62/B sky130_fd_sc_hd__xor2_1_84/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_73 sky130_fd_sc_hd__nor2_1_62/A sky130_fd_sc_hd__or2_0_6/B
+ sky130_fd_sc_hd__fa_2_73/A sky130_fd_sc_hd__fa_2_73/B sky130_fd_sc_hd__fa_2_73/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_84 sky130_fd_sc_hd__fa_2_80/B sky130_fd_sc_hd__fa_2_86/CIN
+ sky130_fd_sc_hd__fa_2_84/A sky130_fd_sc_hd__fa_2_84/B sky130_fd_sc_hd__fa_2_84/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_95 sky130_fd_sc_hd__fa_2_89/A sky130_fd_sc_hd__fa_2_96/B sky130_fd_sc_hd__fa_2_95/A
+ sky130_fd_sc_hd__fa_2_95/B sky130_fd_sc_hd__fa_2_95/CIN vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_210 vccd1 vssd1 la_data_out[80] sky130_fd_sc_hd__xnor2_2_4/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__a21oi_1_12 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_41/Y
+ sky130_fd_sc_hd__a21oi_1_12/Y sky130_fd_sc_hd__dfxtp_1_85/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_23 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_52/Y
+ sky130_fd_sc_hd__a21oi_1_23/Y sky130_fd_sc_hd__dfxtp_1_74/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_34 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_63/Y
+ sky130_fd_sc_hd__a21oi_1_34/Y sky130_fd_sc_hd__dfxtp_1_65/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_45 sky130_fd_sc_hd__a21oi_1_45/A1 sky130_fd_sc_hd__nor2_1_59/A
+ sky130_fd_sc_hd__a21oi_1_45/Y sky130_fd_sc_hd__or2_0_13/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_209 sky130_fd_sc_hd__buf_6_57/X sky130_fd_sc_hd__buf_12_406/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a222oi_1_590 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_396/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_428/Q sky130_fd_sc_hd__clkbuf_1_32/X
+ sky130_fd_sc_hd__clkinv_1_787/A sky130_fd_sc_hd__dfxtp_1_364/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a21oi_1_56 sky130_fd_sc_hd__o21ai_1_360/Y sky130_fd_sc_hd__o21ai_1_341/Y
+ sky130_fd_sc_hd__o21ai_2_7/A2 sky130_fd_sc_hd__nor2_1_82/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_67 sky130_fd_sc_hd__xnor2_1_60/A sky130_fd_sc_hd__a21oi_1_67/B1
+ sky130_fd_sc_hd__a21oi_1_67/Y sky130_fd_sc_hd__or2_0_21/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_78 sky130_fd_sc_hd__a21oi_1_80/A1 sky130_fd_sc_hd__o21ai_1_474/Y
+ sky130_fd_sc_hd__a21oi_1_78/Y sky130_fd_sc_hd__nor2_1_118/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_89 sky130_fd_sc_hd__a21oi_1_89/A1 sky130_fd_sc_hd__a21oi_1_89/B1
+ sky130_fd_sc_hd__a21oi_1_89/Y sky130_fd_sc_hd__nand2_1_434/A vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__nor3_1_4 sky130_fd_sc_hd__nor4_1_1/D sky130_fd_sc_hd__nor3_1_4/Y
+ wbs_ack_o wbs_we_i vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__clkinv_1_409 sky130_fd_sc_hd__nand2_1_252/A sky130_fd_sc_hd__nor2_2_10/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__bufinv_16_1 sky130_fd_sc_hd__bufinv_16_1/A sky130_fd_sc_hd__buf_12_269/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__bufinv_16
Xsky130_fd_sc_hd__decap_12_30 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_41 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_52 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_63 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_74 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_85 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_96 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_30 vccd1 vssd1 sky130_fd_sc_hd__buf_6_30/X sky130_fd_sc_hd__buf_8_99/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_41 vccd1 vssd1 sky130_fd_sc_hd__buf_6_41/X sky130_fd_sc_hd__buf_8_65/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_52 vccd1 vssd1 sky130_fd_sc_hd__buf_6_52/X sky130_fd_sc_hd__buf_8_6/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_63 vccd1 vssd1 sky130_fd_sc_hd__buf_6_63/X sky130_fd_sc_hd__buf_8_87/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_74 vccd1 vssd1 sky130_fd_sc_hd__buf_6_74/X sky130_fd_sc_hd__buf_6_74/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_85 vccd1 vssd1 sky130_fd_sc_hd__buf_6_85/X sky130_fd_sc_hd__buf_8_10/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_10 sky130_fd_sc_hd__conb_1_147/HI vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_21 sky130_fd_sc_hd__clkinv_4_64/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_32 sky130_fd_sc_hd__clkinv_4_75/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_43 sky130_fd_sc_hd__buf_2_189/A vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_54 sky130_fd_sc_hd__buf_2_192/A vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_65 sky130_fd_sc_hd__dfxtp_1_3/D vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a222oi_1_9 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_350/Q sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__a22oi_1_8/B1 sky130_fd_sc_hd__o211ai_1_25/Y sky130_fd_sc_hd__a22oi_1_8/A1
+ sky130_fd_sc_hd__a222oi_1_9/Y sky130_fd_sc_hd__dfxtp_1_301/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__decap_12_405 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_416 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_300 sky130_fd_sc_hd__nand2_1_300/Y sky130_fd_sc_hd__or2_0_23/A
+ sky130_fd_sc_hd__or2_0_23/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_427 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_311 sky130_fd_sc_hd__nand2_1_311/Y sky130_fd_sc_hd__buf_8_0/X
+ sky130_fd_sc_hd__inv_6_0/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_438 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_910 sky130_fd_sc_hd__clkinv_1_910/Y sky130_fd_sc_hd__inv_2_105/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_322 sky130_fd_sc_hd__nand2_1_322/Y sky130_fd_sc_hd__nor2_1_109/Y
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_449 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_921 sky130_fd_sc_hd__clkinv_4_15/A sky130_fd_sc_hd__nand2_2_14/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_333 sky130_fd_sc_hd__xnor2_1_67/B sky130_fd_sc_hd__or2_0_53/A
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_932 sky130_fd_sc_hd__inv_8_0/A sky130_fd_sc_hd__a21o_2_2/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_344 sky130_fd_sc_hd__xor2_1_234/B sky130_fd_sc_hd__nand2_1_345/Y
+ sky130_fd_sc_hd__nand2_1_344/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_943 sky130_fd_sc_hd__inv_2_135/A sky130_fd_sc_hd__buf_8_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_355 sky130_fd_sc_hd__xor2_1_255/B sky130_fd_sc_hd__o21ai_2_11/B1
+ sky130_fd_sc_hd__nand2_1_355/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_954 sky130_fd_sc_hd__clkinv_1_954/Y sky130_fd_sc_hd__clkinv_1_954/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_366 sky130_fd_sc_hd__xor2_1_276/B sky130_fd_sc_hd__nand2_1_367/Y
+ sky130_fd_sc_hd__nand2_1_366/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_965 sky130_fd_sc_hd__clkinv_1_965/Y sky130_fd_sc_hd__inv_2_152/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_377 sky130_fd_sc_hd__xor2_1_296/B sky130_fd_sc_hd__nand2_1_378/Y
+ sky130_fd_sc_hd__nand2_1_377/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_976 sky130_fd_sc_hd__clkinv_1_976/Y sky130_fd_sc_hd__clkinv_4_94/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_388 sky130_fd_sc_hd__xor2_1_313/B sky130_fd_sc_hd__nand2_1_389/Y
+ sky130_fd_sc_hd__nand2_1_388/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_987 sky130_fd_sc_hd__clkinv_1_987/Y sky130_fd_sc_hd__clkinv_4_31/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_399 sky130_fd_sc_hd__nand2_1_399/Y sky130_fd_sc_hd__nor2_2_15/A
+ sky130_fd_sc_hd__nor2_2_15/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_998 sky130_fd_sc_hd__clkinv_1_998/Y sky130_fd_sc_hd__clkinv_1_998/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1404 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1415 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1426 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1437 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_140 sky130_fd_sc_hd__dfxtp_1_140/Q sky130_fd_sc_hd__dfxtp_1_141/CLK
+ sky130_fd_sc_hd__and2_0_175/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1448 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_151 sky130_fd_sc_hd__dfxtp_1_151/Q sky130_fd_sc_hd__dfxtp_1_154/CLK
+ sky130_fd_sc_hd__and2_0_226/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1459 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_162 sky130_fd_sc_hd__dfxtp_1_162/Q sky130_fd_sc_hd__dfxtp_1_176/CLK
+ sky130_fd_sc_hd__and2_0_119/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_173 sky130_fd_sc_hd__dfxtp_1_173/Q sky130_fd_sc_hd__dfxtp_1_177/CLK
+ sky130_fd_sc_hd__and2_0_178/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_184 sky130_fd_sc_hd__dfxtp_1_184/Q sky130_fd_sc_hd__clkinv_4_2/Y
+ sky130_fd_sc_hd__and2_0_227/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_195 sky130_fd_sc_hd__xnor2_1_180/A sky130_fd_sc_hd__dfxtp_2_1/CLK
+ sky130_fd_sc_hd__and2_0_24/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_950 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_961 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_972 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_983 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_994 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o211ai_1_15 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_48/B1
+ sky130_fd_sc_hd__a22oi_1_0/A2 sky130_fd_sc_hd__a22oi_1_62/Y sky130_fd_sc_hd__a22oi_1_63/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_26 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_36/B1
+ sky130_fd_sc_hd__o211ai_1_26/Y sky130_fd_sc_hd__a22oi_1_84/Y sky130_fd_sc_hd__a22oi_1_85/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_37 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o21ai_1_7/A2
+ sky130_fd_sc_hd__fa_2_327/A sky130_fd_sc_hd__nand2_1_57/Y sky130_fd_sc_hd__a21oi_1_8/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_48 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o22ai_1_15/B1
+ sky130_fd_sc_hd__fa_2_389/B sky130_fd_sc_hd__nand2_1_68/Y sky130_fd_sc_hd__a21oi_1_19/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_59 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o22ai_1_4/B1
+ sky130_fd_sc_hd__fa_2_413/A sky130_fd_sc_hd__nand2_1_79/Y sky130_fd_sc_hd__a21oi_1_30/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__clkinv_1_206 sky130_fd_sc_hd__nor2_1_17/A sky130_fd_sc_hd__dfxtp_1_140/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_217 sky130_fd_sc_hd__o22ai_1_9/A2 sky130_fd_sc_hd__dfxtp_1_168/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_228 sky130_fd_sc_hd__o22ai_1_6/B1 sky130_fd_sc_hd__dfxtp_1_101/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_239 sky130_fd_sc_hd__nor2_1_4/A sky130_fd_sc_hd__dfxtp_1_127/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_2_6 sky130_fd_sc_hd__o21ai_2_6/B1 sky130_fd_sc_hd__o21ai_2_6/Y
+ sky130_fd_sc_hd__xor2_1_63/A sky130_fd_sc_hd__nor2_1_58/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__o21ai_2
Xsky130_fd_sc_hd__and3_4_19 sky130_fd_sc_hd__and3_4_19/A sky130_fd_sc_hd__nor2_4_15/B
+ sky130_fd_sc_hd__or2b_2_2/A sky130_fd_sc_hd__and3_4_19/X vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__and3_4
Xsky130_fd_sc_hd__a21oi_1_103 sky130_fd_sc_hd__xor2_1_423/X sky130_fd_sc_hd__clkinv_1_508/Y
+ sky130_fd_sc_hd__o21a_1_3/A1 sky130_fd_sc_hd__or2_0_51/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_114 sky130_fd_sc_hd__clkinv_1_549/Y sky130_fd_sc_hd__clkinv_1_542/Y
+ sky130_fd_sc_hd__a21oi_1_114/Y sky130_fd_sc_hd__nand2_1_540/B vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_125 sky130_fd_sc_hd__xnor2_1_166/B sky130_fd_sc_hd__clkinv_1_513/Y
+ sky130_fd_sc_hd__xor2_1_580/A sky130_fd_sc_hd__nand2_1_602/A vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_136 sky130_fd_sc_hd__xnor2_1_185/A sky130_fd_sc_hd__clkinv_1_608/Y
+ sky130_fd_sc_hd__a21oi_1_136/Y sky130_fd_sc_hd__or2_0_67/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_147 sky130_fd_sc_hd__xnor2_1_197/B sky130_fd_sc_hd__clkinv_1_643/Y
+ sky130_fd_sc_hd__xor2_1_648/A sky130_fd_sc_hd__or2_1_10/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_158 sky130_fd_sc_hd__or2_0_92/X sky130_fd_sc_hd__clkinv_1_675/Y
+ sky130_fd_sc_hd__xor2_1_657/A sky130_fd_sc_hd__xnor2_1_211/A vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_169 sky130_fd_sc_hd__xnor2_1_290/B sky130_fd_sc_hd__clkinv_1_806/Y
+ sky130_fd_sc_hd__a21oi_1_169/Y sky130_fd_sc_hd__or2_0_99/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_540 sky130_fd_sc_hd__buf_12_540/A sky130_fd_sc_hd__buf_12_540/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_551 sky130_fd_sc_hd__buf_12_551/A sky130_fd_sc_hd__buf_12_551/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_562 sky130_fd_sc_hd__buf_12_562/A sky130_fd_sc_hd__buf_12_562/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_573 sky130_fd_sc_hd__buf_12_573/A sky130_fd_sc_hd__buf_12_573/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_202 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_584 sky130_fd_sc_hd__buf_12_584/A sky130_fd_sc_hd__buf_12_584/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_213 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_595 sky130_fd_sc_hd__buf_12_595/A sky130_fd_sc_hd__buf_12_595/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_224 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_235 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_246 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_130 sky130_fd_sc_hd__nand2_1_130/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_131/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_257 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_141 sky130_fd_sc_hd__nand2_1_141/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__xnor2_1_123/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_268 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_740 sky130_fd_sc_hd__nor2b_1_119/A sky130_fd_sc_hd__xnor2_1_303/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_303 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_303/B sky130_fd_sc_hd__xnor2_1_303/Y
+ sky130_fd_sc_hd__nor2b_1_85/Y vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_152 sky130_fd_sc_hd__nand2_1_152/Y sky130_fd_sc_hd__nor2_1_48/Y
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_279 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_751 sky130_fd_sc_hd__fa_2_474/A sky130_fd_sc_hd__clkinv_1_751/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_163 sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__nor2_1_46/Y
+ sky130_fd_sc_hd__nor2_1_54/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_762 sky130_fd_sc_hd__fa_2_485/A sky130_fd_sc_hd__clkinv_1_762/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_174 sky130_fd_sc_hd__nand2_1_174/Y sky130_fd_sc_hd__nor2_2_2/A
+ sky130_fd_sc_hd__nor2_2_2/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_773 sky130_fd_sc_hd__and2_0_334/A sky130_fd_sc_hd__clkinv_1_773/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_185 sky130_fd_sc_hd__o21ai_2_5/B1 sky130_fd_sc_hd__nor2_1_52/A
+ sky130_fd_sc_hd__nor2_1_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_784 sky130_fd_sc_hd__and2_0_323/A sky130_fd_sc_hd__clkinv_1_784/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_196 sky130_fd_sc_hd__o21ai_2_6/B1 sky130_fd_sc_hd__nor2_1_58/A
+ sky130_fd_sc_hd__nor2_1_58/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_795 sky130_fd_sc_hd__and2_0_312/A sky130_fd_sc_hd__clkinv_1_795/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1201 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_1 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__xor3_1_3/C
+ sky130_fd_sc_hd__xor2_1_1/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1212 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1223 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1234 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1245 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1256 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1267 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1278 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_709 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_709/A2 sky130_fd_sc_hd__or2b_2_2/X
+ sky130_fd_sc_hd__o21ai_1_709/B1 sky130_fd_sc_hd__xor2_1_488/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1289 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_16 sky130_fd_sc_hd__xor2_1_9/B sky130_fd_sc_hd__fa_2_2/B
+ sky130_fd_sc_hd__xor2_1_16/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_27 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__xor2_1_27/X
+ sky130_fd_sc_hd__xor2_1_27/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_38 sky130_fd_sc_hd__fa_2_28/A sky130_fd_sc_hd__fa_2_19/B
+ sky130_fd_sc_hd__xor2_1_38/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_49 sky130_fd_sc_hd__fa_2_28/A sky130_fd_sc_hd__and3_1_0/B
+ sky130_fd_sc_hd__xor2_1_49/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_780 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_791 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_503 sky130_fd_sc_hd__fa_2_338/A sky130_fd_sc_hd__xor2_1_503/X
+ sky130_fd_sc_hd__xor2_1_503/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_514 sky130_fd_sc_hd__fah_1_15/A sky130_fd_sc_hd__fa_2_347/A
+ sky130_fd_sc_hd__xor2_1_514/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_525 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__fa_2_349/A
+ sky130_fd_sc_hd__xor2_1_525/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_536 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__xor2_1_536/X
+ sky130_fd_sc_hd__xor2_1_536/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_547 sky130_fd_sc_hd__fah_1_14/A sky130_fd_sc_hd__xor2_1_547/X
+ sky130_fd_sc_hd__xor2_1_547/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_558 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__fa_2_375/A
+ sky130_fd_sc_hd__xor2_1_558/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_569 sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__fa_2_385/A
+ sky130_fd_sc_hd__xor2_1_569/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1790 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__ha_2_10 vssd1 vccd1 sky130_fd_sc_hd__or4_1_1/C sky130_fd_sc_hd__ha_2_5/B
+ sky130_fd_sc_hd__nor2_1_42/B sky130_fd_sc_hd__ha_2_10/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_21 vssd1 vccd1 la_data_out[62] sky130_fd_sc_hd__ha_2_20/B sky130_fd_sc_hd__ha_2_21/SUM
+ sky130_fd_sc_hd__ha_2_21/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_32 vssd1 vccd1 sky130_fd_sc_hd__ha_2_32/A sky130_fd_sc_hd__ha_2_31/B
+ sky130_fd_sc_hd__ha_2_32/SUM la_data_out[39] vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_43 vssd1 vccd1 sky130_fd_sc_hd__ha_2_43/A sky130_fd_sc_hd__ha_2_42/B
+ sky130_fd_sc_hd__ha_2_43/SUM sky130_fd_sc_hd__ha_2_43/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__and2b_4_5 sky130_fd_sc_hd__or2b_2_1/A sky130_fd_sc_hd__and2b_4_5/X
+ sky130_fd_sc_hd__and3_4_9/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__and2b_4
Xsky130_fd_sc_hd__ha_2_54 vssd1 vccd1 sky130_fd_sc_hd__ha_2_54/A sky130_fd_sc_hd__ha_2_57/B
+ sky130_fd_sc_hd__ha_2_54/SUM sky130_fd_sc_hd__ha_2_54/B vssd1 vccd1 sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_6 vssd1 vccd1 sky130_fd_sc_hd__fa_2_281/A sky130_fd_sc_hd__dfxtp_2_5/Q
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__sdlclkp_4_50 sky130_fd_sc_hd__conb_1_148/LO sky130_fd_sc_hd__clkinv_8_67/A
+ sky130_fd_sc_hd__dfxtp_1_489/CLK sky130_fd_sc_hd__o21ai_1_911/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_130 sky130_fd_sc_hd__and3_4_15/A sky130_fd_sc_hd__nor2_1_130/Y
+ sky130_fd_sc_hd__and3_4_15/C vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_141 sky130_fd_sc_hd__nor2_1_145/Y sky130_fd_sc_hd__nor2_1_141/Y
+ sky130_fd_sc_hd__nor2_1_147/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_152 sky130_fd_sc_hd__nor2_1_152/B sky130_fd_sc_hd__nor2_1_152/Y
+ sky130_fd_sc_hd__nor2_1_152/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_1_6 la_data_out[121] sky130_fd_sc_hd__clkinv_1_6/A vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_163 sky130_fd_sc_hd__xor2_1_422/X sky130_fd_sc_hd__o21a_1_3/A2
+ sky130_fd_sc_hd__a211o_1_1/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_50 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__clkbuf_1_25/X
+ sky130_fd_sc_hd__nand2_1_74/B sky130_fd_sc_hd__dfxtp_1_136/Q sky130_fd_sc_hd__a22oi_1_50/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_174 sky130_fd_sc_hd__and3_1_2/B sky130_fd_sc_hd__nor2_1_174/Y
+ sky130_fd_sc_hd__and3_1_2/C vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_185 sky130_fd_sc_hd__nor2_1_73/B sky130_fd_sc_hd__nor2_1_185/Y
+ sky130_fd_sc_hd__buf_4_3/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_61 sky130_fd_sc_hd__clkbuf_1_24/X sky130_fd_sc_hd__clkbuf_1_23/X
+ sky130_fd_sc_hd__dfxtp_1_109/Q sky130_fd_sc_hd__dfxtp_1_77/Q sky130_fd_sc_hd__a22oi_1_61/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_72 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__nor2_4_3/Y
+ sky130_fd_sc_hd__nand2_1_63/B sky130_fd_sc_hd__dfxtp_1_147/Q sky130_fd_sc_hd__a22oi_1_72/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_196 sky130_fd_sc_hd__fah_1_9/SUM sky130_fd_sc_hd__nor2_2_28/A
+ sky130_fd_sc_hd__nor2_1_196/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_83 sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__dfxtp_1_120/Q sky130_fd_sc_hd__dfxtp_1_88/Q sky130_fd_sc_hd__a22oi_1_83/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_94 sky130_fd_sc_hd__buf_2_18/X sky130_fd_sc_hd__nor2_4_3/Y
+ sky130_fd_sc_hd__nand2_1_59/B sky130_fd_sc_hd__dfxtp_1_158/Q sky130_fd_sc_hd__a22oi_1_94/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_370 sky130_fd_sc_hd__buf_12_96/X sky130_fd_sc_hd__buf_12_554/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_381 sky130_fd_sc_hd__buf_12_381/A sky130_fd_sc_hd__buf_12_503/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_392 sky130_fd_sc_hd__buf_12_392/A sky130_fd_sc_hd__buf_12_392/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xnor2_1_100 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_100/B sky130_fd_sc_hd__inv_2_36/A
+ sky130_fd_sc_hd__xnor2_1_100/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_111 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_396/A sky130_fd_sc_hd__and3_4_10/C
+ sky130_fd_sc_hd__xnor2_1_114/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_122 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_124/A sky130_fd_sc_hd__and3_4_12/C
+ sky130_fd_sc_hd__xor2_1_418/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_570 sky130_fd_sc_hd__o21ai_1_780/A2 sky130_fd_sc_hd__xnor2_1_159/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_133 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_133/B sky130_fd_sc_hd__xnor2_1_133/Y
+ sky130_fd_sc_hd__xnor2_1_133/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_581 sky130_fd_sc_hd__nand2_1_600/A sky130_fd_sc_hd__nor2_1_194/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_144 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_504/A sky130_fd_sc_hd__and3_4_23/B
+ sky130_fd_sc_hd__xnor2_1_147/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_592 sky130_fd_sc_hd__nand2_1_617/A sky130_fd_sc_hd__nor2_1_203/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_155 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_155/B sky130_fd_sc_hd__xnor2_1_155/Y
+ sky130_fd_sc_hd__xnor2_1_155/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_166 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_166/B sky130_fd_sc_hd__xnor2_1_166/Y
+ sky130_fd_sc_hd__xnor2_1_166/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_177 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_177/B sky130_fd_sc_hd__inv_2_49/A
+ sky130_fd_sc_hd__xnor2_1_177/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_188 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_188/B sky130_fd_sc_hd__and2_0_277/A
+ sky130_fd_sc_hd__xnor2_1_188/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_4_50 sky130_fd_sc_hd__clkinv_4_50/A sky130_fd_sc_hd__clkinv_4_50/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__xnor2_1_199 vssd1 vccd1 sky130_fd_sc_hd__xnor2_1_199/B sky130_fd_sc_hd__and2_0_255/A
+ sky130_fd_sc_hd__xnor2_1_199/A vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_4_61 sky130_fd_sc_hd__clkinv_4_61/A sky130_fd_sc_hd__clkinv_4_61/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_72 sky130_fd_sc_hd__clkinv_4_72/A sky130_fd_sc_hd__clkinv_4_72/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_83 wbs_dat_i[23] sky130_fd_sc_hd__clkinv_4_83/Y vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_94 sky130_fd_sc_hd__nand2_1_16/Y sky130_fd_sc_hd__clkinv_4_94/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_1020 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1031 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1042 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1053 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1064 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__inv_16_2/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__decap_12_1075 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_506 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_7/X sky130_fd_sc_hd__nand2_1_385/Y
+ sky130_fd_sc_hd__a21oi_1_82/Y sky130_fd_sc_hd__xnor2_1_87/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1086 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_517 vssd1 vccd1 sky130_fd_sc_hd__buf_2_10/X sky130_fd_sc_hd__nand2b_1_14/Y
+ sky130_fd_sc_hd__o21ai_1_517/B1 sky130_fd_sc_hd__xor2_1_315/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_1097 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_528 vssd1 vccd1 sky130_fd_sc_hd__buf_2_7/X sky130_fd_sc_hd__nand2b_1_14/Y
+ sky130_fd_sc_hd__o21ai_1_528/B1 sky130_fd_sc_hd__xor2_1_327/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_539 vssd1 vccd1 sky130_fd_sc_hd__inv_2_31/Y sky130_fd_sc_hd__nand2b_2_3/Y
+ sky130_fd_sc_hd__o21ai_1_539/B1 sky130_fd_sc_hd__xor2_1_337/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_300 sky130_fd_sc_hd__fa_2_250/A sky130_fd_sc_hd__fa_2_207/B
+ sky130_fd_sc_hd__xor2_1_300/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_311 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__fa_2_213/B
+ sky130_fd_sc_hd__xor2_1_311/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_322 sky130_fd_sc_hd__dfxtp_2_5/Q sky130_fd_sc_hd__fa_2_216/A
+ sky130_fd_sc_hd__xor2_1_322/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_333 sky130_fd_sc_hd__or2_0_51/A sky130_fd_sc_hd__xor2_1_333/X
+ sky130_fd_sc_hd__xor2_1_333/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_344 sky130_fd_sc_hd__fa_2_239/A sky130_fd_sc_hd__and3_4_15/A
+ sky130_fd_sc_hd__xor2_1_344/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_355 sky130_fd_sc_hd__fa_2_250/A sky130_fd_sc_hd__fa_2_246/B
+ sky130_fd_sc_hd__xor2_1_355/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_366 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__fa_2_249/A
+ sky130_fd_sc_hd__xor2_1_366/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_377 sky130_fd_sc_hd__fa_2_262/A sky130_fd_sc_hd__fa_2_258/B
+ sky130_fd_sc_hd__xor2_1_377/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_388 sky130_fd_sc_hd__fa_2_281/A sky130_fd_sc_hd__fa_2_266/A
+ sky130_fd_sc_hd__xor2_1_388/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_399 sky130_fd_sc_hd__xor2_1_399/B sky130_fd_sc_hd__xor2_1_399/X
+ sky130_fd_sc_hd__xor2_1_399/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_304 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_88/A sky130_fd_sc_hd__clkbuf_1_304/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_315 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_315/X sky130_fd_sc_hd__clkinv_1_989/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_326 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_326/X sky130_fd_sc_hd__buf_8_61/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_337 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1_5/D sky130_fd_sc_hd__dfxtp_1_6/Q
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_408 vccd1 vssd1 sky130_fd_sc_hd__and3_4_26/X sky130_fd_sc_hd__nor2_1_87/A
+ sky130_fd_sc_hd__nor2_1_85/B sky130_fd_sc_hd__nor2_2_31/Y sky130_fd_sc_hd__nor2_2_10/B
+ sky130_fd_sc_hd__o21ai_1_676/B1 sky130_fd_sc_hd__nor2b_1_12/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_348 vssd1 vccd1 sky130_fd_sc_hd__inv_2_2/A sky130_fd_sc_hd__a222oi_1_8/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_419 vccd1 vssd1 sky130_fd_sc_hd__and3_4_21/X sky130_fd_sc_hd__buf_4_2/X
+ sky130_fd_sc_hd__buf_4_4/X sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__o21ai_1_690/B1 sky130_fd_sc_hd__and2b_4_12/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_359 vssd1 vccd1 la_data_out[37] sky130_fd_sc_hd__nor2_1_277/B
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_30 sky130_fd_sc_hd__dfxtp_1_30/Q sky130_fd_sc_hd__dfxtp_2_7/CLK
+ sky130_fd_sc_hd__and2_0_0/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_41 sky130_fd_sc_hd__nand2_1_73/B sky130_fd_sc_hd__dfxtp_1_62/CLK
+ sky130_fd_sc_hd__dfxtp_1_41/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_52 sky130_fd_sc_hd__nand2_1_62/B sky130_fd_sc_hd__dfxtp_1_57/CLK
+ sky130_fd_sc_hd__dfxtp_1_52/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_63 sky130_fd_sc_hd__dfxtp_1_63/Q sky130_fd_sc_hd__dfxtp_1_65/CLK
+ sky130_fd_sc_hd__dfxtp_1_63/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_74 sky130_fd_sc_hd__dfxtp_1_74/Q sky130_fd_sc_hd__dfxtp_1_81/CLK
+ sky130_fd_sc_hd__dfxtp_1_74/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_85 sky130_fd_sc_hd__dfxtp_1_85/Q sky130_fd_sc_hd__dfxtp_1_85/CLK
+ sky130_fd_sc_hd__dfxtp_1_85/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_96 sky130_fd_sc_hd__dfxtp_1_96/Q sky130_fd_sc_hd__dfxtp_1_97/CLK
+ sky130_fd_sc_hd__dfxtp_1_96/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_302 vccd1 vssd1 sky130_fd_sc_hd__or2_0_95/B sky130_fd_sc_hd__and2_0_302/B
+ sky130_fd_sc_hd__or2_0_98/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_313 vccd1 vssd1 sky130_fd_sc_hd__and2_0_313/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_313/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_324 vccd1 vssd1 sky130_fd_sc_hd__and2_0_324/X sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_324/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_335 vccd1 vssd1 sky130_fd_sc_hd__and2_0_398/A sky130_fd_sc_hd__ha_2_42/SUM
+ sky130_fd_sc_hd__and2_0_342/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_346 vccd1 vssd1 sky130_fd_sc_hd__and2_0_346/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__clkbuf_4_7/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_357 vccd1 vssd1 sky130_fd_sc_hd__and2_0_357/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__buf_2_184/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_368 vccd1 vssd1 sky130_fd_sc_hd__and2_0_368/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_60/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_379 vccd1 vssd1 sky130_fd_sc_hd__and2_0_379/X sky130_fd_sc_hd__buf_6_91/X
+ sky130_fd_sc_hd__a22o_1_58/X vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__inv_2_102 wbs_dat_i[10] sky130_fd_sc_hd__inv_2_102/Y vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_113 sky130_fd_sc_hd__inv_2_113/A sky130_fd_sc_hd__inv_2_113/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__or2_0_4 sky130_fd_sc_hd__or2_0_9/A sky130_fd_sc_hd__or2_0_4/X sky130_fd_sc_hd__or2_0_4/B
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__inv_2_124 sky130_fd_sc_hd__inv_2_124/A sky130_fd_sc_hd__inv_2_169/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_135 sky130_fd_sc_hd__inv_2_135/A sky130_fd_sc_hd__inv_2_135/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_146 sky130_fd_sc_hd__buf_8_25/A sky130_fd_sc_hd__inv_2_147/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_157 sky130_fd_sc_hd__inv_2_157/A sky130_fd_sc_hd__inv_2_157/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_168 sky130_fd_sc_hd__inv_2_168/A sky130_fd_sc_hd__buf_8_64/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_179 sky130_fd_sc_hd__inv_2_179/A sky130_fd_sc_hd__inv_2_179/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__o22ai_1_109 sky130_fd_sc_hd__xnor2_1_264/Y sky130_fd_sc_hd__xnor2_1_258/Y
+ sky130_fd_sc_hd__fa_2_448/CIN sky130_fd_sc_hd__nor2b_1_19/A sky130_fd_sc_hd__o22ai_1_66/B2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o31ai_2_0 sky130_fd_sc_hd__ha_2_9/B sky130_fd_sc_hd__o31ai_2_0/Y
+ sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__nand4_1_0/Y sky130_fd_sc_hd__o31ai_2_0/A2
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o31ai_2
Xsky130_fd_sc_hd__a211o_1_3 vssd1 vccd1 sky130_fd_sc_hd__fa_2_281/B sky130_fd_sc_hd__dfxtp_1_66/Q
+ sky130_fd_sc_hd__nor2_1_7/Y sky130_fd_sc_hd__inv_2_53/Y sky130_fd_sc_hd__o22ai_1_3/Y
+ vssd1 vccd1 sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__o21ai_1_303 vssd1 vccd1 sky130_fd_sc_hd__nand2_4_4/Y sky130_fd_sc_hd__nand2b_1_6/Y
+ sky130_fd_sc_hd__a22oi_1_195/Y sky130_fd_sc_hd__xor2_1_123/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_314 vssd1 vccd1 sky130_fd_sc_hd__a21oi_1_57/Y sky130_fd_sc_hd__nor2_1_74/A
+ sky130_fd_sc_hd__a21oi_1_49/Y sky130_fd_sc_hd__o21ai_1_314/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_325 vssd1 vccd1 sky130_fd_sc_hd__inv_2_22/Y sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__o21ai_1_325/B1 sky130_fd_sc_hd__xor2_1_145/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_336 vssd1 vccd1 sky130_fd_sc_hd__inv_2_18/Y sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__o21ai_1_336/B1 sky130_fd_sc_hd__xor2_1_155/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_347 vssd1 vccd1 sky130_fd_sc_hd__nand2_4_4/Y sky130_fd_sc_hd__nand2b_1_1/Y
+ sky130_fd_sc_hd__a22oi_1_197/Y sky130_fd_sc_hd__xor2_1_164/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_358 vssd1 vccd1 sky130_fd_sc_hd__inv_2_16/Y sky130_fd_sc_hd__nand2b_2_1/Y
+ sky130_fd_sc_hd__o21ai_1_358/B1 sky130_fd_sc_hd__xor2_1_174/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_369 vssd1 vccd1 sky130_fd_sc_hd__inv_2_26/Y sky130_fd_sc_hd__nand2b_2_0/Y
+ sky130_fd_sc_hd__nand2_1_159/Y sky130_fd_sc_hd__xor2_1_182/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nand2_1_707 sky130_fd_sc_hd__nand2_1_707/Y sky130_fd_sc_hd__or2_0_82/A
+ sky130_fd_sc_hd__or2_0_82/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_718 sky130_fd_sc_hd__o22ai_1_78/B2 sky130_fd_sc_hd__nor2b_1_20/A
+ sky130_fd_sc_hd__xor2_1_670/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_16 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_16/A1 sky130_fd_sc_hd__buf_2_94/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__or2_0_76/A vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nand2_1_729 sky130_fd_sc_hd__nand2_1_729/Y sky130_fd_sc_hd__or2_0_87/A
+ sky130_fd_sc_hd__or2_0_87/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__mux2_2_27 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_27/A1 sky130_fd_sc_hd__buf_2_146/X
+ sky130_fd_sc_hd__mux2_8_0/S sky130_fd_sc_hd__mux2_2_27/X vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_38 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_38/A1 sky130_fd_sc_hd__buf_2_151/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__mux2_2_38/X vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_49 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_49/A1 sky130_fd_sc_hd__buf_4_16/X
+ sky130_fd_sc_hd__mux2_4_4/S sky130_fd_sc_hd__mux2_2_49/X vssd1 vccd1 sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__conb_1_102 sky130_fd_sc_hd__conb_1_102/LO sky130_fd_sc_hd__conb_1_102/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_113 sky130_fd_sc_hd__conb_1_113/LO sky130_fd_sc_hd__conb_1_113/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_124 sky130_fd_sc_hd__conb_1_124/LO sky130_fd_sc_hd__conb_1_124/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_135 sky130_fd_sc_hd__conb_1_135/LO sky130_fd_sc_hd__clkinv_1_7/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_146 sky130_fd_sc_hd__buf_6_7/A sky130_fd_sc_hd__conb_1_146/HI
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__xor2_1_130 sky130_fd_sc_hd__fa_2_97/A sky130_fd_sc_hd__fa_2_97/CIN
+ sky130_fd_sc_hd__xor2_1_130/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_141 sky130_fd_sc_hd__fa_2_122/A sky130_fd_sc_hd__fa_2_105/B
+ sky130_fd_sc_hd__xor2_1_141/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_152 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__fa_2_109/B
+ sky130_fd_sc_hd__xor2_1_152/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_503 sky130_fd_sc_hd__or4_1_3/D sky130_fd_sc_hd__dfxtp_1_509/CLK
+ sky130_fd_sc_hd__and2_0_392/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_163 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__fa_2_116/B
+ sky130_fd_sc_hd__xor2_1_163/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_514 sky130_fd_sc_hd__ha_2_56/A sky130_fd_sc_hd__dfxtp_1_515/CLK
+ sky130_fd_sc_hd__and2_0_347/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_174 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__fa_2_124/A
+ sky130_fd_sc_hd__xor2_1_174/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_525 wbs_dat_o[4] sky130_fd_sc_hd__dfxtp_1_533/CLK sky130_fd_sc_hd__nor2b_1_153/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_185 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__fa_2_132/A
+ sky130_fd_sc_hd__xor2_1_185/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_536 wbs_dat_o[15] sky130_fd_sc_hd__dfxtp_1_538/CLK sky130_fd_sc_hd__nor2b_1_142/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_196 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__xor2_1_196/X
+ sky130_fd_sc_hd__xor2_1_196/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_547 wbs_dat_o[26] sky130_fd_sc_hd__dfxtp_1_552/CLK sky130_fd_sc_hd__nor2b_1_131/Y
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_101 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_16/A1 sky130_fd_sc_hd__clkbuf_1_101/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_112 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_112/X sky130_fd_sc_hd__clkinv_1_970/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_123 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1_123/X sky130_fd_sc_hd__inv_2_2/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_134 vssd1 vccd1 sky130_fd_sc_hd__buf_8_133/A sky130_fd_sc_hd__clkbuf_1_52/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_205 vccd1 vssd1 sky130_fd_sc_hd__and3_4_0/X sky130_fd_sc_hd__buf_4_1/X
+ sky130_fd_sc_hd__nor2_2_5/A sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__nor2_2_5/B
+ sky130_fd_sc_hd__o21ai_1_377/B1 sky130_fd_sc_hd__and2b_4_1/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_145 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_18/A1 sky130_fd_sc_hd__clkbuf_1_145/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_216 vccd1 vssd1 sky130_fd_sc_hd__and3_1_1/X sky130_fd_sc_hd__buf_2_32/X
+ sky130_fd_sc_hd__buf_8_0/X sky130_fd_sc_hd__nor2_1_117/Y sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__o21ai_1_404/B1 sky130_fd_sc_hd__nor2b_1_8/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__dfxtp_1_3 sky130_fd_sc_hd__buf_8_79/A sky130_fd_sc_hd__dfxtp_1_3/CLK
+ sky130_fd_sc_hd__dfxtp_1_3/D vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_156 vssd1 vccd1 sky130_fd_sc_hd__mux2_2_24/A1 sky130_fd_sc_hd__clkbuf_1_156/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_227 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__or2_0_61/A
+ sky130_fd_sc_hd__or2_0_42/B sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__or2_0_39/B
+ sky130_fd_sc_hd__o21ai_1_418/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_167 vssd1 vccd1 sky130_fd_sc_hd__buf_8_78/A sky130_fd_sc_hd__buf_2_159/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a222oi_1_238 vccd1 vssd1 sky130_fd_sc_hd__and3_4_12/X sky130_fd_sc_hd__or2_0_60/A
+ sky130_fd_sc_hd__or2_0_61/A sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__or2_0_42/B
+ sky130_fd_sc_hd__o21ai_1_432/B1 sky130_fd_sc_hd__and2b_4_6/X vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_178 vssd1 vccd1 sky130_fd_sc_hd__a22o_1_25/B2 sky130_fd_sc_hd__clkbuf_1_178/A
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o21ai_1_870 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_648/A sky130_fd_sc_hd__nor2_1_229/Y
+ sky130_fd_sc_hd__nand2_1_697/Y sky130_fd_sc_hd__xnor2_1_196/B vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_249 vccd1 vssd1 sky130_fd_sc_hd__and3_4_13/X sky130_fd_sc_hd__buf_2_32/X
+ sky130_fd_sc_hd__buf_8_0/X sky130_fd_sc_hd__nor2_1_121/Y sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__o21ai_1_447/B1 sky130_fd_sc_hd__nor2b_1_9/Y vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__clkbuf_1_189 vssd1 vccd1 sky130_fd_sc_hd__buf_12_12/A sky130_fd_sc_hd__clkbuf_1_51/X
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o21ai_1_881 vssd1 vccd1 sky130_fd_sc_hd__xor2_1_658/B sky130_fd_sc_hd__nor2_1_241/Y
+ sky130_fd_sc_hd__nand2_1_752/Y sky130_fd_sc_hd__xnor2_1_211/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_408 sky130_fd_sc_hd__fa_2_406/B sky130_fd_sc_hd__fa_2_409/A
+ sky130_fd_sc_hd__fa_2_408/A sky130_fd_sc_hd__fa_2_408/B sky130_fd_sc_hd__fa_2_408/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o21ai_1_892 vssd1 vccd1 sky130_fd_sc_hd__nand4_1_0/Y sky130_fd_sc_hd__inv_2_67/A
+ sky130_fd_sc_hd__o31ai_2_0/B1 sky130_fd_sc_hd__o21ai_1_892/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_419 sky130_fd_sc_hd__fa_2_418/CIN sky130_fd_sc_hd__fa_2_419/SUM
+ sky130_fd_sc_hd__fa_2_419/A sky130_fd_sc_hd__fa_2_419/B sky130_fd_sc_hd__fa_2_419/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_4_13 sky130_fd_sc_hd__inv_4_13/Y sky130_fd_sc_hd__inv_4_13/A
+ vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__and2_0_110 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_32/D sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__and2_0_110/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_121 vccd1 vssd1 sky130_fd_sc_hd__and2_0_121/X sky130_fd_sc_hd__o21ai_2_0/B1
+ sky130_fd_sc_hd__and2_0_121/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_8_1 sky130_fd_sc_hd__nand2_8_1/A sky130_fd_sc_hd__nand2_8_1/B
+ sky130_fd_sc_hd__nor2_2_10/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_8
Xsky130_fd_sc_hd__and2_0_132 vccd1 vssd1 sky130_fd_sc_hd__and2_0_132/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_132/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_40 la_data_out[23] sky130_fd_sc_hd__conb_1_102/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_143 vccd1 vssd1 sky130_fd_sc_hd__and2_0_143/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_143/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_51 la_data_out[12] sky130_fd_sc_hd__conb_1_91/HI vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_154 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_41/D sky130_fd_sc_hd__buf_2_16/A
+ sky130_fd_sc_hd__and2_0_154/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_62 la_data_out[1] sky130_fd_sc_hd__conb_1_80/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_165 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_75/D sky130_fd_sc_hd__o21ai_2_0/B1
+ sky130_fd_sc_hd__and2_0_165/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_73 io_out[28] sky130_fd_sc_hd__conb_1_69/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_176 vccd1 vssd1 sky130_fd_sc_hd__and2_0_176/X sky130_fd_sc_hd__o21ai_2_0/B1
+ sky130_fd_sc_hd__and2_0_176/A vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_84 io_out[17] sky130_fd_sc_hd__conb_1_58/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_187 vccd1 vssd1 sky130_fd_sc_hd__and2_0_187/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_93/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_95 io_out[6] sky130_fd_sc_hd__conb_1_47/HI vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_198 vccd1 vssd1 sky130_fd_sc_hd__and2_0_198/X sky130_fd_sc_hd__buf_2_16/X
+ sky130_fd_sc_hd__o21ai_1_84/Y vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__sdlclkp_1_4 sky130_fd_sc_hd__conb_1_145/LO sky130_fd_sc_hd__clkinv_8_7/Y
+ sky130_fd_sc_hd__clkinv_2_14/A sky130_fd_sc_hd__o31ai_2_0/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__sdlclkp_1
Xsky130_fd_sc_hd__o21ai_1_100 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_98/A2 sky130_fd_sc_hd__nand2_2_9/Y
+ sky130_fd_sc_hd__a22oi_1_160/Y sky130_fd_sc_hd__and2_0_177/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_111 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_113/A2 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_123/Y sky130_fd_sc_hd__and2_0_164/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_122 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_125/A2 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nand2_1_128/Y sky130_fd_sc_hd__and2_0_150/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_133 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_133/A2 sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__a22oi_1_177/Y sky130_fd_sc_hd__and2_0_137/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_144 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_145/A2 sky130_fd_sc_hd__inv_2_5/Y
+ sky130_fd_sc_hd__a22oi_1_182/Y sky130_fd_sc_hd__and2_0_123/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_155 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_157/A2 sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_145/Y sky130_fd_sc_hd__and2_0_109/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_166 vssd1 vccd1 sky130_fd_sc_hd__a21oi_1_65/Y sky130_fd_sc_hd__nand2_1_284/Y
+ sky130_fd_sc_hd__a21oi_1_60/Y sky130_fd_sc_hd__inv_2_11/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_177 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_177/A2 sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__a222oi_1_58/Y sky130_fd_sc_hd__xor2_1_10/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_188 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_209/A2 sky130_fd_sc_hd__nor2_1_47/A
+ sky130_fd_sc_hd__a21oi_1_39/Y sky130_fd_sc_hd__o21ai_1_188/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_199 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_199/A2 sky130_fd_sc_hd__or2b_2_0/X
+ sky130_fd_sc_hd__a222oi_1_75/Y sky130_fd_sc_hd__xor2_1_28/A vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_609 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_504 sky130_fd_sc_hd__nand2_1_517/B sky130_fd_sc_hd__nor2_2_22/A
+ sky130_fd_sc_hd__nor2_2_22/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_515 sky130_fd_sc_hd__xnor2_1_133/A sky130_fd_sc_hd__nand2_1_516/Y
+ sky130_fd_sc_hd__or2_0_56/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_526 sky130_fd_sc_hd__nand2_1_526/Y sky130_fd_sc_hd__or2_0_58/A
+ sky130_fd_sc_hd__or2_0_58/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_537 sky130_fd_sc_hd__nand2_1_537/Y sky130_fd_sc_hd__or2_0_61/A
+ sky130_fd_sc_hd__or2_0_61/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_548 sky130_fd_sc_hd__nand2_1_548/Y sky130_fd_sc_hd__or2_0_60/A
+ sky130_fd_sc_hd__or2_0_60/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_559 sky130_fd_sc_hd__nand2_1_559/Y sky130_fd_sc_hd__or2_0_66/A
+ sky130_fd_sc_hd__buf_4_5/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_6 sky130_fd_sc_hd__and3_4_6/C sky130_fd_sc_hd__nor2b_1_6/Y
+ sky130_fd_sc_hd__and3_4_6/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1106 sky130_fd_sc_hd__clkinv_4_49/A sky130_fd_sc_hd__a22o_1_26/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1117 sky130_fd_sc_hd__clkinv_4_60/A sky130_fd_sc_hd__a22o_1_37/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1128 sky130_fd_sc_hd__clkinv_4_71/A sky130_fd_sc_hd__a22o_1_48/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1139 sky130_fd_sc_hd__a22o_1_79/A2 sky130_fd_sc_hd__clkinv_4_85/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_300 sky130_fd_sc_hd__dfxtp_1_300/Q sky130_fd_sc_hd__clkinv_8_6/Y
+ sky130_fd_sc_hd__and2_0_276/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1608 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_311 sky130_fd_sc_hd__or2_0_92/A sky130_fd_sc_hd__dfxtp_1_319/CLK
+ sky130_fd_sc_hd__and2_0_288/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1619 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_322 sky130_fd_sc_hd__nor2_1_235/A sky130_fd_sc_hd__dfxtp_1_323/CLK
+ sky130_fd_sc_hd__and2_0_299/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_333 sky130_fd_sc_hd__dfxtp_1_333/Q sky130_fd_sc_hd__dfxtp_1_339/CLK
+ sky130_fd_sc_hd__and2_0_334/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_344 sky130_fd_sc_hd__dfxtp_1_344/Q sky130_fd_sc_hd__dfxtp_1_354/CLK
+ sky130_fd_sc_hd__and2_0_313/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_355 sky130_fd_sc_hd__dfxtp_1_355/Q sky130_fd_sc_hd__dfxtp_1_356/CLK
+ sky130_fd_sc_hd__and2_0_306/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_366 sky130_fd_sc_hd__dfxtp_1_366/Q sky130_fd_sc_hd__dfxtp_1_371/CLK
+ sky130_fd_sc_hd__nor2b_1_117/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_377 sky130_fd_sc_hd__dfxtp_1_377/Q sky130_fd_sc_hd__dfxtp_1_380/CLK
+ sky130_fd_sc_hd__nor2b_1_106/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_388 sky130_fd_sc_hd__dfxtp_1_388/Q sky130_fd_sc_hd__dfxtp_1_395/CLK
+ sky130_fd_sc_hd__nor2b_1_95/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_8 sky130_fd_sc_hd__nand2_2_0/B sky130_fd_sc_hd__nand2_1_8/B
+ sky130_fd_sc_hd__or2_0_84/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_399 sky130_fd_sc_hd__dfxtp_1_399/Q sky130_fd_sc_hd__clkinv_4_8/Y
+ sky130_fd_sc_hd__nor2b_1_116/Y vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_205 sky130_fd_sc_hd__fa_2_201/B sky130_fd_sc_hd__fa_2_208/CIN
+ sky130_fd_sc_hd__fa_2_205/A sky130_fd_sc_hd__fa_2_205/B sky130_fd_sc_hd__fa_2_205/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_216 sky130_fd_sc_hd__fa_2_212/CIN sky130_fd_sc_hd__fa_2_222/A
+ sky130_fd_sc_hd__fa_2_216/A sky130_fd_sc_hd__fa_2_216/B sky130_fd_sc_hd__fa_2_221/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_227 sky130_fd_sc_hd__fa_2_216/B sky130_fd_sc_hd__fa_2_227/SUM
+ sky130_fd_sc_hd__fa_2_227/A sky130_fd_sc_hd__fa_2_227/B sky130_fd_sc_hd__xor2_1_326/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_238 sky130_fd_sc_hd__fa_2_234/B sky130_fd_sc_hd__fa_2_240/CIN
+ sky130_fd_sc_hd__fa_2_238/A sky130_fd_sc_hd__fa_2_238/B sky130_fd_sc_hd__fa_2_238/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_249 sky130_fd_sc_hd__fah_1_4/CI sky130_fd_sc_hd__fah_1_2/A
+ sky130_fd_sc_hd__fa_2_249/A sky130_fd_sc_hd__fa_2_249/B sky130_fd_sc_hd__xor2_1_364/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_30 sky130_fd_sc_hd__fa_2_23/A sky130_fd_sc_hd__fa_2_29/B sky130_fd_sc_hd__fa_2_30/A
+ sky130_fd_sc_hd__fa_2_30/B sky130_fd_sc_hd__fa_2_30/CIN vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_41 sky130_fd_sc_hd__fa_2_35/B sky130_fd_sc_hd__fa_2_43/CIN
+ sky130_fd_sc_hd__fa_2_41/A sky130_fd_sc_hd__fa_2_41/B sky130_fd_sc_hd__fa_2_41/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_9 vccd1 vssd1 sky130_fd_sc_hd__and2_0_9/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__or2_0_72/B vssd1 vccd1 sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__fa_2_52 sky130_fd_sc_hd__fa_2_47/CIN sky130_fd_sc_hd__fa_2_59/A
+ sky130_fd_sc_hd__fa_2_52/A sky130_fd_sc_hd__fa_2_52/B sky130_fd_sc_hd__fa_2_57/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_63 sky130_fd_sc_hd__fa_2_59/B sky130_fd_sc_hd__fa_2_66/CIN
+ sky130_fd_sc_hd__fa_2_63/A sky130_fd_sc_hd__fa_2_63/B sky130_fd_sc_hd__fa_2_63/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_74 sky130_fd_sc_hd__fa_2_70/CIN sky130_fd_sc_hd__fa_2_80/A
+ sky130_fd_sc_hd__fa_2_74/A sky130_fd_sc_hd__fa_2_74/B sky130_fd_sc_hd__fa_2_79/SUM
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_85 sky130_fd_sc_hd__fa_2_74/B sky130_fd_sc_hd__fa_2_85/SUM
+ sky130_fd_sc_hd__fa_2_85/A sky130_fd_sc_hd__fa_2_85/B sky130_fd_sc_hd__fa_2_85/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_96 sky130_fd_sc_hd__fa_2_92/B sky130_fd_sc_hd__fa_2_98/CIN
+ sky130_fd_sc_hd__fa_2_96/A sky130_fd_sc_hd__fa_2_96/B sky130_fd_sc_hd__fa_2_96/CIN
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_200 vccd1 vssd1 la_data_out[88] sky130_fd_sc_hd__nand2_2_5/Y
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_211 vccd1 vssd1 sky130_fd_sc_hd__buf_2_211/X sky130_fd_sc_hd__or2_0_84/B
+ vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__a21oi_1_13 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_42/Y
+ sky130_fd_sc_hd__a21oi_1_13/Y sky130_fd_sc_hd__dfxtp_1_84/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_24 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__o22ai_1_53/Y
+ sky130_fd_sc_hd__a21oi_1_24/Y sky130_fd_sc_hd__dfxtp_1_73/Q vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_35 sky130_fd_sc_hd__o21ai_1_161/Y sky130_fd_sc_hd__a21oi_1_35/B1
+ sky130_fd_sc_hd__inv_2_25/A sky130_fd_sc_hd__or2_0_0/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_580 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_406/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_438/Q sky130_fd_sc_hd__clkbuf_1_32/X
+ sky130_fd_sc_hd__clkinv_1_777/A sky130_fd_sc_hd__dfxtp_1_374/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a21oi_1_46 sky130_fd_sc_hd__nand2_1_229/Y sky130_fd_sc_hd__o21ai_1_263/Y
+ sky130_fd_sc_hd__o21a_1_0/A2 sky130_fd_sc_hd__nor2_1_64/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_591 vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1_401/Q sky130_fd_sc_hd__nor2_4_19/Y
+ sky130_fd_sc_hd__and2b_4_13/X sky130_fd_sc_hd__dfxtp_1_433/Q sky130_fd_sc_hd__clkbuf_1_32/X
+ sky130_fd_sc_hd__clkinv_1_788/A sky130_fd_sc_hd__dfxtp_1_369/Q vssd1 vccd1 sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a21oi_1_57 sky130_fd_sc_hd__nor2_1_84/Y sky130_fd_sc_hd__nand2_1_261/Y
+ sky130_fd_sc_hd__a21oi_1_57/Y sky130_fd_sc_hd__nand2_1_272/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_68 sky130_fd_sc_hd__xor2_1_211/X sky130_fd_sc_hd__a21oi_1_68/B1
+ sky130_fd_sc_hd__o21a_1_1/A1 sky130_fd_sc_hd__or2_0_24/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_79 sky130_fd_sc_hd__a21oi_1_80/A1 sky130_fd_sc_hd__a21oi_1_79/B1
+ sky130_fd_sc_hd__a21oi_1_79/Y sky130_fd_sc_hd__nand2_1_368/B vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__nor3_1_5 sky130_fd_sc_hd__nor3_1_5/C sky130_fd_sc_hd__nor3_1_5/Y
+ wbs_adr_i[18] wbs_adr_i[0] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__decap_12_20 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_31 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_42 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_53 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_64 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_75 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_86 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_97 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_20 vccd1 vssd1 sky130_fd_sc_hd__buf_6_20/X sky130_fd_sc_hd__buf_6_20/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_31 vccd1 vssd1 sky130_fd_sc_hd__buf_6_31/X sky130_fd_sc_hd__buf_6_31/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_42 vccd1 vssd1 sky130_fd_sc_hd__buf_6_42/X sky130_fd_sc_hd__buf_6_42/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_53 vccd1 vssd1 sky130_fd_sc_hd__buf_6_53/X sky130_fd_sc_hd__buf_8_91/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_64 vccd1 vssd1 sky130_fd_sc_hd__buf_6_64/X sky130_fd_sc_hd__buf_8_79/X
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_75 vccd1 vssd1 sky130_fd_sc_hd__buf_6_75/X sky130_fd_sc_hd__buf_6_75/A
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_86 vccd1 vssd1 sky130_fd_sc_hd__buf_6_86/X sky130_fd_sc_hd__inv_16_6/Y
+ vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_11 la_data_out[62] vssd1 vccd1 vccd1 vssd1 sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_22 sky130_fd_sc_hd__clkinv_4_71/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_33 sky130_fd_sc_hd__clkinv_4_74/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_44 sky130_fd_sc_hd__buf_2_189/A vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_55 sky130_fd_sc_hd__buf_2_192/A vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_66 sky130_fd_sc_hd__nand2_2_3/Y vssd1 vccd1 vccd1 vssd1
+ sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__decap_12_406 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_417 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_301 sky130_fd_sc_hd__nand2_1_301/Y sky130_fd_sc_hd__nand2_1_311/Y
+ sky130_fd_sc_hd__nand2_1_307/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_428 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_900 sky130_fd_sc_hd__clkinv_1_901/A sky130_fd_sc_hd__buf_2_47/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_312 sky130_fd_sc_hd__nand2_1_312/Y sky130_fd_sc_hd__xnor2_1_4/B
+ sky130_fd_sc_hd__nand2_1_316/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_439 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_911 sky130_fd_sc_hd__clkinv_1_911/Y sky130_fd_sc_hd__inv_2_105/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_323 sky130_fd_sc_hd__nand2_1_323/Y sky130_fd_sc_hd__nor2_1_117/Y
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_922 sky130_fd_sc_hd__inv_2_109/A sky130_fd_sc_hd__a21o_2_4/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_334 sky130_fd_sc_hd__or2_0_32/A sky130_fd_sc_hd__nor2_1_107/Y
+ sky130_fd_sc_hd__nor2_1_115/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_933 sky130_fd_sc_hd__inv_12_0/A sky130_fd_sc_hd__o21ai_1_926/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_345 sky130_fd_sc_hd__nand2_1_345/Y sky130_fd_sc_hd__nor2_1_110/A
+ sky130_fd_sc_hd__nor2_1_110/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_944 sky130_fd_sc_hd__inv_2_139/A sky130_fd_sc_hd__buf_8_6/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_356 sky130_fd_sc_hd__o21ai_2_11/B1 sky130_fd_sc_hd__nor2_2_11/A
+ sky130_fd_sc_hd__nor2_2_11/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_955 sky130_fd_sc_hd__clkinv_1_955/Y sky130_fd_sc_hd__inv_2_151/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_367 sky130_fd_sc_hd__nand2_1_367/Y sky130_fd_sc_hd__nor2_2_13/A
+ sky130_fd_sc_hd__nor2_2_13/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_966 sky130_fd_sc_hd__clkinv_2_30/A sky130_fd_sc_hd__buf_2_128/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_378 sky130_fd_sc_hd__nand2_1_378/Y sky130_fd_sc_hd__nor2_2_12/A
+ sky130_fd_sc_hd__nor2_2_12/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_977 sky130_fd_sc_hd__clkinv_1_977/Y sky130_fd_sc_hd__clkinv_4_95/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_389 sky130_fd_sc_hd__nand2_1_389/Y sky130_fd_sc_hd__nor2_1_124/A
+ sky130_fd_sc_hd__nor2_1_124/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_988 sky130_fd_sc_hd__clkinv_1_988/Y sky130_fd_sc_hd__clkinv_4_31/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_999 sky130_fd_sc_hd__clkinv_1_999/Y sky130_fd_sc_hd__inv_4_4/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1405 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1416 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1427 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_130 sky130_fd_sc_hd__dfxtp_1_130/Q sky130_fd_sc_hd__dfxtp_1_146/CLK
+ sky130_fd_sc_hd__and2_0_121/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1438 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_141 sky130_fd_sc_hd__dfxtp_1_141/Q sky130_fd_sc_hd__dfxtp_1_141/CLK
+ sky130_fd_sc_hd__and2_0_186/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_1449 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_152 sky130_fd_sc_hd__dfxtp_1_152/Q sky130_fd_sc_hd__dfxtp_1_152/CLK
+ sky130_fd_sc_hd__and2_0_231/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_163 sky130_fd_sc_hd__dfxtp_1_163/Q sky130_fd_sc_hd__dfxtp_1_170/CLK
+ sky130_fd_sc_hd__and2_0_122/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_174 sky130_fd_sc_hd__dfxtp_1_174/Q sky130_fd_sc_hd__dfxtp_1_176/CLK
+ sky130_fd_sc_hd__and2_0_177/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_185 sky130_fd_sc_hd__dfxtp_1_185/Q sky130_fd_sc_hd__clkinv_4_2/Y
+ sky130_fd_sc_hd__and2_0_232/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_196 sky130_fd_sc_hd__xor2_1_622/A sky130_fd_sc_hd__dfxtp_2_1/CLK
+ sky130_fd_sc_hd__and2_0_15/X vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_12_940 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_951 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_962 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_973 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_984 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_995 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o211ai_1_16 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_47/B1
+ sky130_fd_sc_hd__o211ai_1_16/Y sky130_fd_sc_hd__a22oi_1_64/Y sky130_fd_sc_hd__a22oi_1_65/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_27 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__o22ai_1_34/B1
+ sky130_fd_sc_hd__o211ai_1_27/Y sky130_fd_sc_hd__a22oi_1_86/Y sky130_fd_sc_hd__a22oi_1_87/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_38 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o21ai_1_8/A2
+ sky130_fd_sc_hd__fa_2_338/B sky130_fd_sc_hd__nand2_1_58/Y sky130_fd_sc_hd__a21oi_1_9/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_49 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__o22ai_1_14/B1
+ sky130_fd_sc_hd__fa_2_393/A sky130_fd_sc_hd__nand2_1_69/Y sky130_fd_sc_hd__a21oi_1_20/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o21ai_1_90 vssd1 vccd1 sky130_fd_sc_hd__o21ai_1_93/A2 sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__o21ai_1_90/B1 sky130_fd_sc_hd__o21ai_1_90/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkinv_1_207 sky130_fd_sc_hd__o22ai_1_13/B1 sky130_fd_sc_hd__dfxtp_1_108/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_218 sky130_fd_sc_hd__nor2_1_13/A sky130_fd_sc_hd__dfxtp_1_136/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_229 sky130_fd_sc_hd__o22ai_1_5/A2 sky130_fd_sc_hd__dfxtp_1_164/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_2_7 sky130_fd_sc_hd__o21ai_2_7/B1 sky130_fd_sc_hd__o21ai_2_7/Y
+ sky130_fd_sc_hd__o21ai_2_7/A2 sky130_fd_sc_hd__o21ai_2_7/A1 vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__o21ai_2
Xsky130_fd_sc_hd__a21oi_1_104 sky130_fd_sc_hd__xnor2_1_132/B sky130_fd_sc_hd__clkinv_1_518/Y
+ sky130_fd_sc_hd__a21oi_1_104/Y sky130_fd_sc_hd__or2_1_9/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_115 sky130_fd_sc_hd__clkinv_1_549/Y sky130_fd_sc_hd__nor2_1_176/A
+ sky130_fd_sc_hd__a21oi_1_115/Y sky130_fd_sc_hd__or2_0_59/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_126 sky130_fd_sc_hd__o21ai_1_828/Y sky130_fd_sc_hd__o21ai_1_811/Y
+ sky130_fd_sc_hd__o21ai_2_16/A2 sky130_fd_sc_hd__nor2_1_195/Y vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_137 sky130_fd_sc_hd__xor2_1_636/X sky130_fd_sc_hd__clkinv_1_611/Y
+ sky130_fd_sc_hd__o21a_1_5/A1 sky130_fd_sc_hd__or2_0_70/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_148 sky130_fd_sc_hd__xnor2_1_198/B sky130_fd_sc_hd__clkinv_1_645/Y
+ sky130_fd_sc_hd__xor2_1_649/A sky130_fd_sc_hd__or2_0_81/X vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_159 sky130_fd_sc_hd__or2_0_95/X sky130_fd_sc_hd__clkinv_1_676/Y
+ sky130_fd_sc_hd__xor2_1_658/B sky130_fd_sc_hd__xnor2_1_212/A vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_530 sky130_fd_sc_hd__buf_12_530/A sky130_fd_sc_hd__buf_12_530/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_541 sky130_fd_sc_hd__buf_12_541/A sky130_fd_sc_hd__buf_12_541/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_552 sky130_fd_sc_hd__buf_12_552/A sky130_fd_sc_hd__buf_12_552/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_563 sky130_fd_sc_hd__buf_12_563/A sky130_fd_sc_hd__buf_12_563/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_8_0 sky130_fd_sc_hd__buf_2_140/A sky130_fd_sc_hd__buf_6_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_8
Xsky130_fd_sc_hd__buf_12_574 sky130_fd_sc_hd__buf_12_574/A sky130_fd_sc_hd__buf_12_574/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_203 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_585 sky130_fd_sc_hd__buf_12_585/A sky130_fd_sc_hd__buf_12_585/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_214 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_596 sky130_fd_sc_hd__buf_12_596/A sky130_fd_sc_hd__buf_12_596/X
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_225 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_236 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_120 sky130_fd_sc_hd__nand2_1_120/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__xnor2_1_104/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_247 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_131 sky130_fd_sc_hd__nand2_1_131/Y sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nand2_1_131/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_258 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_730 sky130_fd_sc_hd__nor2b_1_109/A sky130_fd_sc_hd__xnor2_1_298/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_142 sky130_fd_sc_hd__nand2_1_142/Y sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__xor2_1_419/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_269 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_741 sky130_fd_sc_hd__fa_2_461/A sky130_fd_sc_hd__clkinv_1_741/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_304 vssd1 vccd1 sky130_fd_sc_hd__maj3_1_1/A sky130_fd_sc_hd__nand4_1_2/D
+ la_data_out[41] vssd1 vccd1 sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_153 sky130_fd_sc_hd__nand2_1_153/Y sky130_fd_sc_hd__nor2_1_56/Y
+ sky130_fd_sc_hd__or2_0_52/B vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_752 sky130_fd_sc_hd__fa_2_475/A sky130_fd_sc_hd__clkinv_1_752/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_164 sky130_fd_sc_hd__nor2_1_46/A sky130_fd_sc_hd__or2_0_9/X
+ sky130_fd_sc_hd__or2_0_10/X vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_763 sky130_fd_sc_hd__fa_2_486/A sky130_fd_sc_hd__clkinv_1_763/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_175 sky130_fd_sc_hd__nand2_1_175/Y sky130_fd_sc_hd__nor2_1_50/Y
+ sky130_fd_sc_hd__nand2_1_203/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_774 sky130_fd_sc_hd__and2_0_333/A sky130_fd_sc_hd__clkinv_1_774/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_186 sky130_fd_sc_hd__nand2_1_186/Y sky130_fd_sc_hd__nor2_1_54/Y
+ sky130_fd_sc_hd__nand2_1_203/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_785 sky130_fd_sc_hd__and2_0_322/A sky130_fd_sc_hd__clkinv_1_785/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_197 sky130_fd_sc_hd__nand2_1_197/Y sky130_fd_sc_hd__nand2_1_197/B
+ sky130_fd_sc_hd__nand2_1_203/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_796 sky130_fd_sc_hd__and2_0_311/A sky130_fd_sc_hd__clkinv_1_796/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1202 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_2 sky130_fd_sc_hd__fa_2_56/A sky130_fd_sc_hd__xor3_1_4/C
+ sky130_fd_sc_hd__xor2_1_2/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_1213 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1224 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1235 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1246 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1257 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1268 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1279 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_8_0 sky130_fd_sc_hd__clkinv_8_1/A sky130_fd_sc_hd__clkinv_8_2/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__xor2_1_17 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__fa_2_2/A
+ sky130_fd_sc_hd__xor2_1_17/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_28 sky130_fd_sc_hd__or2_0_24/A sky130_fd_sc_hd__fa_2_11/B
+ sky130_fd_sc_hd__xor2_1_28/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_39 sky130_fd_sc_hd__xor2_1_9/B sky130_fd_sc_hd__fa_2_21/A
+ sky130_fd_sc_hd__xor2_1_39/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_12_770 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_781 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_792 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__xor2_1_504 sky130_fd_sc_hd__fa_2_338/A sky130_fd_sc_hd__and3_4_23/A
+ sky130_fd_sc_hd__xor2_1_504/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_515 sky130_fd_sc_hd__fah_1_14/A sky130_fd_sc_hd__xor2_1_515/X
+ sky130_fd_sc_hd__xor2_1_515/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_526 sky130_fd_sc_hd__xor2_1_526/B sky130_fd_sc_hd__inv_2_61/A
+ sky130_fd_sc_hd__xor2_1_526/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_537 sky130_fd_sc_hd__fah_1_14/A sky130_fd_sc_hd__fa_2_365/B
+ sky130_fd_sc_hd__xor2_1_537/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_548 sky130_fd_sc_hd__xor2_1_548/B sky130_fd_sc_hd__fa_2_373/B
+ sky130_fd_sc_hd__xor2_1_548/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_559 sky130_fd_sc_hd__xor2_1_559/B sky130_fd_sc_hd__xor2_1_559/X
+ sky130_fd_sc_hd__xor2_1_559/A vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__xor2_1
.ends

