magic
tech sky130A
magscale 1 2
timestamp 1655789722
<< metal1 >>
rect 3878 700748 3884 700800
rect 3936 700788 3942 700800
rect 8110 700788 8116 700800
rect 3936 700760 8116 700788
rect 3936 700748 3942 700760
rect 8110 700748 8116 700760
rect 8168 700748 8174 700800
rect 102042 700748 102048 700800
rect 102100 700788 102106 700800
rect 105446 700788 105452 700800
rect 102100 700760 105452 700788
rect 102100 700748 102106 700760
rect 105446 700748 105452 700760
rect 105504 700748 105510 700800
rect 200022 700748 200028 700800
rect 200080 700788 200086 700800
rect 202782 700788 202788 700800
rect 200080 700760 202788 700788
rect 200080 700748 200086 700760
rect 202782 700748 202788 700760
rect 202840 700748 202846 700800
rect 314470 700748 314476 700800
rect 314528 700788 314534 700800
rect 316310 700788 316316 700800
rect 314528 700760 316316 700788
rect 314528 700748 314534 700760
rect 316310 700748 316316 700760
rect 316368 700748 316374 700800
rect 363506 700408 363512 700460
rect 363564 700448 363570 700460
rect 364978 700448 364984 700460
rect 363564 700420 364984 700448
rect 363564 700408 363570 700420
rect 364978 700408 364984 700420
rect 365036 700408 365042 700460
rect 412450 700408 412456 700460
rect 412508 700448 412514 700460
rect 413646 700448 413652 700460
rect 412508 700420 413652 700448
rect 412508 700408 412514 700420
rect 413646 700408 413652 700420
rect 413704 700408 413710 700460
rect 20346 700204 20352 700256
rect 20404 700244 20410 700256
rect 24302 700244 24308 700256
rect 20404 700216 24308 700244
rect 20404 700204 20410 700216
rect 24302 700204 24308 700216
rect 24360 700204 24366 700256
rect 36722 700204 36728 700256
rect 36780 700244 36786 700256
rect 40494 700244 40500 700256
rect 36780 700216 40500 700244
rect 36780 700204 36786 700216
rect 40494 700204 40500 700216
rect 40552 700204 40558 700256
rect 69382 700204 69388 700256
rect 69440 700244 69446 700256
rect 72970 700244 72976 700256
rect 69440 700216 72976 700244
rect 69440 700204 69446 700216
rect 72970 700204 72976 700216
rect 73028 700204 73034 700256
rect 85758 700204 85764 700256
rect 85816 700244 85822 700256
rect 89162 700244 89168 700256
rect 85816 700216 89168 700244
rect 85816 700204 85822 700216
rect 89162 700204 89168 700216
rect 89220 700204 89226 700256
rect 134702 700204 134708 700256
rect 134760 700244 134766 700256
rect 137830 700244 137836 700256
rect 134760 700216 137836 700244
rect 134760 700204 134766 700216
rect 137830 700204 137836 700216
rect 137888 700204 137894 700256
rect 167362 700204 167368 700256
rect 167420 700244 167426 700256
rect 170306 700244 170312 700256
rect 167420 700216 170312 700244
rect 167420 700204 167426 700216
rect 170306 700204 170312 700216
rect 170364 700204 170370 700256
rect 183738 700204 183744 700256
rect 183796 700244 183802 700256
rect 186498 700244 186504 700256
rect 183796 700216 186504 700244
rect 183796 700204 183802 700216
rect 186498 700204 186504 700216
rect 186556 700204 186562 700256
rect 232774 700204 232780 700256
rect 232832 700244 232838 700256
rect 235166 700244 235172 700256
rect 232832 700216 235172 700244
rect 232832 700204 232838 700216
rect 235166 700204 235172 700216
rect 235224 700204 235230 700256
rect 249058 700204 249064 700256
rect 249116 700244 249122 700256
rect 251450 700244 251456 700256
rect 249116 700216 251456 700244
rect 249116 700204 249122 700216
rect 251450 700204 251456 700216
rect 251508 700204 251514 700256
rect 265434 700204 265440 700256
rect 265492 700244 265498 700256
rect 267642 700244 267648 700256
rect 265492 700216 267648 700244
rect 265492 700204 265498 700216
rect 267642 700204 267648 700216
rect 267700 700204 267706 700256
rect 281810 700204 281816 700256
rect 281868 700244 281874 700256
rect 283834 700244 283840 700256
rect 281868 700216 283840 700244
rect 281868 700204 281874 700216
rect 283834 700204 283840 700216
rect 283892 700204 283898 700256
rect 330754 700204 330760 700256
rect 330812 700244 330818 700256
rect 332502 700244 332508 700256
rect 330812 700216 332508 700244
rect 330812 700204 330818 700216
rect 332502 700204 332508 700216
rect 332560 700204 332566 700256
rect 347130 700204 347136 700256
rect 347188 700244 347194 700256
rect 348786 700244 348792 700256
rect 347188 700216 348792 700244
rect 347188 700204 347194 700216
rect 348786 700204 348792 700216
rect 348844 700204 348850 700256
rect 396166 700204 396172 700256
rect 396224 700244 396230 700256
rect 397454 700244 397460 700256
rect 396224 700216 397460 700244
rect 396224 700204 396230 700216
rect 397454 700204 397460 700216
rect 397512 700204 397518 700256
rect 428826 700204 428832 700256
rect 428884 700244 428890 700256
rect 429838 700244 429844 700256
rect 428884 700216 429844 700244
rect 428884 700204 428890 700216
rect 429838 700204 429844 700216
rect 429896 700204 429902 700256
rect 445202 700204 445208 700256
rect 445260 700244 445266 700256
rect 446122 700244 446128 700256
rect 445260 700216 446128 700244
rect 445260 700204 445266 700216
rect 446122 700204 446128 700216
rect 446180 700204 446186 700256
rect 461486 700204 461492 700256
rect 461544 700244 461550 700256
rect 462314 700244 462320 700256
rect 461544 700216 462320 700244
rect 461544 700204 461550 700216
rect 462314 700204 462320 700216
rect 462372 700204 462378 700256
rect 118418 700136 118424 700188
rect 118476 700176 118482 700188
rect 121638 700176 121644 700188
rect 118476 700148 121644 700176
rect 118476 700136 118482 700148
rect 121638 700136 121644 700148
rect 121696 700136 121702 700188
rect 151078 700136 151084 700188
rect 151136 700176 151142 700188
rect 154114 700176 154120 700188
rect 151136 700148 154120 700176
rect 151136 700136 151142 700148
rect 154114 700136 154120 700148
rect 154172 700136 154178 700188
rect 216398 700136 216404 700188
rect 216456 700176 216462 700188
rect 218974 700176 218980 700188
rect 216456 700148 218980 700176
rect 216456 700136 216462 700148
rect 218974 700136 218980 700148
rect 219032 700136 219038 700188
rect 298002 700136 298008 700188
rect 298060 700176 298066 700188
rect 300118 700176 300124 700188
rect 298060 700148 300124 700176
rect 298060 700136 298066 700148
rect 300118 700136 300124 700148
rect 300176 700136 300182 700188
rect 477862 700136 477868 700188
rect 477920 700176 477926 700188
rect 478506 700176 478512 700188
rect 477920 700148 478512 700176
rect 477920 700136 477926 700148
rect 478506 700136 478512 700148
rect 478564 700136 478570 700188
rect 494238 700136 494244 700188
rect 494296 700176 494302 700188
rect 494790 700176 494796 700188
rect 494296 700148 494796 700176
rect 494296 700136 494302 700148
rect 494790 700136 494796 700148
rect 494848 700136 494854 700188
rect 53006 700000 53012 700052
rect 53064 700040 53070 700052
rect 56778 700040 56784 700052
rect 53064 700012 56784 700040
rect 53064 700000 53070 700012
rect 56778 700000 56784 700012
rect 56836 700000 56842 700052
rect 379790 699864 379796 699916
rect 379848 699904 379854 699916
rect 381170 699904 381176 699916
rect 379848 699876 381176 699904
rect 379848 699864 379854 699876
rect 381170 699864 381176 699876
rect 381228 699864 381234 699916
rect 578326 644512 578332 644564
rect 578384 644552 578390 644564
rect 580902 644552 580908 644564
rect 578384 644524 580908 644552
rect 578384 644512 578390 644524
rect 580902 644512 580908 644524
rect 580960 644512 580966 644564
rect 578878 257796 578884 257848
rect 578936 257836 578942 257848
rect 580902 257836 580908 257848
rect 578936 257808 580908 257836
rect 578936 257796 578942 257808
rect 580902 257796 580908 257808
rect 580960 257796 580966 257848
rect 578510 151444 578516 151496
rect 578568 151484 578574 151496
rect 580902 151484 580908 151496
rect 578568 151456 580908 151484
rect 578568 151444 578574 151456
rect 580902 151444 580908 151456
rect 580960 151444 580966 151496
rect 578326 44956 578332 45008
rect 578384 44996 578390 45008
rect 579982 44996 579988 45008
rect 578384 44968 579988 44996
rect 578384 44956 578390 44968
rect 579982 44956 579988 44968
rect 580040 44956 580046 45008
rect 11146 3884 11152 3936
rect 11204 3924 11210 3936
rect 14502 3924 14508 3936
rect 11204 3896 14508 3924
rect 11204 3884 11210 3896
rect 14502 3884 14508 3896
rect 14560 3884 14566 3936
rect 14734 3884 14740 3936
rect 14792 3924 14798 3936
rect 17998 3924 18004 3936
rect 14792 3896 18004 3924
rect 14792 3884 14798 3896
rect 17998 3884 18004 3896
rect 18056 3884 18062 3936
rect 20622 3884 20628 3936
rect 20680 3924 20686 3936
rect 23794 3924 23800 3936
rect 20680 3896 23800 3924
rect 20680 3884 20686 3896
rect 23794 3884 23800 3896
rect 23852 3884 23858 3936
rect 24210 3884 24216 3936
rect 24268 3924 24274 3936
rect 27290 3924 27296 3936
rect 24268 3896 27296 3924
rect 24268 3884 24274 3896
rect 27290 3884 27296 3896
rect 27348 3884 27354 3936
rect 27706 3884 27712 3936
rect 27764 3924 27770 3936
rect 30694 3924 30700 3936
rect 27764 3896 30700 3924
rect 27764 3884 27770 3896
rect 30694 3884 30700 3896
rect 30752 3884 30758 3936
rect 32398 3884 32404 3936
rect 32456 3924 32462 3936
rect 35386 3924 35392 3936
rect 32456 3896 35392 3924
rect 32456 3884 32462 3896
rect 35386 3884 35392 3896
rect 35444 3884 35450 3936
rect 38378 3884 38384 3936
rect 38436 3924 38442 3936
rect 41182 3924 41188 3936
rect 38436 3896 41188 3924
rect 38436 3884 38442 3896
rect 41182 3884 41188 3896
rect 41240 3884 41246 3936
rect 43070 3884 43076 3936
rect 43128 3924 43134 3936
rect 45782 3924 45788 3936
rect 43128 3896 45788 3924
rect 43128 3884 43134 3896
rect 45782 3884 45788 3896
rect 45840 3884 45846 3936
rect 46658 3884 46664 3936
rect 46716 3924 46722 3936
rect 49278 3924 49284 3936
rect 46716 3896 49284 3924
rect 46716 3884 46722 3896
rect 49278 3884 49284 3896
rect 49336 3884 49342 3936
rect 50154 3884 50160 3936
rect 50212 3924 50218 3936
rect 52774 3924 52780 3936
rect 50212 3896 52780 3924
rect 50212 3884 50218 3896
rect 52774 3884 52780 3896
rect 52832 3884 52838 3936
rect 56042 3884 56048 3936
rect 56100 3924 56106 3936
rect 58570 3924 58576 3936
rect 56100 3896 58576 3924
rect 56100 3884 56106 3896
rect 58570 3884 58576 3896
rect 58628 3884 58634 3936
rect 72602 3884 72608 3936
rect 72660 3924 72666 3936
rect 74854 3924 74860 3936
rect 72660 3896 74860 3924
rect 72660 3884 72666 3896
rect 74854 3884 74860 3896
rect 74912 3884 74918 3936
rect 247630 3884 247636 3936
rect 247688 3924 247694 3936
rect 248598 3924 248604 3936
rect 247688 3896 248604 3924
rect 247688 3884 247694 3896
rect 248598 3884 248604 3896
rect 248656 3884 248662 3936
rect 285902 3884 285908 3936
rect 285960 3924 285966 3936
rect 287790 3924 287796 3936
rect 285960 3896 287796 3924
rect 285960 3884 285966 3896
rect 287790 3884 287796 3896
rect 287848 3884 287854 3936
rect 1670 3816 1676 3868
rect 1728 3856 1734 3868
rect 5210 3856 5216 3868
rect 1728 3828 5216 3856
rect 1728 3816 1734 3828
rect 5210 3816 5216 3828
rect 5268 3816 5274 3868
rect 13538 3816 13544 3868
rect 13596 3856 13602 3868
rect 16802 3856 16808 3868
rect 13596 3828 16808 3856
rect 13596 3816 13602 3828
rect 16802 3816 16808 3828
rect 16860 3816 16866 3868
rect 19426 3816 19432 3868
rect 19484 3856 19490 3868
rect 22598 3856 22604 3868
rect 19484 3828 22604 3856
rect 19484 3816 19490 3828
rect 22598 3816 22604 3828
rect 22656 3816 22662 3868
rect 23014 3816 23020 3868
rect 23072 3856 23078 3868
rect 26094 3856 26100 3868
rect 23072 3828 26100 3856
rect 23072 3816 23078 3828
rect 26094 3816 26100 3828
rect 26152 3816 26158 3868
rect 26510 3816 26516 3868
rect 26568 3856 26574 3868
rect 29590 3856 29596 3868
rect 26568 3828 29596 3856
rect 26568 3816 26574 3828
rect 29590 3816 29596 3828
rect 29648 3816 29654 3868
rect 30098 3816 30104 3868
rect 30156 3856 30162 3868
rect 33086 3856 33092 3868
rect 30156 3828 33092 3856
rect 30156 3816 30162 3828
rect 33086 3816 33092 3828
rect 33144 3816 33150 3868
rect 33594 3816 33600 3868
rect 33652 3856 33658 3868
rect 36582 3856 36588 3868
rect 33652 3828 36588 3856
rect 33652 3816 33658 3828
rect 36582 3816 36588 3828
rect 36640 3816 36646 3868
rect 37182 3816 37188 3868
rect 37240 3856 37246 3868
rect 39986 3856 39992 3868
rect 37240 3828 39992 3856
rect 37240 3816 37246 3828
rect 39986 3816 39992 3828
rect 40044 3816 40050 3868
rect 41874 3816 41880 3868
rect 41932 3856 41938 3868
rect 44678 3856 44684 3868
rect 41932 3828 44684 3856
rect 41932 3816 41938 3828
rect 44678 3816 44684 3828
rect 44736 3816 44742 3868
rect 45462 3816 45468 3868
rect 45520 3856 45526 3868
rect 48174 3856 48180 3868
rect 45520 3828 48180 3856
rect 45520 3816 45526 3828
rect 48174 3816 48180 3828
rect 48232 3816 48238 3868
rect 48958 3816 48964 3868
rect 49016 3856 49022 3868
rect 51578 3856 51584 3868
rect 49016 3828 51584 3856
rect 49016 3816 49022 3828
rect 51578 3816 51584 3828
rect 51636 3816 51642 3868
rect 53742 3816 53748 3868
rect 53800 3856 53806 3868
rect 56270 3856 56276 3868
rect 53800 3828 56276 3856
rect 53800 3816 53806 3828
rect 56270 3816 56276 3828
rect 56328 3816 56334 3868
rect 57238 3816 57244 3868
rect 57296 3856 57302 3868
rect 59766 3856 59772 3868
rect 57296 3828 59772 3856
rect 57296 3816 57302 3828
rect 59766 3816 59772 3828
rect 59824 3816 59830 3868
rect 71498 3816 71504 3868
rect 71556 3856 71562 3868
rect 73658 3856 73664 3868
rect 71556 3828 73664 3856
rect 71556 3816 71562 3828
rect 73658 3816 73664 3828
rect 73716 3816 73722 3868
rect 78582 3816 78588 3868
rect 78640 3856 78646 3868
rect 80650 3856 80656 3868
rect 78640 3828 80656 3856
rect 78640 3816 78646 3828
rect 80650 3816 80656 3828
rect 80708 3816 80714 3868
rect 80882 3816 80888 3868
rect 80940 3856 80946 3868
rect 82950 3856 82956 3868
rect 80940 3828 82956 3856
rect 80940 3816 80946 3828
rect 82950 3816 82956 3828
rect 83008 3816 83014 3868
rect 87966 3816 87972 3868
rect 88024 3856 88030 3868
rect 89942 3856 89948 3868
rect 88024 3828 89948 3856
rect 88024 3816 88030 3828
rect 89942 3816 89948 3828
rect 90000 3816 90006 3868
rect 96246 3816 96252 3868
rect 96304 3856 96310 3868
rect 98038 3856 98044 3868
rect 96304 3828 98044 3856
rect 96304 3816 96310 3828
rect 98038 3816 98044 3828
rect 98096 3816 98102 3868
rect 244134 3816 244140 3868
rect 244192 3856 244198 3868
rect 245194 3856 245200 3868
rect 244192 3828 245200 3856
rect 244192 3816 244198 3828
rect 245194 3816 245200 3828
rect 245252 3816 245258 3868
rect 256922 3816 256928 3868
rect 256980 3856 256986 3868
rect 258258 3856 258264 3868
rect 256980 3828 258264 3856
rect 256980 3816 256986 3828
rect 258258 3816 258264 3828
rect 258316 3816 258322 3868
rect 259222 3816 259228 3868
rect 259280 3856 259286 3868
rect 260650 3856 260656 3868
rect 259280 3828 260656 3856
rect 259280 3816 259286 3828
rect 260650 3816 260656 3828
rect 260708 3816 260714 3868
rect 261614 3816 261620 3868
rect 261672 3856 261678 3868
rect 262950 3856 262956 3868
rect 261672 3828 262956 3856
rect 261672 3816 261678 3828
rect 262950 3816 262956 3828
rect 263008 3816 263014 3868
rect 263914 3816 263920 3868
rect 263972 3856 263978 3868
rect 265342 3856 265348 3868
rect 263972 3828 265348 3856
rect 263972 3816 263978 3828
rect 265342 3816 265348 3828
rect 265400 3816 265406 3868
rect 268514 3816 268520 3868
rect 268572 3856 268578 3868
rect 270034 3856 270040 3868
rect 268572 3828 270040 3856
rect 268572 3816 268578 3828
rect 270034 3816 270040 3828
rect 270092 3816 270098 3868
rect 270814 3816 270820 3868
rect 270872 3856 270878 3868
rect 272426 3856 272432 3868
rect 270872 3828 272432 3856
rect 270872 3816 270878 3828
rect 272426 3816 272432 3828
rect 272484 3816 272490 3868
rect 275506 3816 275512 3868
rect 275564 3856 275570 3868
rect 277118 3856 277124 3868
rect 275564 3828 277124 3856
rect 275564 3816 275570 3828
rect 277118 3816 277124 3828
rect 277176 3816 277182 3868
rect 277806 3816 277812 3868
rect 277864 3856 277870 3868
rect 279510 3856 279516 3868
rect 277864 3828 279516 3856
rect 277864 3816 277870 3828
rect 279510 3816 279516 3828
rect 279568 3816 279574 3868
rect 284798 3816 284804 3868
rect 284856 3856 284862 3868
rect 286594 3856 286600 3868
rect 284856 3828 286600 3856
rect 284856 3816 284862 3828
rect 286594 3816 286600 3828
rect 286652 3816 286658 3868
rect 292894 3816 292900 3868
rect 292952 3856 292958 3868
rect 294874 3856 294880 3868
rect 292952 3828 294880 3856
rect 292952 3816 292958 3828
rect 294874 3816 294880 3828
rect 294932 3816 294938 3868
rect 299886 3816 299892 3868
rect 299944 3856 299950 3868
rect 301958 3856 301964 3868
rect 299944 3828 301964 3856
rect 299944 3816 299950 3828
rect 301958 3816 301964 3828
rect 302016 3816 302022 3868
rect 306786 3816 306792 3868
rect 306844 3856 306850 3868
rect 309042 3856 309048 3868
rect 306844 3828 309048 3856
rect 306844 3816 306850 3828
rect 309042 3816 309048 3828
rect 309100 3816 309106 3868
rect 566 3748 572 3800
rect 624 3788 630 3800
rect 4106 3788 4112 3800
rect 624 3760 4112 3788
rect 624 3748 630 3760
rect 4106 3748 4112 3760
rect 4164 3748 4170 3800
rect 7650 3748 7656 3800
rect 7708 3788 7714 3800
rect 11006 3788 11012 3800
rect 7708 3760 11012 3788
rect 7708 3748 7714 3760
rect 11006 3748 11012 3760
rect 11064 3748 11070 3800
rect 12342 3748 12348 3800
rect 12400 3788 12406 3800
rect 15698 3788 15704 3800
rect 12400 3760 15704 3788
rect 12400 3748 12406 3760
rect 15698 3748 15704 3760
rect 15756 3748 15762 3800
rect 15930 3748 15936 3800
rect 15988 3788 15994 3800
rect 19102 3788 19108 3800
rect 15988 3760 19108 3788
rect 15988 3748 15994 3760
rect 19102 3748 19108 3760
rect 19160 3748 19166 3800
rect 21818 3748 21824 3800
rect 21876 3788 21882 3800
rect 24898 3788 24904 3800
rect 21876 3760 24904 3788
rect 21876 3748 21882 3760
rect 24898 3748 24904 3760
rect 24956 3748 24962 3800
rect 25314 3748 25320 3800
rect 25372 3788 25378 3800
rect 28394 3788 28400 3800
rect 25372 3760 28400 3788
rect 25372 3748 25378 3760
rect 28394 3748 28400 3760
rect 28452 3748 28458 3800
rect 31294 3748 31300 3800
rect 31352 3788 31358 3800
rect 34190 3788 34196 3800
rect 31352 3760 34196 3788
rect 31352 3748 31358 3760
rect 34190 3748 34196 3760
rect 34248 3748 34254 3800
rect 34790 3748 34796 3800
rect 34848 3788 34854 3800
rect 37686 3788 37692 3800
rect 34848 3760 37692 3788
rect 34848 3748 34854 3760
rect 37686 3748 37692 3760
rect 37744 3748 37750 3800
rect 40678 3748 40684 3800
rect 40736 3788 40742 3800
rect 43482 3788 43488 3800
rect 40736 3760 43488 3788
rect 40736 3748 40742 3760
rect 43482 3748 43488 3760
rect 43540 3748 43546 3800
rect 44266 3748 44272 3800
rect 44324 3788 44330 3800
rect 46978 3788 46984 3800
rect 44324 3760 46984 3788
rect 44324 3748 44330 3760
rect 46978 3748 46984 3760
rect 47036 3748 47042 3800
rect 47854 3748 47860 3800
rect 47912 3788 47918 3800
rect 50474 3788 50480 3800
rect 47912 3760 50480 3788
rect 47912 3748 47918 3760
rect 50474 3748 50480 3760
rect 50532 3748 50538 3800
rect 51350 3748 51356 3800
rect 51408 3788 51414 3800
rect 53970 3788 53976 3800
rect 51408 3760 53976 3788
rect 51408 3748 51414 3760
rect 53970 3748 53976 3760
rect 54028 3748 54034 3800
rect 54938 3748 54944 3800
rect 54996 3788 55002 3800
rect 57374 3788 57380 3800
rect 54996 3760 57380 3788
rect 54996 3748 55002 3760
rect 57374 3748 57380 3760
rect 57432 3748 57438 3800
rect 58434 3748 58440 3800
rect 58492 3788 58498 3800
rect 60870 3788 60876 3800
rect 58492 3760 60876 3788
rect 58492 3748 58498 3760
rect 60870 3748 60876 3760
rect 60928 3748 60934 3800
rect 64322 3748 64328 3800
rect 64380 3788 64386 3800
rect 66666 3788 66672 3800
rect 64380 3760 66672 3788
rect 64380 3748 64386 3760
rect 66666 3748 66672 3760
rect 66724 3748 66730 3800
rect 67082 3748 67088 3800
rect 67140 3788 67146 3800
rect 69058 3788 69064 3800
rect 67140 3760 69064 3788
rect 67140 3748 67146 3760
rect 69058 3748 69064 3760
rect 69116 3748 69122 3800
rect 70302 3748 70308 3800
rect 70360 3788 70366 3800
rect 72462 3788 72468 3800
rect 70360 3760 72468 3788
rect 70360 3748 70366 3760
rect 72462 3748 72468 3760
rect 72520 3748 72526 3800
rect 73798 3748 73804 3800
rect 73856 3788 73862 3800
rect 75958 3788 75964 3800
rect 73856 3760 75964 3788
rect 73856 3748 73862 3760
rect 75958 3748 75964 3760
rect 76016 3748 76022 3800
rect 79686 3748 79692 3800
rect 79744 3788 79750 3800
rect 81754 3788 81760 3800
rect 79744 3760 81760 3788
rect 79744 3748 79750 3760
rect 81754 3748 81760 3760
rect 81812 3748 81818 3800
rect 86862 3748 86868 3800
rect 86920 3788 86926 3800
rect 88746 3788 88752 3800
rect 86920 3760 88752 3788
rect 86920 3748 86926 3760
rect 88746 3748 88752 3760
rect 88804 3748 88810 3800
rect 95142 3748 95148 3800
rect 95200 3788 95206 3800
rect 96842 3788 96848 3800
rect 95200 3760 96848 3788
rect 95200 3748 95206 3760
rect 96842 3748 96848 3760
rect 96900 3748 96906 3800
rect 103330 3748 103336 3800
rect 103388 3788 103394 3800
rect 104938 3788 104944 3800
rect 103388 3760 104944 3788
rect 103388 3748 103394 3760
rect 104938 3748 104944 3760
rect 104996 3748 105002 3800
rect 216350 3748 216356 3800
rect 216408 3788 216414 3800
rect 216858 3788 216864 3800
rect 216408 3760 216864 3788
rect 216408 3748 216414 3760
rect 216858 3748 216864 3760
rect 216916 3748 216922 3800
rect 222146 3748 222152 3800
rect 222204 3788 222210 3800
rect 222746 3788 222752 3800
rect 222204 3760 222752 3788
rect 222204 3748 222210 3760
rect 222746 3748 222752 3760
rect 222804 3748 222810 3800
rect 224446 3748 224452 3800
rect 224504 3788 224510 3800
rect 225138 3788 225144 3800
rect 224504 3760 225144 3788
rect 224504 3748 224510 3760
rect 225138 3748 225144 3760
rect 225196 3748 225202 3800
rect 230242 3748 230248 3800
rect 230300 3788 230306 3800
rect 231026 3788 231032 3800
rect 230300 3760 231032 3788
rect 230300 3748 230306 3760
rect 231026 3748 231032 3760
rect 231084 3748 231090 3800
rect 231438 3748 231444 3800
rect 231496 3788 231502 3800
rect 232222 3788 232228 3800
rect 231496 3760 232228 3788
rect 231496 3748 231502 3760
rect 232222 3748 232228 3760
rect 232280 3748 232286 3800
rect 232542 3748 232548 3800
rect 232600 3788 232606 3800
rect 233418 3788 233424 3800
rect 232600 3760 233424 3788
rect 232600 3748 232606 3760
rect 233418 3748 233424 3760
rect 233476 3748 233482 3800
rect 233738 3748 233744 3800
rect 233796 3788 233802 3800
rect 234614 3788 234620 3800
rect 233796 3760 234620 3788
rect 233796 3748 233802 3760
rect 234614 3748 234620 3760
rect 234672 3748 234678 3800
rect 237234 3748 237240 3800
rect 237292 3788 237298 3800
rect 238110 3788 238116 3800
rect 237292 3760 238116 3788
rect 237292 3748 237298 3760
rect 238110 3748 238116 3760
rect 238168 3748 238174 3800
rect 238338 3748 238344 3800
rect 238396 3788 238402 3800
rect 239306 3788 239312 3800
rect 238396 3760 239312 3788
rect 238396 3748 238402 3760
rect 239306 3748 239312 3760
rect 239364 3748 239370 3800
rect 239534 3748 239540 3800
rect 239592 3788 239598 3800
rect 240502 3788 240508 3800
rect 239592 3760 240508 3788
rect 239592 3748 239598 3760
rect 240502 3748 240508 3760
rect 240560 3748 240566 3800
rect 240730 3748 240736 3800
rect 240788 3788 240794 3800
rect 241698 3788 241704 3800
rect 240788 3760 241704 3788
rect 240788 3748 240794 3760
rect 241698 3748 241704 3760
rect 241756 3748 241762 3800
rect 241834 3748 241840 3800
rect 241892 3788 241898 3800
rect 242894 3788 242900 3800
rect 241892 3760 242900 3788
rect 241892 3748 241898 3760
rect 242894 3748 242900 3760
rect 242952 3748 242958 3800
rect 245330 3748 245336 3800
rect 245388 3788 245394 3800
rect 246390 3788 246396 3800
rect 245388 3760 246396 3788
rect 245388 3748 245394 3760
rect 246390 3748 246396 3760
rect 246448 3748 246454 3800
rect 246526 3748 246532 3800
rect 246584 3788 246590 3800
rect 247586 3788 247592 3800
rect 246584 3760 247592 3788
rect 246584 3748 246590 3760
rect 247586 3748 247592 3760
rect 247644 3748 247650 3800
rect 250022 3748 250028 3800
rect 250080 3788 250086 3800
rect 251174 3788 251180 3800
rect 250080 3760 251180 3788
rect 250080 3748 250086 3760
rect 251174 3748 251180 3760
rect 251232 3748 251238 3800
rect 252322 3748 252328 3800
rect 252380 3788 252386 3800
rect 253474 3788 253480 3800
rect 252380 3760 253480 3788
rect 252380 3748 252386 3760
rect 253474 3748 253480 3760
rect 253532 3748 253538 3800
rect 255818 3748 255824 3800
rect 255876 3788 255882 3800
rect 257062 3788 257068 3800
rect 255876 3760 257068 3788
rect 255876 3748 255882 3760
rect 257062 3748 257068 3760
rect 257120 3748 257126 3800
rect 258118 3748 258124 3800
rect 258176 3788 258182 3800
rect 259454 3788 259460 3800
rect 258176 3760 259460 3788
rect 258176 3748 258182 3760
rect 259454 3748 259460 3760
rect 259512 3748 259518 3800
rect 260418 3748 260424 3800
rect 260476 3788 260482 3800
rect 261754 3788 261760 3800
rect 260476 3760 261760 3788
rect 260476 3748 260482 3760
rect 261754 3748 261760 3760
rect 261812 3748 261818 3800
rect 262718 3748 262724 3800
rect 262776 3788 262782 3800
rect 264146 3788 264152 3800
rect 262776 3760 264152 3788
rect 262776 3748 262782 3760
rect 264146 3748 264152 3760
rect 264204 3748 264210 3800
rect 265018 3748 265024 3800
rect 265076 3788 265082 3800
rect 266538 3788 266544 3800
rect 265076 3760 266544 3788
rect 265076 3748 265082 3760
rect 266538 3748 266544 3760
rect 266596 3748 266602 3800
rect 267410 3748 267416 3800
rect 267468 3788 267474 3800
rect 268838 3788 268844 3800
rect 267468 3760 268844 3788
rect 267468 3748 267474 3760
rect 268838 3748 268844 3760
rect 268896 3748 268902 3800
rect 269710 3748 269716 3800
rect 269768 3788 269774 3800
rect 271230 3788 271236 3800
rect 269768 3760 271236 3788
rect 269768 3748 269774 3760
rect 271230 3748 271236 3760
rect 271288 3748 271294 3800
rect 272010 3748 272016 3800
rect 272068 3788 272074 3800
rect 273622 3788 273628 3800
rect 272068 3760 273628 3788
rect 272068 3748 272074 3760
rect 273622 3748 273628 3760
rect 273680 3748 273686 3800
rect 276702 3748 276708 3800
rect 276760 3788 276766 3800
rect 278314 3788 278320 3800
rect 276760 3760 278320 3788
rect 276760 3748 276766 3760
rect 278314 3748 278320 3760
rect 278372 3748 278378 3800
rect 279002 3748 279008 3800
rect 279060 3788 279066 3800
rect 280706 3788 280712 3800
rect 279060 3760 280712 3788
rect 279060 3748 279066 3760
rect 280706 3748 280712 3760
rect 280764 3748 280770 3800
rect 283602 3748 283608 3800
rect 283660 3788 283666 3800
rect 285398 3788 285404 3800
rect 283660 3760 285404 3788
rect 283660 3748 283666 3760
rect 285398 3748 285404 3760
rect 285456 3748 285462 3800
rect 287098 3748 287104 3800
rect 287156 3788 287162 3800
rect 288986 3788 288992 3800
rect 287156 3760 288992 3788
rect 287156 3748 287162 3760
rect 288986 3748 288992 3760
rect 289044 3748 289050 3800
rect 291698 3748 291704 3800
rect 291756 3788 291762 3800
rect 293678 3788 293684 3800
rect 291756 3760 293684 3788
rect 291756 3748 291762 3760
rect 293678 3748 293684 3760
rect 293736 3748 293742 3800
rect 294090 3748 294096 3800
rect 294148 3788 294154 3800
rect 296070 3788 296076 3800
rect 294148 3760 296076 3788
rect 294148 3748 294154 3760
rect 296070 3748 296076 3760
rect 296128 3748 296134 3800
rect 298690 3748 298696 3800
rect 298748 3788 298754 3800
rect 300762 3788 300768 3800
rect 298748 3760 300768 3788
rect 298748 3748 298754 3760
rect 300762 3748 300768 3760
rect 300820 3748 300826 3800
rect 300990 3748 300996 3800
rect 301048 3788 301054 3800
rect 303154 3788 303160 3800
rect 301048 3760 303160 3788
rect 301048 3748 301054 3760
rect 303154 3748 303160 3760
rect 303212 3748 303218 3800
rect 307982 3748 307988 3800
rect 308040 3788 308046 3800
rect 310238 3788 310244 3800
rect 308040 3760 310244 3788
rect 308040 3748 308046 3760
rect 310238 3748 310244 3760
rect 310296 3748 310302 3800
rect 316078 3748 316084 3800
rect 316136 3788 316142 3800
rect 318518 3788 318524 3800
rect 316136 3760 318524 3788
rect 316136 3748 316142 3760
rect 318518 3748 318524 3760
rect 318576 3748 318582 3800
rect 323070 3748 323076 3800
rect 323128 3788 323134 3800
rect 325602 3788 325608 3800
rect 323128 3760 325608 3788
rect 323128 3748 323134 3760
rect 325602 3748 325608 3760
rect 325660 3748 325666 3800
rect 63218 3000 63224 3052
rect 63276 3040 63282 3052
rect 65518 3040 65524 3052
rect 63276 3012 65524 3040
rect 63276 3000 63282 3012
rect 65518 3000 65524 3012
rect 65576 3000 65582 3052
rect 4062 2864 4068 2916
rect 4120 2904 4126 2916
rect 7466 2904 7472 2916
rect 4120 2876 7472 2904
rect 4120 2864 4126 2876
rect 7466 2864 7472 2876
rect 7524 2864 7530 2916
rect 18230 2864 18236 2916
rect 18288 2904 18294 2916
rect 21450 2904 21456 2916
rect 18288 2876 21456 2904
rect 18288 2864 18294 2876
rect 21450 2864 21456 2876
rect 21508 2864 21514 2916
rect 253382 2864 253388 2916
rect 253440 2904 253446 2916
rect 254670 2904 254676 2916
rect 253440 2876 254676 2904
rect 253440 2864 253446 2876
rect 254670 2864 254676 2876
rect 254728 2864 254734 2916
rect 6454 2796 6460 2848
rect 6512 2836 6518 2848
rect 9858 2836 9864 2848
rect 6512 2808 9864 2836
rect 6512 2796 6518 2808
rect 9858 2796 9864 2808
rect 9916 2796 9922 2848
rect 9950 2796 9956 2848
rect 10008 2836 10014 2848
rect 13262 2836 13268 2848
rect 10008 2808 13268 2836
rect 10008 2796 10014 2808
rect 13262 2796 13268 2808
rect 13320 2796 13326 2848
rect 17034 2796 17040 2848
rect 17092 2836 17098 2848
rect 20254 2836 20260 2848
rect 17092 2808 20260 2836
rect 17092 2796 17098 2808
rect 20254 2796 20260 2808
rect 20312 2796 20318 2848
rect 28902 2796 28908 2848
rect 28960 2836 28966 2848
rect 31846 2836 31852 2848
rect 28960 2808 31852 2836
rect 28960 2796 28966 2808
rect 31846 2796 31852 2808
rect 31904 2796 31910 2848
rect 35986 2796 35992 2848
rect 36044 2836 36050 2848
rect 38838 2836 38844 2848
rect 36044 2808 38844 2836
rect 36044 2796 36050 2808
rect 38838 2796 38844 2808
rect 38896 2796 38902 2848
rect 39574 2796 39580 2848
rect 39632 2836 39638 2848
rect 42334 2836 42340 2848
rect 39632 2808 42340 2836
rect 39632 2796 39638 2808
rect 42334 2796 42340 2808
rect 42392 2796 42398 2848
rect 62022 2796 62028 2848
rect 62080 2836 62086 2848
rect 64414 2836 64420 2848
rect 62080 2808 64420 2836
rect 62080 2796 62086 2808
rect 64414 2796 64420 2808
rect 64472 2796 64478 2848
rect 65518 2796 65524 2848
rect 65576 2836 65582 2848
rect 67818 2836 67824 2848
rect 65576 2808 67824 2836
rect 65576 2796 65582 2808
rect 67818 2796 67824 2808
rect 67876 2796 67882 2848
rect 248874 2796 248880 2848
rect 248932 2836 248938 2848
rect 249978 2836 249984 2848
rect 248932 2808 249984 2836
rect 248932 2796 248938 2808
rect 249978 2796 249984 2808
rect 250036 2796 250042 2848
rect 251082 2796 251088 2848
rect 251140 2836 251146 2848
rect 252370 2836 252376 2848
rect 251140 2808 252376 2836
rect 251140 2796 251146 2808
rect 252370 2796 252376 2808
rect 252428 2796 252434 2848
rect 254578 2796 254584 2848
rect 254636 2836 254642 2848
rect 255866 2836 255872 2848
rect 254636 2808 255872 2836
rect 254636 2796 254642 2808
rect 255866 2796 255872 2808
rect 255924 2796 255930 2848
rect 309226 2796 309232 2848
rect 309284 2836 309290 2848
rect 311434 2836 311440 2848
rect 309284 2808 311440 2836
rect 309284 2796 309290 2808
rect 311434 2796 311440 2808
rect 311492 2796 311498 2848
rect 315022 2796 315028 2848
rect 315080 2836 315086 2848
rect 317322 2836 317328 2848
rect 315080 2808 317328 2836
rect 315080 2796 315086 2808
rect 317322 2796 317328 2808
rect 317380 2796 317386 2848
rect 411162 2796 411168 2848
rect 411220 2836 411226 2848
rect 415486 2836 415492 2848
rect 411220 2808 415492 2836
rect 411220 2796 411226 2808
rect 415486 2796 415492 2808
rect 415544 2796 415550 2848
rect 440142 2796 440148 2848
rect 440200 2836 440206 2848
rect 445018 2836 445024 2848
rect 440200 2808 445024 2836
rect 440200 2796 440206 2808
rect 445018 2796 445024 2808
rect 445076 2796 445082 2848
rect 449526 2796 449532 2848
rect 449584 2836 449590 2848
rect 454494 2836 454500 2848
rect 449584 2808 454500 2836
rect 449584 2796 449590 2808
rect 454494 2796 454500 2808
rect 454552 2796 454558 2848
rect 478506 2796 478512 2848
rect 478564 2836 478570 2848
rect 484026 2836 484032 2848
rect 478564 2808 484032 2836
rect 478564 2796 478570 2808
rect 484026 2796 484032 2808
rect 484084 2796 484090 2848
rect 487798 2796 487804 2848
rect 487856 2836 487862 2848
rect 493502 2836 493508 2848
rect 487856 2808 493508 2836
rect 487856 2796 487862 2808
rect 493502 2796 493508 2808
rect 493560 2796 493566 2848
rect 3234 1300 3240 1352
rect 3292 1340 3298 1352
rect 6362 1340 6368 1352
rect 3292 1312 6368 1340
rect 3292 1300 3298 1312
rect 6362 1300 6368 1312
rect 6420 1300 6426 1352
rect 60826 1300 60832 1352
rect 60884 1340 60890 1352
rect 63310 1340 63316 1352
rect 60884 1312 63316 1340
rect 60884 1300 60890 1312
rect 63310 1300 63316 1312
rect 63368 1300 63374 1352
rect 67910 1300 67916 1352
rect 67968 1340 67974 1352
rect 70118 1340 70124 1352
rect 67968 1312 70124 1340
rect 67968 1300 67974 1312
rect 70118 1300 70124 1312
rect 70176 1300 70182 1352
rect 76190 1300 76196 1352
rect 76248 1340 76254 1352
rect 78214 1340 78220 1352
rect 76248 1312 78220 1340
rect 76248 1300 76254 1312
rect 78214 1300 78220 1312
rect 78272 1300 78278 1352
rect 83274 1300 83280 1352
rect 83332 1340 83338 1352
rect 85206 1340 85212 1352
rect 83332 1312 85212 1340
rect 83332 1300 83338 1312
rect 85206 1300 85212 1312
rect 85264 1300 85270 1352
rect 85666 1300 85672 1352
rect 85724 1340 85730 1352
rect 87506 1340 87512 1352
rect 85724 1312 87512 1340
rect 85724 1300 85730 1312
rect 87506 1300 87512 1312
rect 87564 1300 87570 1352
rect 89162 1300 89168 1352
rect 89220 1340 89226 1352
rect 91002 1340 91008 1352
rect 89220 1312 91008 1340
rect 89220 1300 89226 1312
rect 91002 1300 91008 1312
rect 91060 1300 91066 1352
rect 91554 1300 91560 1352
rect 91612 1340 91618 1352
rect 93302 1340 93308 1352
rect 91612 1312 93308 1340
rect 91612 1300 91618 1312
rect 93302 1300 93308 1312
rect 93360 1300 93366 1352
rect 93946 1300 93952 1352
rect 94004 1340 94010 1352
rect 95694 1340 95700 1352
rect 94004 1312 95700 1340
rect 94004 1300 94010 1312
rect 95694 1300 95700 1312
rect 95752 1300 95758 1352
rect 97442 1300 97448 1352
rect 97500 1340 97506 1352
rect 99098 1340 99104 1352
rect 97500 1312 99104 1340
rect 97500 1300 97506 1312
rect 99098 1300 99104 1312
rect 99156 1300 99162 1352
rect 101030 1300 101036 1352
rect 101088 1340 101094 1352
rect 102594 1340 102600 1352
rect 101088 1312 102600 1340
rect 101088 1300 101094 1312
rect 102594 1300 102600 1312
rect 102652 1300 102658 1352
rect 104526 1300 104532 1352
rect 104584 1340 104590 1352
rect 106090 1340 106096 1352
rect 104584 1312 106096 1340
rect 104584 1300 104590 1312
rect 106090 1300 106096 1312
rect 106148 1300 106154 1352
rect 106918 1300 106924 1352
rect 106976 1340 106982 1352
rect 108390 1340 108396 1352
rect 106976 1312 108396 1340
rect 106976 1300 106982 1312
rect 108390 1300 108396 1312
rect 108448 1300 108454 1352
rect 109310 1300 109316 1352
rect 109368 1340 109374 1352
rect 110690 1340 110696 1352
rect 109368 1312 110696 1340
rect 109368 1300 109374 1312
rect 110690 1300 110696 1312
rect 110748 1300 110754 1352
rect 112806 1300 112812 1352
rect 112864 1340 112870 1352
rect 114186 1340 114192 1352
rect 112864 1312 114192 1340
rect 112864 1300 112870 1312
rect 114186 1300 114192 1312
rect 114244 1300 114250 1352
rect 116394 1300 116400 1352
rect 116452 1340 116458 1352
rect 117682 1340 117688 1352
rect 116452 1312 117688 1340
rect 116452 1300 116458 1312
rect 117682 1300 117688 1312
rect 117740 1300 117746 1352
rect 119890 1300 119896 1352
rect 119948 1340 119954 1352
rect 121178 1340 121184 1352
rect 119948 1312 121184 1340
rect 119948 1300 119954 1312
rect 121178 1300 121184 1312
rect 121236 1300 121242 1352
rect 125870 1300 125876 1352
rect 125928 1340 125934 1352
rect 126974 1340 126980 1352
rect 125928 1312 126980 1340
rect 125928 1300 125934 1312
rect 126974 1300 126980 1312
rect 127032 1300 127038 1352
rect 129366 1300 129372 1352
rect 129424 1340 129430 1352
rect 130470 1340 130476 1352
rect 129424 1312 130476 1340
rect 129424 1300 129430 1312
rect 130470 1300 130476 1312
rect 130528 1300 130534 1352
rect 130562 1300 130568 1352
rect 130620 1340 130626 1352
rect 131574 1340 131580 1352
rect 130620 1312 131580 1340
rect 130620 1300 130626 1312
rect 131574 1300 131580 1312
rect 131632 1300 131638 1352
rect 131758 1300 131764 1352
rect 131816 1340 131822 1352
rect 132770 1340 132776 1352
rect 131816 1312 132776 1340
rect 131816 1300 131822 1312
rect 132770 1300 132776 1312
rect 132828 1300 132834 1352
rect 132954 1300 132960 1352
rect 133012 1340 133018 1352
rect 133966 1340 133972 1352
rect 133012 1312 133972 1340
rect 133012 1300 133018 1312
rect 133966 1300 133972 1312
rect 134024 1300 134030 1352
rect 137646 1300 137652 1352
rect 137704 1340 137710 1352
rect 138566 1340 138572 1352
rect 137704 1312 138572 1340
rect 137704 1300 137710 1312
rect 138566 1300 138572 1312
rect 138624 1300 138630 1352
rect 144730 1300 144736 1352
rect 144788 1340 144794 1352
rect 145558 1340 145564 1352
rect 144788 1312 145564 1340
rect 144788 1300 144794 1312
rect 145558 1300 145564 1312
rect 145616 1300 145622 1352
rect 145926 1300 145932 1352
rect 145984 1340 145990 1352
rect 146662 1340 146668 1352
rect 145984 1312 146668 1340
rect 145984 1300 145990 1312
rect 146662 1300 146668 1312
rect 146720 1300 146726 1352
rect 148318 1300 148324 1352
rect 148376 1340 148382 1352
rect 149054 1340 149060 1352
rect 148376 1312 149060 1340
rect 148376 1300 148382 1312
rect 149054 1300 149060 1312
rect 149112 1300 149118 1352
rect 154206 1300 154212 1352
rect 154264 1340 154270 1352
rect 154850 1340 154856 1352
rect 154264 1312 154856 1340
rect 154264 1300 154270 1312
rect 154850 1300 154856 1312
rect 154908 1300 154914 1352
rect 162486 1300 162492 1352
rect 162544 1340 162550 1352
rect 162946 1340 162952 1352
rect 162544 1312 162952 1340
rect 162544 1300 162550 1312
rect 162946 1300 162952 1312
rect 163004 1300 163010 1352
rect 266262 1300 266268 1352
rect 266320 1340 266326 1352
rect 267734 1340 267740 1352
rect 266320 1312 267740 1340
rect 266320 1300 266326 1312
rect 267734 1300 267740 1312
rect 267792 1300 267798 1352
rect 273162 1300 273168 1352
rect 273220 1340 273226 1352
rect 274818 1340 274824 1352
rect 273220 1312 274824 1340
rect 273220 1300 273226 1312
rect 274818 1300 274824 1312
rect 274876 1300 274882 1352
rect 280062 1300 280068 1352
rect 280120 1340 280126 1352
rect 281902 1340 281908 1352
rect 280120 1312 281908 1340
rect 280120 1300 280126 1312
rect 281902 1300 281908 1312
rect 281960 1300 281966 1352
rect 282546 1300 282552 1352
rect 282604 1340 282610 1352
rect 284294 1340 284300 1352
rect 282604 1312 284300 1340
rect 282604 1300 282610 1312
rect 284294 1300 284300 1312
rect 284352 1300 284358 1352
rect 288342 1300 288348 1352
rect 288400 1340 288406 1352
rect 290182 1340 290188 1352
rect 288400 1312 290188 1340
rect 288400 1300 288406 1312
rect 290182 1300 290188 1312
rect 290240 1300 290246 1352
rect 295242 1300 295248 1352
rect 295300 1340 295306 1352
rect 297266 1340 297272 1352
rect 295300 1312 297272 1340
rect 295300 1300 295306 1312
rect 297266 1300 297272 1312
rect 297324 1300 297330 1352
rect 297542 1300 297548 1352
rect 297600 1340 297606 1352
rect 299658 1340 299664 1352
rect 297600 1312 299664 1340
rect 297600 1300 297606 1312
rect 299658 1300 299664 1312
rect 299716 1300 299722 1352
rect 302142 1300 302148 1352
rect 302200 1340 302206 1352
rect 304350 1340 304356 1352
rect 302200 1312 304356 1340
rect 302200 1300 302206 1312
rect 304350 1300 304356 1312
rect 304408 1300 304414 1352
rect 305730 1300 305736 1352
rect 305788 1340 305794 1352
rect 307938 1340 307944 1352
rect 305788 1312 307944 1340
rect 305788 1300 305794 1312
rect 307938 1300 307944 1312
rect 307996 1300 308002 1352
rect 310330 1300 310336 1352
rect 310388 1340 310394 1352
rect 312630 1340 312636 1352
rect 310388 1312 312636 1340
rect 310388 1300 310394 1312
rect 312630 1300 312636 1312
rect 312688 1300 312694 1352
rect 313826 1300 313832 1352
rect 313884 1340 313890 1352
rect 316218 1340 316224 1352
rect 313884 1312 316224 1340
rect 313884 1300 313890 1312
rect 316218 1300 316224 1312
rect 316276 1300 316282 1352
rect 317230 1300 317236 1352
rect 317288 1340 317294 1352
rect 319714 1340 319720 1352
rect 317288 1312 319720 1340
rect 317288 1300 317294 1312
rect 319714 1300 319720 1312
rect 319772 1300 319778 1352
rect 321922 1300 321928 1352
rect 321980 1340 321986 1352
rect 324406 1340 324412 1352
rect 321980 1312 324412 1340
rect 321980 1300 321986 1312
rect 324406 1300 324412 1312
rect 324464 1300 324470 1352
rect 326614 1300 326620 1352
rect 326672 1340 326678 1352
rect 329190 1340 329196 1352
rect 326672 1312 329196 1340
rect 326672 1300 326678 1312
rect 329190 1300 329196 1312
rect 329248 1300 329254 1352
rect 332410 1300 332416 1352
rect 332468 1340 332474 1352
rect 335078 1340 335084 1352
rect 332468 1312 335084 1340
rect 332468 1300 332474 1312
rect 335078 1300 335084 1312
rect 335136 1300 335142 1352
rect 335906 1300 335912 1352
rect 335964 1340 335970 1352
rect 338666 1340 338672 1352
rect 335964 1312 338672 1340
rect 335964 1300 335970 1312
rect 338666 1300 338672 1312
rect 338724 1300 338730 1352
rect 339310 1300 339316 1352
rect 339368 1340 339374 1352
rect 342162 1340 342168 1352
rect 339368 1312 342168 1340
rect 339368 1300 339374 1312
rect 342162 1300 342168 1312
rect 342220 1300 342226 1352
rect 345106 1300 345112 1352
rect 345164 1340 345170 1352
rect 348050 1340 348056 1352
rect 345164 1312 348056 1340
rect 345164 1300 345170 1312
rect 348050 1300 348056 1312
rect 348108 1300 348114 1352
rect 349798 1300 349804 1352
rect 349856 1340 349862 1352
rect 352834 1340 352840 1352
rect 349856 1312 352840 1340
rect 349856 1300 349862 1312
rect 352834 1300 352840 1312
rect 352892 1300 352898 1352
rect 353202 1300 353208 1352
rect 353260 1340 353266 1352
rect 356330 1340 356336 1352
rect 353260 1312 356336 1340
rect 353260 1300 353266 1312
rect 356330 1300 356336 1312
rect 356388 1300 356394 1352
rect 356698 1300 356704 1352
rect 356756 1340 356762 1352
rect 359918 1340 359924 1352
rect 356756 1312 359924 1340
rect 356756 1300 356762 1312
rect 359918 1300 359924 1312
rect 359976 1300 359982 1352
rect 362586 1300 362592 1352
rect 362644 1340 362650 1352
rect 365806 1340 365812 1352
rect 362644 1312 365812 1340
rect 362644 1300 362650 1312
rect 365806 1300 365812 1312
rect 365864 1300 365870 1352
rect 367186 1300 367192 1352
rect 367244 1340 367250 1352
rect 370590 1340 370596 1352
rect 367244 1312 370596 1340
rect 367244 1300 367250 1312
rect 370590 1300 370596 1312
rect 370648 1300 370654 1352
rect 370682 1300 370688 1352
rect 370740 1340 370746 1352
rect 374086 1340 374092 1352
rect 370740 1312 374092 1340
rect 370740 1300 370746 1312
rect 374086 1300 374092 1312
rect 374144 1300 374150 1352
rect 376386 1300 376392 1352
rect 376444 1340 376450 1352
rect 379974 1340 379980 1352
rect 376444 1312 379980 1340
rect 376444 1300 376450 1312
rect 379974 1300 379980 1312
rect 380032 1300 380038 1352
rect 385770 1300 385776 1352
rect 385828 1340 385834 1352
rect 389450 1340 389456 1352
rect 385828 1312 389456 1340
rect 385828 1300 385834 1312
rect 389450 1300 389456 1312
rect 389508 1300 389514 1352
rect 395062 1300 395068 1352
rect 395120 1340 395126 1352
rect 398926 1340 398932 1352
rect 395120 1312 398932 1340
rect 395120 1300 395126 1312
rect 398926 1300 398932 1312
rect 398984 1300 398990 1352
rect 399662 1300 399668 1352
rect 399720 1340 399726 1352
rect 403618 1340 403624 1352
rect 399720 1312 403624 1340
rect 399720 1300 399726 1312
rect 403618 1300 403624 1312
rect 403676 1300 403682 1352
rect 405458 1300 405464 1352
rect 405516 1340 405522 1352
rect 409598 1340 409604 1352
rect 405516 1312 409604 1340
rect 405516 1300 405522 1312
rect 409598 1300 409604 1312
rect 409656 1300 409662 1352
rect 413554 1300 413560 1352
rect 413612 1340 413618 1352
rect 417878 1340 417884 1352
rect 413612 1312 417884 1340
rect 413612 1300 413618 1312
rect 417878 1300 417884 1312
rect 417936 1300 417942 1352
rect 422846 1300 422852 1352
rect 422904 1340 422910 1352
rect 427262 1340 427268 1352
rect 422904 1312 427268 1340
rect 422904 1300 422910 1312
rect 427262 1300 427268 1312
rect 427320 1300 427326 1352
rect 427538 1300 427544 1352
rect 427596 1340 427602 1352
rect 431862 1340 431868 1352
rect 427596 1312 431868 1340
rect 427596 1300 427602 1312
rect 431862 1300 431868 1312
rect 431920 1300 431926 1352
rect 433242 1300 433248 1352
rect 433300 1340 433306 1352
rect 437842 1340 437848 1352
rect 433300 1312 437848 1340
rect 433300 1300 433306 1312
rect 437842 1300 437848 1312
rect 437900 1300 437906 1352
rect 441430 1300 441436 1352
rect 441488 1340 441494 1352
rect 445846 1340 445852 1352
rect 441488 1312 445852 1340
rect 441488 1300 441494 1312
rect 445846 1300 445852 1312
rect 445904 1300 445910 1352
rect 447226 1300 447232 1352
rect 447284 1340 447290 1352
rect 452102 1340 452108 1352
rect 447284 1312 452108 1340
rect 447284 1300 447290 1312
rect 452102 1300 452108 1312
rect 452160 1300 452166 1352
rect 453022 1300 453028 1352
rect 453080 1340 453086 1352
rect 458082 1340 458088 1352
rect 453080 1312 458088 1340
rect 453080 1300 453086 1312
rect 458082 1300 458088 1312
rect 458140 1300 458146 1352
rect 458818 1300 458824 1352
rect 458876 1340 458882 1352
rect 463970 1340 463976 1352
rect 458876 1312 463976 1340
rect 458876 1300 458882 1312
rect 463970 1300 463976 1312
rect 464028 1300 464034 1352
rect 471606 1300 471612 1352
rect 471664 1340 471670 1352
rect 476574 1340 476580 1352
rect 471664 1312 476580 1340
rect 471664 1300 471670 1312
rect 476574 1300 476580 1312
rect 476632 1300 476638 1352
rect 477402 1300 477408 1352
rect 477460 1340 477466 1352
rect 482462 1340 482468 1352
rect 477460 1312 482468 1340
rect 477460 1300 477466 1312
rect 482462 1300 482468 1312
rect 482520 1300 482526 1352
rect 483198 1300 483204 1352
rect 483256 1340 483262 1352
rect 488810 1340 488816 1352
rect 483256 1312 488816 1340
rect 483256 1300 483262 1312
rect 488810 1300 488816 1312
rect 488868 1300 488874 1352
rect 490098 1300 490104 1352
rect 490156 1340 490162 1352
rect 495526 1340 495532 1352
rect 490156 1312 495532 1340
rect 490156 1300 490162 1312
rect 495526 1300 495532 1312
rect 495584 1300 495590 1352
rect 497090 1300 497096 1352
rect 497148 1340 497154 1352
rect 502978 1340 502984 1352
rect 497148 1312 502984 1340
rect 497148 1300 497154 1312
rect 502978 1300 502984 1312
rect 503036 1300 503042 1352
rect 504082 1300 504088 1352
rect 504140 1340 504146 1352
rect 509694 1340 509700 1352
rect 504140 1312 509700 1340
rect 504140 1300 504146 1312
rect 509694 1300 509700 1312
rect 509752 1300 509758 1352
rect 509878 1300 509884 1352
rect 509936 1340 509942 1352
rect 515766 1340 515772 1352
rect 509936 1312 515772 1340
rect 509936 1300 509942 1312
rect 515766 1300 515772 1312
rect 515824 1300 515830 1352
rect 519170 1300 519176 1352
rect 519228 1340 519234 1352
rect 525426 1340 525432 1352
rect 519228 1312 525432 1340
rect 519228 1300 519234 1312
rect 525426 1300 525432 1312
rect 525484 1300 525490 1352
rect 526070 1300 526076 1352
rect 526128 1340 526134 1352
rect 532142 1340 532148 1352
rect 526128 1312 532148 1340
rect 526128 1300 526134 1312
rect 532142 1300 532148 1312
rect 532200 1300 532206 1352
rect 534258 1300 534264 1352
rect 534316 1340 534322 1352
rect 540422 1340 540428 1352
rect 534316 1312 540428 1340
rect 534316 1300 534322 1312
rect 540422 1300 540428 1312
rect 540480 1300 540486 1352
rect 542262 1300 542268 1352
rect 542320 1340 542326 1352
rect 549070 1340 549076 1352
rect 542320 1312 549076 1340
rect 542320 1300 542326 1312
rect 549070 1300 549076 1312
rect 549128 1300 549134 1352
rect 551646 1300 551652 1352
rect 551704 1340 551710 1352
rect 558546 1340 558552 1352
rect 551704 1312 558552 1340
rect 551704 1300 551710 1312
rect 558546 1300 558552 1312
rect 558604 1300 558610 1352
rect 560938 1300 560944 1352
rect 560996 1340 561002 1352
rect 568022 1340 568028 1352
rect 560996 1312 568028 1340
rect 560996 1300 561002 1312
rect 568022 1300 568028 1312
rect 568080 1300 568086 1352
rect 571242 1300 571248 1352
rect 571300 1340 571306 1352
rect 578602 1340 578608 1352
rect 571300 1312 578608 1340
rect 571300 1300 571306 1312
rect 578602 1300 578608 1312
rect 578660 1300 578666 1352
rect 74994 1232 75000 1284
rect 75052 1272 75058 1284
rect 77110 1272 77116 1284
rect 75052 1244 77116 1272
rect 75052 1232 75058 1244
rect 77110 1232 77116 1244
rect 77168 1232 77174 1284
rect 77386 1232 77392 1284
rect 77444 1272 77450 1284
rect 79410 1272 79416 1284
rect 77444 1244 79416 1272
rect 77444 1232 77450 1244
rect 79410 1232 79416 1244
rect 79468 1232 79474 1284
rect 82078 1232 82084 1284
rect 82136 1272 82142 1284
rect 84010 1272 84016 1284
rect 82136 1244 84016 1272
rect 82136 1232 82142 1244
rect 84010 1232 84016 1244
rect 84068 1232 84074 1284
rect 84470 1232 84476 1284
rect 84528 1272 84534 1284
rect 86402 1272 86408 1284
rect 84528 1244 86408 1272
rect 84528 1232 84534 1244
rect 86402 1232 86408 1244
rect 86460 1232 86466 1284
rect 90358 1232 90364 1284
rect 90416 1272 90422 1284
rect 92198 1272 92204 1284
rect 90416 1244 92204 1272
rect 90416 1232 90422 1244
rect 92198 1232 92204 1244
rect 92256 1232 92262 1284
rect 92750 1232 92756 1284
rect 92808 1272 92814 1284
rect 94498 1272 94504 1284
rect 92808 1244 94504 1272
rect 92808 1232 92814 1244
rect 94498 1232 94504 1244
rect 94556 1232 94562 1284
rect 98638 1232 98644 1284
rect 98696 1272 98702 1284
rect 100294 1272 100300 1284
rect 98696 1244 100300 1272
rect 98696 1232 98702 1244
rect 100294 1232 100300 1244
rect 100352 1232 100358 1284
rect 102226 1232 102232 1284
rect 102284 1272 102290 1284
rect 103790 1272 103796 1284
rect 102284 1244 103796 1272
rect 102284 1232 102290 1244
rect 103790 1232 103796 1244
rect 103848 1232 103854 1284
rect 108114 1232 108120 1284
rect 108172 1272 108178 1284
rect 109586 1272 109592 1284
rect 108172 1244 109592 1272
rect 108172 1232 108178 1244
rect 109586 1232 109592 1244
rect 109644 1232 109650 1284
rect 110506 1232 110512 1284
rect 110564 1272 110570 1284
rect 111886 1272 111892 1284
rect 110564 1244 111892 1272
rect 110564 1232 110570 1244
rect 111886 1232 111892 1244
rect 111944 1232 111950 1284
rect 115198 1232 115204 1284
rect 115256 1272 115262 1284
rect 116578 1272 116584 1284
rect 115256 1244 116584 1272
rect 115256 1232 115262 1244
rect 116578 1232 116584 1244
rect 116636 1232 116642 1284
rect 117590 1232 117596 1284
rect 117648 1272 117654 1284
rect 118878 1272 118884 1284
rect 117648 1244 118884 1272
rect 117648 1232 117654 1244
rect 118878 1232 118884 1244
rect 118936 1232 118942 1284
rect 122282 1232 122288 1284
rect 122340 1272 122346 1284
rect 123478 1272 123484 1284
rect 122340 1244 123484 1272
rect 122340 1232 122346 1244
rect 123478 1232 123484 1244
rect 123536 1232 123542 1284
rect 124674 1232 124680 1284
rect 124732 1272 124738 1284
rect 125778 1272 125784 1284
rect 124732 1244 125784 1272
rect 124732 1232 124738 1244
rect 125778 1232 125784 1244
rect 125836 1232 125842 1284
rect 128170 1232 128176 1284
rect 128228 1272 128234 1284
rect 129274 1272 129280 1284
rect 128228 1244 129280 1272
rect 128228 1232 128234 1244
rect 129274 1232 129280 1244
rect 129332 1232 129338 1284
rect 136450 1232 136456 1284
rect 136508 1272 136514 1284
rect 137370 1272 137376 1284
rect 136508 1244 137376 1272
rect 136508 1232 136514 1244
rect 137370 1232 137376 1244
rect 137428 1232 137434 1284
rect 138842 1232 138848 1284
rect 138900 1272 138906 1284
rect 139762 1272 139768 1284
rect 138900 1244 139768 1272
rect 138900 1232 138906 1244
rect 139762 1232 139768 1244
rect 139820 1232 139826 1284
rect 140038 1232 140044 1284
rect 140096 1272 140102 1284
rect 140866 1272 140872 1284
rect 140096 1244 140872 1272
rect 140096 1232 140102 1244
rect 140866 1232 140872 1244
rect 140924 1232 140930 1284
rect 281350 1232 281356 1284
rect 281408 1272 281414 1284
rect 283098 1272 283104 1284
rect 281408 1244 283104 1272
rect 281408 1232 281414 1244
rect 283098 1232 283104 1244
rect 283156 1232 283162 1284
rect 289446 1232 289452 1284
rect 289504 1272 289510 1284
rect 291378 1272 291384 1284
rect 289504 1244 291384 1272
rect 289504 1232 289510 1244
rect 291378 1232 291384 1244
rect 291436 1232 291442 1284
rect 296438 1232 296444 1284
rect 296496 1272 296502 1284
rect 298462 1272 298468 1284
rect 296496 1244 298468 1272
rect 296496 1232 296502 1244
rect 298462 1232 298468 1244
rect 298520 1232 298526 1284
rect 303338 1232 303344 1284
rect 303396 1272 303402 1284
rect 305546 1272 305552 1284
rect 303396 1244 305552 1272
rect 303396 1232 303402 1244
rect 305546 1232 305552 1244
rect 305604 1232 305610 1284
rect 312538 1232 312544 1284
rect 312596 1272 312602 1284
rect 315022 1272 315028 1284
rect 312596 1244 315028 1272
rect 312596 1232 312602 1244
rect 315022 1232 315028 1244
rect 315080 1232 315086 1284
rect 318426 1232 318432 1284
rect 318484 1272 318490 1284
rect 320910 1272 320916 1284
rect 318484 1244 320916 1272
rect 318484 1232 318490 1244
rect 320910 1232 320916 1244
rect 320968 1232 320974 1284
rect 328914 1232 328920 1284
rect 328972 1272 328978 1284
rect 331582 1272 331588 1284
rect 328972 1244 331588 1272
rect 328972 1232 328978 1244
rect 331582 1232 331588 1244
rect 331640 1232 331646 1284
rect 334710 1232 334716 1284
rect 334768 1272 334774 1284
rect 337470 1272 337476 1284
rect 334768 1244 337476 1272
rect 334768 1232 334774 1244
rect 337470 1232 337476 1244
rect 337528 1232 337534 1284
rect 340506 1232 340512 1284
rect 340564 1272 340570 1284
rect 343358 1272 343364 1284
rect 340564 1244 343364 1272
rect 340564 1232 340570 1244
rect 343358 1232 343364 1244
rect 343416 1232 343422 1284
rect 344002 1232 344008 1284
rect 344060 1272 344066 1284
rect 346946 1272 346952 1284
rect 344060 1244 346952 1272
rect 344060 1232 344066 1244
rect 346946 1232 346952 1244
rect 347004 1232 347010 1284
rect 348602 1232 348608 1284
rect 348660 1272 348666 1284
rect 351638 1272 351644 1284
rect 348660 1244 351644 1272
rect 348660 1232 348666 1244
rect 351638 1232 351644 1244
rect 351696 1232 351702 1284
rect 352098 1232 352104 1284
rect 352156 1272 352162 1284
rect 355226 1272 355232 1284
rect 352156 1244 355232 1272
rect 352156 1232 352162 1244
rect 355226 1232 355232 1244
rect 355284 1232 355290 1284
rect 355594 1232 355600 1284
rect 355652 1272 355658 1284
rect 358722 1272 358728 1284
rect 355652 1244 358728 1272
rect 355652 1232 355658 1244
rect 358722 1232 358728 1244
rect 358780 1232 358786 1284
rect 359090 1232 359096 1284
rect 359148 1272 359154 1284
rect 362310 1272 362316 1284
rect 359148 1244 362316 1272
rect 359148 1232 359154 1244
rect 362310 1232 362316 1244
rect 362368 1232 362374 1284
rect 363690 1232 363696 1284
rect 363748 1272 363754 1284
rect 367002 1272 367008 1284
rect 363748 1244 367008 1272
rect 363748 1232 363754 1244
rect 367002 1232 367008 1244
rect 367060 1232 367066 1284
rect 372982 1232 372988 1284
rect 373040 1272 373046 1284
rect 376478 1272 376484 1284
rect 373040 1244 376484 1272
rect 373040 1232 373046 1244
rect 376478 1232 376484 1244
rect 376536 1232 376542 1284
rect 377582 1232 377588 1284
rect 377640 1272 377646 1284
rect 381170 1272 381176 1284
rect 377640 1244 381176 1272
rect 377640 1232 377646 1244
rect 381170 1232 381176 1244
rect 381228 1232 381234 1284
rect 388070 1232 388076 1284
rect 388128 1272 388134 1284
rect 391842 1272 391848 1284
rect 388128 1244 391848 1272
rect 388128 1232 388134 1244
rect 391842 1232 391848 1244
rect 391900 1232 391906 1284
rect 393866 1232 393872 1284
rect 393924 1272 393930 1284
rect 397730 1272 397736 1284
rect 393924 1244 397736 1272
rect 393924 1232 393930 1244
rect 397730 1232 397736 1244
rect 397788 1232 397794 1284
rect 403158 1232 403164 1284
rect 403216 1272 403222 1284
rect 407206 1272 407212 1284
rect 403216 1244 407212 1272
rect 403216 1232 403222 1244
rect 407206 1232 407212 1244
rect 407264 1232 407270 1284
rect 410058 1232 410064 1284
rect 410116 1272 410122 1284
rect 414290 1272 414296 1284
rect 410116 1244 414296 1272
rect 410116 1232 410122 1244
rect 414290 1232 414296 1244
rect 414348 1232 414354 1284
rect 418246 1232 418252 1284
rect 418304 1272 418310 1284
rect 422570 1272 422576 1284
rect 418304 1244 422576 1272
rect 418304 1232 418310 1244
rect 422570 1232 422576 1244
rect 422628 1232 422634 1284
rect 426342 1232 426348 1284
rect 426400 1272 426406 1284
rect 430850 1272 430856 1284
rect 426400 1244 430856 1272
rect 426400 1232 426406 1244
rect 430850 1232 430856 1244
rect 430908 1232 430914 1284
rect 435634 1232 435640 1284
rect 435692 1272 435698 1284
rect 439958 1272 439964 1284
rect 435692 1244 439964 1272
rect 435692 1232 435698 1244
rect 439958 1232 439964 1244
rect 440016 1232 440022 1284
rect 442626 1232 442632 1284
rect 442684 1272 442690 1284
rect 447410 1272 447416 1284
rect 442684 1244 447416 1272
rect 442684 1232 442690 1244
rect 447410 1232 447416 1244
rect 447468 1232 447474 1284
rect 457622 1232 457628 1284
rect 457680 1272 457686 1284
rect 462406 1272 462412 1284
rect 457680 1244 462412 1272
rect 457680 1232 457686 1244
rect 462406 1232 462412 1244
rect 462464 1232 462470 1284
rect 468110 1232 468116 1284
rect 468168 1272 468174 1284
rect 473078 1272 473084 1284
rect 468168 1244 473084 1272
rect 468168 1232 468174 1244
rect 473078 1232 473084 1244
rect 473136 1232 473142 1284
rect 475102 1232 475108 1284
rect 475160 1272 475166 1284
rect 480530 1272 480536 1284
rect 475160 1244 480536 1272
rect 475160 1232 475166 1244
rect 480530 1232 480536 1244
rect 480588 1232 480594 1284
rect 485498 1232 485504 1284
rect 485556 1272 485562 1284
rect 490742 1272 490748 1284
rect 485556 1244 490748 1272
rect 485556 1232 485562 1244
rect 490742 1232 490748 1244
rect 490800 1232 490806 1284
rect 492490 1232 492496 1284
rect 492548 1272 492554 1284
rect 498194 1272 498200 1284
rect 492548 1244 498200 1272
rect 492548 1232 492554 1244
rect 498194 1232 498200 1244
rect 498252 1232 498258 1284
rect 498286 1232 498292 1284
rect 498344 1272 498350 1284
rect 503806 1272 503812 1284
rect 498344 1244 503812 1272
rect 498344 1232 498350 1244
rect 503806 1232 503812 1244
rect 503864 1232 503870 1284
rect 510982 1232 510988 1284
rect 511040 1272 511046 1284
rect 517146 1272 517152 1284
rect 511040 1244 517152 1272
rect 511040 1232 511046 1244
rect 517146 1232 517152 1244
rect 517204 1232 517210 1284
rect 517974 1232 517980 1284
rect 518032 1272 518038 1284
rect 523862 1272 523868 1284
rect 518032 1244 523868 1272
rect 518032 1232 518038 1244
rect 523862 1232 523868 1244
rect 523920 1232 523926 1284
rect 527266 1232 527272 1284
rect 527324 1272 527330 1284
rect 533706 1272 533712 1284
rect 527324 1244 533712 1272
rect 527324 1232 527330 1244
rect 533706 1232 533712 1244
rect 533764 1232 533770 1284
rect 541158 1232 541164 1284
rect 541216 1272 541222 1284
rect 547874 1272 547880 1284
rect 541216 1244 547880 1272
rect 541216 1232 541222 1244
rect 547874 1232 547880 1244
rect 547932 1232 547938 1284
rect 548150 1232 548156 1284
rect 548208 1272 548214 1284
rect 554958 1272 554964 1284
rect 548208 1244 554964 1272
rect 548208 1232 548214 1244
rect 554958 1232 554964 1244
rect 555016 1232 555022 1284
rect 562042 1232 562048 1284
rect 562100 1272 562106 1284
rect 569126 1272 569132 1284
rect 562100 1244 569132 1272
rect 562100 1232 562106 1244
rect 569126 1232 569132 1244
rect 569184 1232 569190 1284
rect 570138 1232 570144 1284
rect 570196 1272 570202 1284
rect 577406 1272 577412 1284
rect 570196 1244 577412 1272
rect 570196 1232 570202 1244
rect 577406 1232 577412 1244
rect 577464 1232 577470 1284
rect 99834 1164 99840 1216
rect 99892 1204 99898 1216
rect 101490 1204 101496 1216
rect 99892 1176 101496 1204
rect 99892 1164 99898 1176
rect 101490 1164 101496 1176
rect 101548 1164 101554 1216
rect 114002 1164 114008 1216
rect 114060 1204 114066 1216
rect 115382 1204 115388 1216
rect 114060 1176 115388 1204
rect 114060 1164 114066 1176
rect 115382 1164 115388 1176
rect 115440 1164 115446 1216
rect 311526 1164 311532 1216
rect 311584 1204 311590 1216
rect 313826 1204 313832 1216
rect 311584 1176 313832 1204
rect 311584 1164 311590 1176
rect 313826 1164 313832 1176
rect 313884 1164 313890 1216
rect 319622 1164 319628 1216
rect 319680 1204 319686 1216
rect 322106 1204 322112 1216
rect 319680 1176 322112 1204
rect 319680 1164 319686 1176
rect 322106 1164 322112 1176
rect 322164 1164 322170 1216
rect 330018 1164 330024 1216
rect 330076 1204 330082 1216
rect 332686 1204 332692 1216
rect 330076 1176 332692 1204
rect 330076 1164 330082 1176
rect 332686 1164 332692 1176
rect 332744 1164 332750 1216
rect 337010 1164 337016 1216
rect 337068 1204 337074 1216
rect 339862 1204 339868 1216
rect 337068 1176 339868 1204
rect 337068 1164 337074 1176
rect 339862 1164 339868 1176
rect 339920 1164 339926 1216
rect 341702 1164 341708 1216
rect 341760 1204 341766 1216
rect 344554 1204 344560 1216
rect 341760 1176 344560 1204
rect 341760 1164 341766 1176
rect 344554 1164 344560 1176
rect 344612 1164 344618 1216
rect 357894 1164 357900 1216
rect 357952 1204 357958 1216
rect 361114 1204 361120 1216
rect 357952 1176 361120 1204
rect 357952 1164 357958 1176
rect 361114 1164 361120 1176
rect 361172 1164 361178 1216
rect 364886 1164 364892 1216
rect 364944 1204 364950 1216
rect 368198 1204 368204 1216
rect 364944 1176 368204 1204
rect 364944 1164 364950 1176
rect 368198 1164 368204 1176
rect 368256 1164 368262 1216
rect 375282 1164 375288 1216
rect 375340 1204 375346 1216
rect 378870 1204 378876 1216
rect 375340 1176 378876 1204
rect 375340 1164 375346 1176
rect 378870 1164 378876 1176
rect 378928 1164 378934 1216
rect 381078 1164 381084 1216
rect 381136 1204 381142 1216
rect 384758 1204 384764 1216
rect 381136 1176 384764 1204
rect 381136 1164 381142 1176
rect 384758 1164 384764 1176
rect 384816 1164 384822 1216
rect 390370 1164 390376 1216
rect 390428 1204 390434 1216
rect 394234 1204 394240 1216
rect 390428 1176 394240 1204
rect 390428 1164 390434 1176
rect 394234 1164 394240 1176
rect 394292 1164 394298 1216
rect 396166 1164 396172 1216
rect 396224 1204 396230 1216
rect 400122 1204 400128 1216
rect 396224 1176 400128 1204
rect 396224 1164 396230 1176
rect 400122 1164 400128 1176
rect 400180 1164 400186 1216
rect 400858 1164 400864 1216
rect 400916 1204 400922 1216
rect 404814 1204 404820 1216
rect 400916 1176 404820 1204
rect 400916 1164 400922 1176
rect 404814 1164 404820 1176
rect 404872 1164 404878 1216
rect 407758 1164 407764 1216
rect 407816 1204 407822 1216
rect 411898 1204 411904 1216
rect 407816 1176 411904 1204
rect 407816 1164 407822 1176
rect 411898 1164 411904 1176
rect 411956 1164 411962 1216
rect 420546 1164 420552 1216
rect 420604 1204 420610 1216
rect 424962 1204 424968 1216
rect 420604 1176 424968 1204
rect 420604 1164 420610 1176
rect 424962 1164 424968 1176
rect 425020 1164 425026 1216
rect 425146 1164 425152 1216
rect 425204 1204 425210 1216
rect 429654 1204 429660 1216
rect 425204 1176 429660 1204
rect 425204 1164 425210 1176
rect 429654 1164 429660 1176
rect 429712 1164 429718 1216
rect 436738 1164 436744 1216
rect 436796 1204 436802 1216
rect 441522 1204 441528 1216
rect 436796 1176 441528 1204
rect 436796 1164 436802 1176
rect 441522 1164 441528 1176
rect 441580 1164 441586 1216
rect 444926 1164 444932 1216
rect 444984 1204 444990 1216
rect 449802 1204 449808 1216
rect 444984 1176 449808 1204
rect 444984 1164 444990 1176
rect 449802 1164 449808 1176
rect 449860 1164 449866 1216
rect 450722 1164 450728 1216
rect 450780 1204 450786 1216
rect 455690 1204 455696 1216
rect 450780 1176 455696 1204
rect 450780 1164 450786 1176
rect 455690 1164 455696 1176
rect 455748 1164 455754 1216
rect 456518 1164 456524 1216
rect 456576 1204 456582 1216
rect 461578 1204 461584 1216
rect 456576 1176 461584 1204
rect 456576 1164 456582 1176
rect 461578 1164 461584 1176
rect 461636 1164 461642 1216
rect 462222 1164 462228 1216
rect 462280 1204 462286 1216
rect 467466 1204 467472 1216
rect 462280 1176 467472 1204
rect 462280 1164 462286 1176
rect 467466 1164 467472 1176
rect 467524 1164 467530 1216
rect 472710 1164 472716 1216
rect 472768 1204 472774 1216
rect 478138 1204 478144 1216
rect 472768 1176 478144 1204
rect 472768 1164 472774 1176
rect 478138 1164 478144 1176
rect 478196 1164 478202 1216
rect 480898 1164 480904 1216
rect 480956 1204 480962 1216
rect 486418 1204 486424 1216
rect 480956 1176 486424 1204
rect 480956 1164 480962 1176
rect 486418 1164 486424 1176
rect 486476 1164 486482 1216
rect 486694 1164 486700 1216
rect 486752 1204 486758 1216
rect 492306 1204 492312 1216
rect 486752 1176 492312 1204
rect 486752 1164 486758 1176
rect 492306 1164 492312 1176
rect 492364 1164 492370 1216
rect 493594 1164 493600 1216
rect 493652 1204 493658 1216
rect 499390 1204 499396 1216
rect 493652 1176 499396 1204
rect 493652 1164 493658 1176
rect 499390 1164 499396 1176
rect 499448 1164 499454 1216
rect 500586 1164 500592 1216
rect 500644 1204 500650 1216
rect 506474 1204 506480 1216
rect 500644 1176 506480 1204
rect 500644 1164 500650 1176
rect 506474 1164 506480 1176
rect 506532 1164 506538 1216
rect 522666 1164 522672 1216
rect 522724 1204 522730 1216
rect 529014 1204 529020 1216
rect 522724 1176 529020 1204
rect 522724 1164 522730 1176
rect 529014 1164 529020 1176
rect 529072 1164 529078 1216
rect 530762 1164 530768 1216
rect 530820 1204 530826 1216
rect 537202 1204 537208 1216
rect 530820 1176 537208 1204
rect 530820 1164 530826 1176
rect 537202 1164 537208 1176
rect 537260 1164 537266 1216
rect 538858 1164 538864 1216
rect 538916 1204 538922 1216
rect 545482 1204 545488 1216
rect 538916 1176 545488 1204
rect 538916 1164 538922 1176
rect 545482 1164 545488 1176
rect 545540 1164 545546 1216
rect 550450 1164 550456 1216
rect 550508 1204 550514 1216
rect 557350 1204 557356 1216
rect 550508 1176 557356 1204
rect 550508 1164 550514 1176
rect 557350 1164 557356 1176
rect 557408 1164 557414 1216
rect 558454 1164 558460 1216
rect 558512 1204 558518 1216
rect 565630 1204 565636 1216
rect 558512 1176 565636 1204
rect 558512 1164 558518 1176
rect 565630 1164 565636 1176
rect 565688 1164 565694 1216
rect 569034 1164 569040 1216
rect 569092 1204 569098 1216
rect 576302 1204 576308 1216
rect 569092 1176 576308 1204
rect 569092 1164 569098 1176
rect 576302 1164 576308 1176
rect 576360 1164 576366 1216
rect 5626 1096 5632 1148
rect 5684 1136 5690 1148
rect 8662 1136 8668 1148
rect 5684 1108 8668 1136
rect 5684 1096 5690 1108
rect 8662 1096 8668 1108
rect 8720 1096 8726 1148
rect 111610 1096 111616 1148
rect 111668 1136 111674 1148
rect 113082 1136 113088 1148
rect 111668 1108 113088 1136
rect 111668 1096 111674 1108
rect 113082 1096 113088 1108
rect 113140 1096 113146 1148
rect 123478 1096 123484 1148
rect 123536 1136 123542 1148
rect 124766 1136 124772 1148
rect 123536 1108 124772 1136
rect 123536 1096 123542 1108
rect 124766 1096 124772 1108
rect 124824 1096 124830 1148
rect 320818 1096 320824 1148
rect 320876 1136 320882 1148
rect 323302 1136 323308 1148
rect 320876 1108 323308 1136
rect 320876 1096 320882 1108
rect 323302 1096 323308 1108
rect 323360 1096 323366 1148
rect 331122 1096 331128 1148
rect 331180 1136 331186 1148
rect 333882 1136 333888 1148
rect 331180 1108 333888 1136
rect 331180 1096 331186 1108
rect 333882 1096 333888 1108
rect 333940 1096 333946 1148
rect 360102 1096 360108 1148
rect 360160 1136 360166 1148
rect 363506 1136 363512 1148
rect 360160 1108 363512 1136
rect 360160 1096 360166 1108
rect 363506 1096 363512 1108
rect 363564 1096 363570 1148
rect 382182 1096 382188 1148
rect 382240 1136 382246 1148
rect 385954 1136 385960 1148
rect 382240 1108 385960 1136
rect 382240 1096 382246 1108
rect 385954 1096 385960 1108
rect 386012 1096 386018 1148
rect 389266 1096 389272 1148
rect 389324 1136 389330 1148
rect 393038 1136 393044 1148
rect 389324 1108 393044 1136
rect 389324 1096 389330 1108
rect 393038 1096 393044 1108
rect 393096 1096 393102 1148
rect 398466 1096 398472 1148
rect 398524 1136 398530 1148
rect 402514 1136 402520 1148
rect 398524 1108 402520 1136
rect 398524 1096 398530 1108
rect 402514 1096 402520 1108
rect 402572 1096 402578 1148
rect 404262 1096 404268 1148
rect 404320 1136 404326 1148
rect 408402 1136 408408 1148
rect 404320 1108 408408 1136
rect 404320 1096 404326 1108
rect 408402 1096 408408 1108
rect 408460 1096 408466 1148
rect 408954 1096 408960 1148
rect 409012 1136 409018 1148
rect 413094 1136 413100 1148
rect 409012 1108 413100 1136
rect 409012 1096 409018 1108
rect 413094 1096 413100 1108
rect 413152 1096 413158 1148
rect 415946 1096 415952 1148
rect 416004 1136 416010 1148
rect 420178 1136 420184 1148
rect 416004 1108 420184 1136
rect 416004 1096 416010 1108
rect 420178 1096 420184 1108
rect 420236 1096 420242 1148
rect 428642 1096 428648 1148
rect 428700 1136 428706 1148
rect 433242 1136 433248 1148
rect 428700 1108 433248 1136
rect 428700 1096 428706 1108
rect 433242 1096 433248 1108
rect 433300 1096 433306 1148
rect 439130 1096 439136 1148
rect 439188 1136 439194 1148
rect 443822 1136 443828 1148
rect 439188 1108 443828 1136
rect 439188 1096 439194 1108
rect 443822 1096 443828 1108
rect 443880 1096 443886 1148
rect 448422 1096 448428 1148
rect 448480 1136 448486 1148
rect 453298 1136 453304 1148
rect 448480 1108 453304 1136
rect 448480 1096 448486 1108
rect 453298 1096 453304 1108
rect 453356 1096 453362 1148
rect 454218 1096 454224 1148
rect 454276 1136 454282 1148
rect 459186 1136 459192 1148
rect 454276 1108 459192 1136
rect 454276 1096 454282 1108
rect 459186 1096 459192 1108
rect 459244 1096 459250 1148
rect 465810 1096 465816 1148
rect 465868 1136 465874 1148
rect 470686 1136 470692 1148
rect 465868 1108 470692 1136
rect 465868 1096 465874 1108
rect 470686 1096 470692 1108
rect 470744 1096 470750 1148
rect 482002 1096 482008 1148
rect 482060 1136 482066 1148
rect 487246 1136 487252 1148
rect 482060 1108 487252 1136
rect 482060 1096 482066 1108
rect 487246 1096 487252 1108
rect 487304 1096 487310 1148
rect 488994 1096 489000 1148
rect 489052 1136 489058 1148
rect 494698 1136 494704 1148
rect 489052 1108 494704 1136
rect 489052 1096 489058 1108
rect 494698 1096 494704 1108
rect 494756 1096 494762 1148
rect 501782 1096 501788 1148
rect 501840 1136 501846 1148
rect 507302 1136 507308 1148
rect 501840 1108 507308 1136
rect 501840 1096 501846 1108
rect 507302 1096 507308 1108
rect 507360 1096 507366 1148
rect 513282 1096 513288 1148
rect 513340 1136 513346 1148
rect 519538 1136 519544 1148
rect 513340 1108 519544 1136
rect 513340 1096 513346 1108
rect 519538 1096 519544 1108
rect 519596 1096 519602 1148
rect 523770 1096 523776 1148
rect 523828 1136 523834 1148
rect 530118 1136 530124 1148
rect 523828 1108 530124 1136
rect 523828 1096 523834 1108
rect 530118 1096 530124 1108
rect 530176 1096 530182 1148
rect 533062 1096 533068 1148
rect 533120 1136 533126 1148
rect 539594 1136 539600 1148
rect 533120 1108 539600 1136
rect 533120 1096 533126 1108
rect 539594 1096 539600 1108
rect 539652 1096 539658 1148
rect 543458 1096 543464 1148
rect 543516 1136 543522 1148
rect 550266 1136 550272 1148
rect 543516 1108 550272 1136
rect 543516 1096 543522 1108
rect 550266 1096 550272 1108
rect 550324 1096 550330 1148
rect 552750 1096 552756 1148
rect 552808 1136 552814 1148
rect 559742 1136 559748 1148
rect 552808 1108 559748 1136
rect 552808 1096 552814 1108
rect 559742 1096 559748 1108
rect 559800 1096 559806 1148
rect 567838 1096 567844 1148
rect 567896 1136 567902 1148
rect 575106 1136 575112 1148
rect 567896 1108 575112 1136
rect 567896 1096 567902 1108
rect 575106 1096 575112 1108
rect 575164 1096 575170 1148
rect 378778 1028 378784 1080
rect 378836 1068 378842 1080
rect 382366 1068 382372 1080
rect 378836 1040 382372 1068
rect 378836 1028 378842 1040
rect 382366 1028 382372 1040
rect 382424 1028 382430 1080
rect 386874 1028 386880 1080
rect 386932 1068 386938 1080
rect 390646 1068 390652 1080
rect 386932 1040 390652 1068
rect 386932 1028 386938 1040
rect 390646 1028 390652 1040
rect 390704 1028 390710 1080
rect 417050 1028 417056 1080
rect 417108 1068 417114 1080
rect 421374 1068 421380 1080
rect 417108 1040 421380 1068
rect 417108 1028 417114 1040
rect 421374 1028 421380 1040
rect 421432 1028 421438 1080
rect 437934 1028 437940 1080
rect 437992 1068 437998 1080
rect 442626 1068 442632 1080
rect 437992 1040 442632 1068
rect 437992 1028 437998 1040
rect 442626 1028 442632 1040
rect 442684 1028 442690 1080
rect 446030 1028 446036 1080
rect 446088 1068 446094 1080
rect 450906 1068 450912 1080
rect 446088 1040 450912 1068
rect 446088 1028 446094 1040
rect 450906 1028 450912 1040
rect 450964 1028 450970 1080
rect 455322 1028 455328 1080
rect 455380 1068 455386 1080
rect 460106 1068 460112 1080
rect 455380 1040 460112 1068
rect 455380 1028 455386 1040
rect 460106 1028 460112 1040
rect 460164 1028 460170 1080
rect 461118 1028 461124 1080
rect 461176 1068 461182 1080
rect 466270 1068 466276 1080
rect 461176 1040 466276 1068
rect 461176 1028 461182 1040
rect 466270 1028 466276 1040
rect 466328 1028 466334 1080
rect 466914 1028 466920 1080
rect 466972 1068 466978 1080
rect 472250 1068 472256 1080
rect 466972 1040 472256 1068
rect 466972 1028 466978 1040
rect 472250 1028 472256 1040
rect 472308 1028 472314 1080
rect 479702 1028 479708 1080
rect 479760 1068 479766 1080
rect 484854 1068 484860 1080
rect 479760 1040 484860 1068
rect 479760 1028 479766 1040
rect 484854 1028 484860 1040
rect 484912 1028 484918 1080
rect 491202 1028 491208 1080
rect 491260 1068 491266 1080
rect 497090 1068 497096 1080
rect 491260 1040 497096 1068
rect 491260 1028 491266 1040
rect 497090 1028 497096 1040
rect 497148 1028 497154 1080
rect 505186 1028 505192 1080
rect 505244 1068 505250 1080
rect 511258 1068 511264 1080
rect 505244 1040 511264 1068
rect 505244 1028 505250 1040
rect 511258 1028 511264 1040
rect 511316 1028 511322 1080
rect 512178 1028 512184 1080
rect 512236 1068 512242 1080
rect 517974 1068 517980 1080
rect 512236 1040 517980 1068
rect 512236 1028 512242 1040
rect 517974 1028 517980 1040
rect 518032 1028 518038 1080
rect 520182 1028 520188 1080
rect 520240 1068 520246 1080
rect 526622 1068 526628 1080
rect 520240 1040 526628 1068
rect 520240 1028 520246 1040
rect 526622 1028 526628 1040
rect 526680 1028 526686 1080
rect 529566 1028 529572 1080
rect 529624 1068 529630 1080
rect 536098 1068 536104 1080
rect 529624 1040 536104 1068
rect 529624 1028 529630 1040
rect 536098 1028 536104 1040
rect 536156 1028 536162 1080
rect 545850 1028 545856 1080
rect 545908 1068 545914 1080
rect 552658 1068 552664 1080
rect 545908 1040 552664 1068
rect 545908 1028 545914 1040
rect 552658 1028 552664 1040
rect 552716 1028 552722 1080
rect 559650 1028 559656 1080
rect 559708 1068 559714 1080
rect 566826 1068 566832 1080
rect 559708 1040 566832 1068
rect 559708 1028 559714 1040
rect 566826 1028 566832 1040
rect 566884 1028 566890 1080
rect 325418 960 325424 1012
rect 325476 1000 325482 1012
rect 327994 1000 328000 1012
rect 325476 972 328000 1000
rect 325476 960 325482 972
rect 327994 960 328000 972
rect 328052 960 328058 1012
rect 374178 960 374184 1012
rect 374236 1000 374242 1012
rect 377674 1000 377680 1012
rect 374236 972 377680 1000
rect 374236 960 374242 972
rect 377674 960 377680 972
rect 377732 960 377738 1012
rect 379882 960 379888 1012
rect 379940 1000 379946 1012
rect 383562 1000 383568 1012
rect 379940 972 383568 1000
rect 379940 960 379946 972
rect 383562 960 383568 972
rect 383620 960 383626 1012
rect 414750 960 414756 1012
rect 414808 1000 414814 1012
rect 418982 1000 418988 1012
rect 414808 972 418988 1000
rect 414808 960 414814 972
rect 418982 960 418988 972
rect 419040 960 419046 1012
rect 424042 960 424048 1012
rect 424100 1000 424106 1012
rect 428458 1000 428464 1012
rect 424100 972 428464 1000
rect 424100 960 424106 972
rect 428458 960 428464 972
rect 428516 960 428522 1012
rect 432138 960 432144 1012
rect 432196 1000 432202 1012
rect 436738 1000 436744 1012
rect 432196 972 436744 1000
rect 432196 960 432202 972
rect 436738 960 436744 972
rect 436796 960 436802 1012
rect 464614 960 464620 1012
rect 464672 1000 464678 1012
rect 469858 1000 469864 1012
rect 464672 972 469864 1000
rect 464672 960 464678 972
rect 469858 960 469864 972
rect 469916 960 469922 1012
rect 473906 960 473912 1012
rect 473964 1000 473970 1012
rect 479334 1000 479340 1012
rect 473964 972 479340 1000
rect 473964 960 473970 972
rect 479334 960 479340 972
rect 479392 960 479398 1012
rect 495986 960 495992 1012
rect 496044 1000 496050 1012
rect 501782 1000 501788 1012
rect 496044 972 501788 1000
rect 496044 960 496050 972
rect 501782 960 501788 972
rect 501840 960 501846 1012
rect 502886 960 502892 1012
rect 502944 1000 502950 1012
rect 508866 1000 508872 1012
rect 502944 972 508872 1000
rect 502944 960 502950 972
rect 508866 960 508872 972
rect 508924 960 508930 1012
rect 540054 960 540060 1012
rect 540112 1000 540118 1012
rect 546678 1000 546684 1012
rect 540112 972 546684 1000
rect 540112 960 540118 972
rect 546678 960 546684 972
rect 546736 960 546742 1012
rect 8754 892 8760 944
rect 8812 932 8818 944
rect 12158 932 12164 944
rect 8812 904 12164 932
rect 8812 892 8818 904
rect 12158 892 12164 904
rect 12216 892 12222 944
rect 121086 892 121092 944
rect 121144 932 121150 944
rect 122374 932 122380 944
rect 121144 904 122380 932
rect 121144 892 121150 904
rect 122374 892 122380 904
rect 122432 892 122438 944
rect 434346 892 434352 944
rect 434404 932 434410 944
rect 439130 932 439136 944
rect 434404 904 439136 932
rect 434404 892 434410 904
rect 439130 892 439136 904
rect 439188 892 439194 944
rect 463418 892 463424 944
rect 463476 932 463482 944
rect 468662 932 468668 944
rect 463476 904 468668 932
rect 463476 892 463482 904
rect 468662 892 468668 904
rect 468720 892 468726 944
rect 484302 892 484308 944
rect 484360 932 484366 944
rect 489914 932 489920 944
rect 484360 904 489920 932
rect 484360 892 484366 904
rect 489914 892 489920 904
rect 489972 892 489978 944
rect 347498 824 347504 876
rect 347556 864 347562 876
rect 350442 864 350448 876
rect 347556 836 350448 864
rect 347556 824 347562 836
rect 350442 824 350448 836
rect 350500 824 350506 876
rect 361390 824 361396 876
rect 361448 864 361454 876
rect 364610 864 364616 876
rect 361448 836 364616 864
rect 361448 824 361454 836
rect 364610 824 364616 836
rect 364668 824 364674 876
rect 368382 824 368388 876
rect 368440 864 368446 876
rect 371694 864 371700 876
rect 368440 836 371700 864
rect 368440 824 368446 836
rect 371694 824 371700 836
rect 371752 824 371758 876
rect 371786 824 371792 876
rect 371844 864 371850 876
rect 375282 864 375288 876
rect 371844 836 375288 864
rect 371844 824 371850 836
rect 375282 824 375288 836
rect 375340 824 375346 876
rect 384574 824 384580 876
rect 384632 864 384638 876
rect 388254 864 388260 876
rect 384632 836 388260 864
rect 384632 824 384638 836
rect 388254 824 388260 836
rect 388312 824 388318 876
rect 391566 824 391572 876
rect 391624 864 391630 876
rect 395338 864 395344 876
rect 391624 836 395344 864
rect 391624 824 391630 836
rect 395338 824 395344 836
rect 395396 824 395402 876
rect 397362 824 397368 876
rect 397420 864 397426 876
rect 401318 864 401324 876
rect 397420 836 401324 864
rect 397420 824 397426 836
rect 401318 824 401324 836
rect 401376 824 401382 876
rect 406654 824 406660 876
rect 406712 864 406718 876
rect 410794 864 410800 876
rect 406712 836 410800 864
rect 406712 824 406718 836
rect 410794 824 410800 836
rect 410852 824 410858 876
rect 419350 824 419356 876
rect 419408 864 419414 876
rect 423398 864 423404 876
rect 419408 836 423404 864
rect 419408 824 419414 836
rect 423398 824 423404 836
rect 423456 824 423462 876
rect 429838 824 429844 876
rect 429896 864 429902 876
rect 434438 864 434444 876
rect 429896 836 434444 864
rect 429896 824 429902 836
rect 434438 824 434444 836
rect 434496 824 434502 876
rect 443730 824 443736 876
rect 443788 864 443794 876
rect 448238 864 448244 876
rect 443788 836 448244 864
rect 443788 824 443794 836
rect 448238 824 448244 836
rect 448296 824 448302 876
rect 451826 824 451832 876
rect 451884 864 451890 876
rect 456518 864 456524 876
rect 451884 836 456524 864
rect 451884 824 451890 836
rect 456518 824 456524 836
rect 456576 824 456582 876
rect 476206 824 476212 876
rect 476264 864 476270 876
rect 481358 864 481364 876
rect 476264 836 481364 864
rect 476264 824 476270 836
rect 481358 824 481364 836
rect 481416 824 481422 876
rect 514478 824 514484 876
rect 514536 864 514542 876
rect 520734 864 520740 876
rect 514536 836 520740 864
rect 514536 824 514542 836
rect 520734 824 520740 836
rect 520792 824 520798 876
rect 521470 824 521476 876
rect 521528 864 521534 876
rect 527818 864 527824 876
rect 521528 836 527824 864
rect 521528 824 521534 836
rect 527818 824 527824 836
rect 527876 824 527882 876
rect 52546 688 52552 740
rect 52604 728 52610 740
rect 55030 728 55036 740
rect 52604 700 55036 728
rect 52604 688 52610 700
rect 55030 688 55036 700
rect 55088 688 55094 740
rect 59630 688 59636 740
rect 59688 728 59694 740
rect 61930 728 61936 740
rect 59688 700 61936 728
rect 59688 688 59694 700
rect 61930 688 61936 700
rect 61988 688 61994 740
rect 105722 688 105728 740
rect 105780 728 105786 740
rect 107286 728 107292 740
rect 105780 700 107292 728
rect 105780 688 105786 700
rect 107286 688 107292 700
rect 107344 688 107350 740
rect 274358 688 274364 740
rect 274416 728 274422 740
rect 276014 728 276020 740
rect 274416 700 276020 728
rect 274416 688 274422 700
rect 276014 688 276020 700
rect 276072 688 276078 740
rect 333514 688 333520 740
rect 333572 728 333578 740
rect 336274 728 336280 740
rect 333572 700 336280 728
rect 333572 688 333578 700
rect 336274 688 336280 700
rect 336332 688 336338 740
rect 338206 688 338212 740
rect 338264 728 338270 740
rect 340966 728 340972 740
rect 338264 700 340972 728
rect 338264 688 338270 700
rect 340966 688 340972 700
rect 341024 688 341030 740
rect 342806 688 342812 740
rect 342864 728 342870 740
rect 345750 728 345756 740
rect 342864 700 345756 728
rect 342864 688 342870 700
rect 345750 688 345756 700
rect 345808 688 345814 740
rect 346302 688 346308 740
rect 346360 728 346366 740
rect 349246 728 349252 740
rect 346360 700 349252 728
rect 346360 688 346366 700
rect 349246 688 349252 700
rect 349304 688 349310 740
rect 350902 688 350908 740
rect 350960 728 350966 740
rect 354030 728 354036 740
rect 350960 700 354036 728
rect 350960 688 350966 700
rect 354030 688 354036 700
rect 354088 688 354094 740
rect 365990 688 365996 740
rect 366048 728 366054 740
rect 369394 728 369400 740
rect 366048 700 369400 728
rect 366048 688 366054 700
rect 369394 688 369400 700
rect 369452 688 369458 740
rect 369486 688 369492 740
rect 369544 728 369550 740
rect 372890 728 372896 740
rect 369544 700 372896 728
rect 369544 688 369550 700
rect 372890 688 372896 700
rect 372948 688 372954 740
rect 544654 688 544660 740
rect 544712 728 544718 740
rect 551462 728 551468 740
rect 544712 700 551468 728
rect 544712 688 544718 700
rect 551462 688 551468 700
rect 551520 688 551526 740
rect 555142 688 555148 740
rect 555200 728 555206 740
rect 562042 728 562048 740
rect 555200 700 562048 728
rect 555200 688 555206 700
rect 562042 688 562048 700
rect 562100 688 562106 740
rect 494790 620 494796 672
rect 494848 660 494854 672
rect 500586 660 500592 672
rect 494848 632 500592 660
rect 494848 620 494854 632
rect 500586 620 500592 632
rect 500644 620 500650 672
rect 556246 620 556252 672
rect 556304 660 556310 672
rect 563146 660 563152 672
rect 556304 632 563152 660
rect 556304 620 556310 632
rect 563146 620 563152 632
rect 563204 620 563210 672
rect 69106 552 69112 604
rect 69164 592 69170 604
rect 71314 592 71320 604
rect 69164 564 71320 592
rect 69164 552 69170 564
rect 71314 552 71320 564
rect 71372 552 71378 604
rect 290642 552 290648 604
rect 290700 592 290706 604
rect 292574 592 292580 604
rect 290700 564 292580 592
rect 290700 552 290706 564
rect 292574 552 292580 564
rect 292632 552 292638 604
rect 304534 552 304540 604
rect 304592 592 304598 604
rect 306742 592 306748 604
rect 304592 564 306748 592
rect 304592 552 304598 564
rect 306742 552 306748 564
rect 306800 552 306806 604
rect 324222 552 324228 604
rect 324280 592 324286 604
rect 326798 592 326804 604
rect 324280 564 326804 592
rect 324280 552 324286 564
rect 326798 552 326804 564
rect 326856 552 326862 604
rect 327718 552 327724 604
rect 327776 592 327782 604
rect 330386 592 330392 604
rect 327776 564 330392 592
rect 327776 552 327782 564
rect 330386 552 330392 564
rect 330444 552 330450 604
rect 531866 552 531872 604
rect 531924 592 531930 604
rect 538398 592 538404 604
rect 531924 564 538404 592
rect 531924 552 531930 564
rect 538398 552 538404 564
rect 538456 552 538462 604
rect 544378 552 544384 604
rect 544436 552 544442 604
rect 549346 552 549352 604
rect 549404 592 549410 604
rect 556154 592 556160 604
rect 549404 564 556160 592
rect 549404 552 549410 564
rect 556154 552 556160 564
rect 556212 552 556218 604
rect 563330 552 563336 604
rect 563388 592 563394 604
rect 570322 592 570328 604
rect 563388 564 570328 592
rect 563388 552 563394 564
rect 570322 552 570328 564
rect 570380 552 570386 604
rect 537662 484 537668 536
rect 537720 524 537726 536
rect 544396 524 544424 552
rect 537720 496 544424 524
rect 537720 484 537726 496
rect 557534 484 557540 536
rect 557592 524 557598 536
rect 564618 524 564624 536
rect 557592 496 564624 524
rect 557592 484 557598 496
rect 564618 484 564624 496
rect 564676 484 564682 536
rect 535362 416 535368 468
rect 535420 456 535426 468
rect 542170 456 542176 468
rect 535420 428 542176 456
rect 535420 416 535426 428
rect 542170 416 542176 428
rect 542228 416 542234 468
rect 566642 416 566648 468
rect 566700 456 566706 468
rect 573726 456 573732 468
rect 566700 428 573732 456
rect 566700 416 566706 428
rect 573726 416 573732 428
rect 573784 416 573790 468
rect 383378 280 383384 332
rect 383436 320 383442 332
rect 386782 320 386788 332
rect 383436 292 386788 320
rect 383436 280 383442 292
rect 386782 280 386788 292
rect 386840 280 386846 332
rect 565446 280 565452 332
rect 565504 320 565510 332
rect 572898 320 572904 332
rect 565504 292 572904 320
rect 565504 280 565510 292
rect 572898 280 572904 292
rect 572956 280 572962 332
rect 576118 280 576124 332
rect 576176 320 576182 332
rect 583570 320 583576 332
rect 576176 292 583576 320
rect 576176 280 576182 292
rect 583570 280 583576 292
rect 583628 280 583634 332
rect 469306 212 469312 264
rect 469364 252 469370 264
rect 474182 252 474188 264
rect 469364 224 474188 252
rect 469364 212 469370 224
rect 474182 212 474188 224
rect 474240 212 474246 264
rect 508682 212 508688 264
rect 508740 252 508746 264
rect 514938 252 514944 264
rect 508740 224 514944 252
rect 508740 212 508746 224
rect 514938 212 514944 224
rect 514996 212 515002 264
rect 516778 212 516784 264
rect 516836 252 516842 264
rect 523218 252 523224 264
rect 516836 224 523224 252
rect 516836 212 516842 224
rect 523218 212 523224 224
rect 523276 212 523282 264
rect 553946 212 553952 264
rect 554004 252 554010 264
rect 560478 252 560484 264
rect 554004 224 560484 252
rect 554004 212 554010 224
rect 560478 212 560484 224
rect 560536 212 560542 264
rect 564250 212 564256 264
rect 564308 252 564314 264
rect 571334 252 571340 264
rect 564308 224 571340 252
rect 564308 212 564314 224
rect 571334 212 571340 224
rect 571392 212 571398 264
rect 574830 212 574836 264
rect 574888 252 574894 264
rect 581822 252 581828 264
rect 574888 224 581828 252
rect 574888 212 574894 224
rect 581822 212 581828 224
rect 581880 212 581886 264
rect 412450 144 412456 196
rect 412508 184 412514 196
rect 416866 184 416872 196
rect 412508 156 416872 184
rect 412508 144 412514 156
rect 416866 144 416872 156
rect 416924 144 416930 196
rect 470410 144 470416 196
rect 470468 184 470474 196
rect 475930 184 475936 196
rect 470468 156 475936 184
rect 470468 144 470474 156
rect 475930 144 475936 156
rect 475988 144 475994 196
rect 507486 144 507492 196
rect 507544 184 507550 196
rect 513374 184 513380 196
rect 507544 156 513380 184
rect 507544 144 507550 156
rect 513374 144 513380 156
rect 513432 144 513438 196
rect 392670 76 392676 128
rect 392728 116 392734 128
rect 396166 116 396172 128
rect 392728 88 396172 116
rect 392728 76 392734 88
rect 396166 76 396172 88
rect 396224 76 396230 128
rect 401962 76 401968 128
rect 402020 116 402026 128
rect 406194 116 406200 128
rect 402020 88 406200 116
rect 402020 76 402026 88
rect 406194 76 406200 88
rect 406252 76 406258 128
rect 421742 76 421748 128
rect 421800 116 421806 128
rect 425790 116 425796 128
rect 421800 88 425796 116
rect 421800 76 421806 88
rect 425790 76 425796 88
rect 425848 76 425854 128
rect 431034 76 431040 128
rect 431092 116 431098 128
rect 435174 116 435180 128
rect 431092 88 435180 116
rect 431092 76 431098 88
rect 435174 76 435180 88
rect 435232 76 435238 128
rect 460014 76 460020 128
rect 460072 116 460078 128
rect 464982 116 464988 128
rect 460072 88 464988 116
rect 460072 76 460078 88
rect 464982 76 464988 88
rect 465040 76 465046 128
rect 515674 76 515680 128
rect 515732 116 515738 128
rect 521654 116 521660 128
rect 515732 88 521660 116
rect 515732 76 515738 88
rect 521654 76 521660 88
rect 521712 76 521718 128
rect 524966 76 524972 128
rect 525024 116 525030 128
rect 531498 116 531504 128
rect 525024 88 531504 116
rect 525024 76 525030 88
rect 531498 76 531504 88
rect 531556 76 531562 128
rect 573634 76 573640 128
rect 573692 116 573698 128
rect 581178 116 581184 128
rect 573692 88 581184 116
rect 573692 76 573698 88
rect 581178 76 581184 88
rect 581236 76 581242 128
rect 354398 8 354404 60
rect 354456 48 354462 60
rect 357342 48 357348 60
rect 354456 20 357348 48
rect 354456 8 354462 20
rect 357342 8 357348 20
rect 357400 8 357406 60
rect 499206 8 499212 60
rect 499264 48 499270 60
rect 505554 48 505560 60
rect 499264 20 505560 48
rect 499264 8 499270 20
rect 505554 8 505560 20
rect 505612 8 505618 60
rect 506290 8 506296 60
rect 506348 48 506354 60
rect 512086 48 512092 60
rect 506348 20 512092 48
rect 506348 8 506354 20
rect 512086 8 512092 20
rect 512144 8 512150 60
rect 528462 8 528468 60
rect 528520 48 528526 60
rect 534534 48 534540 60
rect 528520 20 534540 48
rect 528520 8 528526 20
rect 534534 8 534540 20
rect 534592 8 534598 60
rect 536558 8 536564 60
rect 536616 48 536622 60
rect 542814 48 542820 60
rect 536616 20 542820 48
rect 536616 8 536622 20
rect 542814 8 542820 20
rect 542872 8 542878 60
rect 546954 8 546960 60
rect 547012 48 547018 60
rect 553946 48 553952 60
rect 547012 20 553952 48
rect 547012 8 547018 20
rect 553946 8 553952 20
rect 554004 8 554010 60
rect 572530 8 572536 60
rect 572588 48 572594 60
rect 579614 48 579620 60
rect 572588 20 579620 48
rect 572588 8 572594 20
rect 579614 8 579620 20
rect 579672 8 579678 60
<< via1 >>
rect 3884 700748 3936 700800
rect 8116 700748 8168 700800
rect 102048 700748 102100 700800
rect 105452 700748 105504 700800
rect 200028 700748 200080 700800
rect 202788 700748 202840 700800
rect 314476 700748 314528 700800
rect 316316 700748 316368 700800
rect 363512 700408 363564 700460
rect 364984 700408 365036 700460
rect 412456 700408 412508 700460
rect 413652 700408 413704 700460
rect 20352 700204 20404 700256
rect 24308 700204 24360 700256
rect 36728 700204 36780 700256
rect 40500 700204 40552 700256
rect 69388 700204 69440 700256
rect 72976 700204 73028 700256
rect 85764 700204 85816 700256
rect 89168 700204 89220 700256
rect 134708 700204 134760 700256
rect 137836 700204 137888 700256
rect 167368 700204 167420 700256
rect 170312 700204 170364 700256
rect 183744 700204 183796 700256
rect 186504 700204 186556 700256
rect 232780 700204 232832 700256
rect 235172 700204 235224 700256
rect 249064 700204 249116 700256
rect 251456 700204 251508 700256
rect 265440 700204 265492 700256
rect 267648 700204 267700 700256
rect 281816 700204 281868 700256
rect 283840 700204 283892 700256
rect 330760 700204 330812 700256
rect 332508 700204 332560 700256
rect 347136 700204 347188 700256
rect 348792 700204 348844 700256
rect 396172 700204 396224 700256
rect 397460 700204 397512 700256
rect 428832 700204 428884 700256
rect 429844 700204 429896 700256
rect 445208 700204 445260 700256
rect 446128 700204 446180 700256
rect 461492 700204 461544 700256
rect 462320 700204 462372 700256
rect 118424 700136 118476 700188
rect 121644 700136 121696 700188
rect 151084 700136 151136 700188
rect 154120 700136 154172 700188
rect 216404 700136 216456 700188
rect 218980 700136 219032 700188
rect 298008 700136 298060 700188
rect 300124 700136 300176 700188
rect 477868 700136 477920 700188
rect 478512 700136 478564 700188
rect 494244 700136 494296 700188
rect 494796 700136 494848 700188
rect 53012 700000 53064 700052
rect 56784 700000 56836 700052
rect 379796 699864 379848 699916
rect 381176 699864 381228 699916
rect 578332 644512 578384 644564
rect 580908 644512 580960 644564
rect 578884 257796 578936 257848
rect 580908 257796 580960 257848
rect 578516 151444 578568 151496
rect 580908 151444 580960 151496
rect 578332 44956 578384 45008
rect 579988 44956 580040 45008
rect 11152 3884 11204 3936
rect 14508 3884 14560 3936
rect 14740 3884 14792 3936
rect 18004 3884 18056 3936
rect 20628 3884 20680 3936
rect 23800 3884 23852 3936
rect 24216 3884 24268 3936
rect 27296 3884 27348 3936
rect 27712 3884 27764 3936
rect 30700 3884 30752 3936
rect 32404 3884 32456 3936
rect 35392 3884 35444 3936
rect 38384 3884 38436 3936
rect 41188 3884 41240 3936
rect 43076 3884 43128 3936
rect 45788 3884 45840 3936
rect 46664 3884 46716 3936
rect 49284 3884 49336 3936
rect 50160 3884 50212 3936
rect 52780 3884 52832 3936
rect 56048 3884 56100 3936
rect 58576 3884 58628 3936
rect 72608 3884 72660 3936
rect 74860 3884 74912 3936
rect 247636 3884 247688 3936
rect 248604 3884 248656 3936
rect 285908 3884 285960 3936
rect 287796 3884 287848 3936
rect 1676 3816 1728 3868
rect 5216 3816 5268 3868
rect 13544 3816 13596 3868
rect 16808 3816 16860 3868
rect 19432 3816 19484 3868
rect 22604 3816 22656 3868
rect 23020 3816 23072 3868
rect 26100 3816 26152 3868
rect 26516 3816 26568 3868
rect 29596 3816 29648 3868
rect 30104 3816 30156 3868
rect 33092 3816 33144 3868
rect 33600 3816 33652 3868
rect 36588 3816 36640 3868
rect 37188 3816 37240 3868
rect 39992 3816 40044 3868
rect 41880 3816 41932 3868
rect 44684 3816 44736 3868
rect 45468 3816 45520 3868
rect 48180 3816 48232 3868
rect 48964 3816 49016 3868
rect 51584 3816 51636 3868
rect 53748 3816 53800 3868
rect 56276 3816 56328 3868
rect 57244 3816 57296 3868
rect 59772 3816 59824 3868
rect 71504 3816 71556 3868
rect 73664 3816 73716 3868
rect 78588 3816 78640 3868
rect 80656 3816 80708 3868
rect 80888 3816 80940 3868
rect 82956 3816 83008 3868
rect 87972 3816 88024 3868
rect 89948 3816 90000 3868
rect 96252 3816 96304 3868
rect 98044 3816 98096 3868
rect 244140 3816 244192 3868
rect 245200 3816 245252 3868
rect 256928 3816 256980 3868
rect 258264 3816 258316 3868
rect 259228 3816 259280 3868
rect 260656 3816 260708 3868
rect 261620 3816 261672 3868
rect 262956 3816 263008 3868
rect 263920 3816 263972 3868
rect 265348 3816 265400 3868
rect 268520 3816 268572 3868
rect 270040 3816 270092 3868
rect 270820 3816 270872 3868
rect 272432 3816 272484 3868
rect 275512 3816 275564 3868
rect 277124 3816 277176 3868
rect 277812 3816 277864 3868
rect 279516 3816 279568 3868
rect 284804 3816 284856 3868
rect 286600 3816 286652 3868
rect 292900 3816 292952 3868
rect 294880 3816 294932 3868
rect 299892 3816 299944 3868
rect 301964 3816 302016 3868
rect 306792 3816 306844 3868
rect 309048 3816 309100 3868
rect 572 3748 624 3800
rect 4112 3748 4164 3800
rect 7656 3748 7708 3800
rect 11012 3748 11064 3800
rect 12348 3748 12400 3800
rect 15704 3748 15756 3800
rect 15936 3748 15988 3800
rect 19108 3748 19160 3800
rect 21824 3748 21876 3800
rect 24904 3748 24956 3800
rect 25320 3748 25372 3800
rect 28400 3748 28452 3800
rect 31300 3748 31352 3800
rect 34196 3748 34248 3800
rect 34796 3748 34848 3800
rect 37692 3748 37744 3800
rect 40684 3748 40736 3800
rect 43488 3748 43540 3800
rect 44272 3748 44324 3800
rect 46984 3748 47036 3800
rect 47860 3748 47912 3800
rect 50480 3748 50532 3800
rect 51356 3748 51408 3800
rect 53976 3748 54028 3800
rect 54944 3748 54996 3800
rect 57380 3748 57432 3800
rect 58440 3748 58492 3800
rect 60876 3748 60928 3800
rect 64328 3748 64380 3800
rect 66672 3748 66724 3800
rect 67088 3748 67140 3800
rect 69064 3748 69116 3800
rect 70308 3748 70360 3800
rect 72468 3748 72520 3800
rect 73804 3748 73856 3800
rect 75964 3748 76016 3800
rect 79692 3748 79744 3800
rect 81760 3748 81812 3800
rect 86868 3748 86920 3800
rect 88752 3748 88804 3800
rect 95148 3748 95200 3800
rect 96848 3748 96900 3800
rect 103336 3748 103388 3800
rect 104944 3748 104996 3800
rect 216356 3748 216408 3800
rect 216864 3748 216916 3800
rect 222152 3748 222204 3800
rect 222752 3748 222804 3800
rect 224452 3748 224504 3800
rect 225144 3748 225196 3800
rect 230248 3748 230300 3800
rect 231032 3748 231084 3800
rect 231444 3748 231496 3800
rect 232228 3748 232280 3800
rect 232548 3748 232600 3800
rect 233424 3748 233476 3800
rect 233744 3748 233796 3800
rect 234620 3748 234672 3800
rect 237240 3748 237292 3800
rect 238116 3748 238168 3800
rect 238344 3748 238396 3800
rect 239312 3748 239364 3800
rect 239540 3748 239592 3800
rect 240508 3748 240560 3800
rect 240736 3748 240788 3800
rect 241704 3748 241756 3800
rect 241840 3748 241892 3800
rect 242900 3748 242952 3800
rect 245336 3748 245388 3800
rect 246396 3748 246448 3800
rect 246532 3748 246584 3800
rect 247592 3748 247644 3800
rect 250028 3748 250080 3800
rect 251180 3748 251232 3800
rect 252328 3748 252380 3800
rect 253480 3748 253532 3800
rect 255824 3748 255876 3800
rect 257068 3748 257120 3800
rect 258124 3748 258176 3800
rect 259460 3748 259512 3800
rect 260424 3748 260476 3800
rect 261760 3748 261812 3800
rect 262724 3748 262776 3800
rect 264152 3748 264204 3800
rect 265024 3748 265076 3800
rect 266544 3748 266596 3800
rect 267416 3748 267468 3800
rect 268844 3748 268896 3800
rect 269716 3748 269768 3800
rect 271236 3748 271288 3800
rect 272016 3748 272068 3800
rect 273628 3748 273680 3800
rect 276708 3748 276760 3800
rect 278320 3748 278372 3800
rect 279008 3748 279060 3800
rect 280712 3748 280764 3800
rect 283608 3748 283660 3800
rect 285404 3748 285456 3800
rect 287104 3748 287156 3800
rect 288992 3748 289044 3800
rect 291704 3748 291756 3800
rect 293684 3748 293736 3800
rect 294096 3748 294148 3800
rect 296076 3748 296128 3800
rect 298696 3748 298748 3800
rect 300768 3748 300820 3800
rect 300996 3748 301048 3800
rect 303160 3748 303212 3800
rect 307988 3748 308040 3800
rect 310244 3748 310296 3800
rect 316084 3748 316136 3800
rect 318524 3748 318576 3800
rect 323076 3748 323128 3800
rect 325608 3748 325660 3800
rect 63224 3000 63276 3052
rect 65524 3000 65576 3052
rect 4068 2864 4120 2916
rect 7472 2864 7524 2916
rect 18236 2864 18288 2916
rect 21456 2864 21508 2916
rect 253388 2864 253440 2916
rect 254676 2864 254728 2916
rect 6460 2796 6512 2848
rect 9864 2796 9916 2848
rect 9956 2796 10008 2848
rect 13268 2796 13320 2848
rect 17040 2796 17092 2848
rect 20260 2796 20312 2848
rect 28908 2796 28960 2848
rect 31852 2796 31904 2848
rect 35992 2796 36044 2848
rect 38844 2796 38896 2848
rect 39580 2796 39632 2848
rect 42340 2796 42392 2848
rect 62028 2796 62080 2848
rect 64420 2796 64472 2848
rect 65524 2796 65576 2848
rect 67824 2796 67876 2848
rect 248880 2796 248932 2848
rect 249984 2796 250036 2848
rect 251088 2796 251140 2848
rect 252376 2796 252428 2848
rect 254584 2796 254636 2848
rect 255872 2796 255924 2848
rect 309232 2796 309284 2848
rect 311440 2796 311492 2848
rect 315028 2796 315080 2848
rect 317328 2796 317380 2848
rect 411168 2796 411220 2848
rect 415492 2796 415544 2848
rect 440148 2796 440200 2848
rect 445024 2796 445076 2848
rect 449532 2796 449584 2848
rect 454500 2796 454552 2848
rect 478512 2796 478564 2848
rect 484032 2796 484084 2848
rect 487804 2796 487856 2848
rect 493508 2796 493560 2848
rect 3240 1300 3292 1352
rect 6368 1300 6420 1352
rect 60832 1300 60884 1352
rect 63316 1300 63368 1352
rect 67916 1300 67968 1352
rect 70124 1300 70176 1352
rect 76196 1300 76248 1352
rect 78220 1300 78272 1352
rect 83280 1300 83332 1352
rect 85212 1300 85264 1352
rect 85672 1300 85724 1352
rect 87512 1300 87564 1352
rect 89168 1300 89220 1352
rect 91008 1300 91060 1352
rect 91560 1300 91612 1352
rect 93308 1300 93360 1352
rect 93952 1300 94004 1352
rect 95700 1300 95752 1352
rect 97448 1300 97500 1352
rect 99104 1300 99156 1352
rect 101036 1300 101088 1352
rect 102600 1300 102652 1352
rect 104532 1300 104584 1352
rect 106096 1300 106148 1352
rect 106924 1300 106976 1352
rect 108396 1300 108448 1352
rect 109316 1300 109368 1352
rect 110696 1300 110748 1352
rect 112812 1300 112864 1352
rect 114192 1300 114244 1352
rect 116400 1300 116452 1352
rect 117688 1300 117740 1352
rect 119896 1300 119948 1352
rect 121184 1300 121236 1352
rect 125876 1300 125928 1352
rect 126980 1300 127032 1352
rect 129372 1300 129424 1352
rect 130476 1300 130528 1352
rect 130568 1300 130620 1352
rect 131580 1300 131632 1352
rect 131764 1300 131816 1352
rect 132776 1300 132828 1352
rect 132960 1300 133012 1352
rect 133972 1300 134024 1352
rect 137652 1300 137704 1352
rect 138572 1300 138624 1352
rect 144736 1300 144788 1352
rect 145564 1300 145616 1352
rect 145932 1300 145984 1352
rect 146668 1300 146720 1352
rect 148324 1300 148376 1352
rect 149060 1300 149112 1352
rect 154212 1300 154264 1352
rect 154856 1300 154908 1352
rect 162492 1300 162544 1352
rect 162952 1300 163004 1352
rect 266268 1300 266320 1352
rect 267740 1300 267792 1352
rect 273168 1300 273220 1352
rect 274824 1300 274876 1352
rect 280068 1300 280120 1352
rect 281908 1300 281960 1352
rect 282552 1300 282604 1352
rect 284300 1300 284352 1352
rect 288348 1300 288400 1352
rect 290188 1300 290240 1352
rect 295248 1300 295300 1352
rect 297272 1300 297324 1352
rect 297548 1300 297600 1352
rect 299664 1300 299716 1352
rect 302148 1300 302200 1352
rect 304356 1300 304408 1352
rect 305736 1300 305788 1352
rect 307944 1300 307996 1352
rect 310336 1300 310388 1352
rect 312636 1300 312688 1352
rect 313832 1300 313884 1352
rect 316224 1300 316276 1352
rect 317236 1300 317288 1352
rect 319720 1300 319772 1352
rect 321928 1300 321980 1352
rect 324412 1300 324464 1352
rect 326620 1300 326672 1352
rect 329196 1300 329248 1352
rect 332416 1300 332468 1352
rect 335084 1300 335136 1352
rect 335912 1300 335964 1352
rect 338672 1300 338724 1352
rect 339316 1300 339368 1352
rect 342168 1300 342220 1352
rect 345112 1300 345164 1352
rect 348056 1300 348108 1352
rect 349804 1300 349856 1352
rect 352840 1300 352892 1352
rect 353208 1300 353260 1352
rect 356336 1300 356388 1352
rect 356704 1300 356756 1352
rect 359924 1300 359976 1352
rect 362592 1300 362644 1352
rect 365812 1300 365864 1352
rect 367192 1300 367244 1352
rect 370596 1300 370648 1352
rect 370688 1300 370740 1352
rect 374092 1300 374144 1352
rect 376392 1300 376444 1352
rect 379980 1300 380032 1352
rect 385776 1300 385828 1352
rect 389456 1300 389508 1352
rect 395068 1300 395120 1352
rect 398932 1300 398984 1352
rect 399668 1300 399720 1352
rect 403624 1300 403676 1352
rect 405464 1300 405516 1352
rect 409604 1300 409656 1352
rect 413560 1300 413612 1352
rect 417884 1300 417936 1352
rect 422852 1300 422904 1352
rect 427268 1300 427320 1352
rect 427544 1300 427596 1352
rect 431868 1300 431920 1352
rect 433248 1300 433300 1352
rect 437848 1300 437900 1352
rect 441436 1300 441488 1352
rect 445852 1300 445904 1352
rect 447232 1300 447284 1352
rect 452108 1300 452160 1352
rect 453028 1300 453080 1352
rect 458088 1300 458140 1352
rect 458824 1300 458876 1352
rect 463976 1300 464028 1352
rect 471612 1300 471664 1352
rect 476580 1300 476632 1352
rect 477408 1300 477460 1352
rect 482468 1300 482520 1352
rect 483204 1300 483256 1352
rect 488816 1300 488868 1352
rect 490104 1300 490156 1352
rect 495532 1300 495584 1352
rect 497096 1300 497148 1352
rect 502984 1300 503036 1352
rect 504088 1300 504140 1352
rect 509700 1300 509752 1352
rect 509884 1300 509936 1352
rect 515772 1300 515824 1352
rect 519176 1300 519228 1352
rect 525432 1300 525484 1352
rect 526076 1300 526128 1352
rect 532148 1300 532200 1352
rect 534264 1300 534316 1352
rect 540428 1300 540480 1352
rect 542268 1300 542320 1352
rect 549076 1300 549128 1352
rect 551652 1300 551704 1352
rect 558552 1300 558604 1352
rect 560944 1300 560996 1352
rect 568028 1300 568080 1352
rect 571248 1300 571300 1352
rect 578608 1300 578660 1352
rect 75000 1232 75052 1284
rect 77116 1232 77168 1284
rect 77392 1232 77444 1284
rect 79416 1232 79468 1284
rect 82084 1232 82136 1284
rect 84016 1232 84068 1284
rect 84476 1232 84528 1284
rect 86408 1232 86460 1284
rect 90364 1232 90416 1284
rect 92204 1232 92256 1284
rect 92756 1232 92808 1284
rect 94504 1232 94556 1284
rect 98644 1232 98696 1284
rect 100300 1232 100352 1284
rect 102232 1232 102284 1284
rect 103796 1232 103848 1284
rect 108120 1232 108172 1284
rect 109592 1232 109644 1284
rect 110512 1232 110564 1284
rect 111892 1232 111944 1284
rect 115204 1232 115256 1284
rect 116584 1232 116636 1284
rect 117596 1232 117648 1284
rect 118884 1232 118936 1284
rect 122288 1232 122340 1284
rect 123484 1232 123536 1284
rect 124680 1232 124732 1284
rect 125784 1232 125836 1284
rect 128176 1232 128228 1284
rect 129280 1232 129332 1284
rect 136456 1232 136508 1284
rect 137376 1232 137428 1284
rect 138848 1232 138900 1284
rect 139768 1232 139820 1284
rect 140044 1232 140096 1284
rect 140872 1232 140924 1284
rect 281356 1232 281408 1284
rect 283104 1232 283156 1284
rect 289452 1232 289504 1284
rect 291384 1232 291436 1284
rect 296444 1232 296496 1284
rect 298468 1232 298520 1284
rect 303344 1232 303396 1284
rect 305552 1232 305604 1284
rect 312544 1232 312596 1284
rect 315028 1232 315080 1284
rect 318432 1232 318484 1284
rect 320916 1232 320968 1284
rect 328920 1232 328972 1284
rect 331588 1232 331640 1284
rect 334716 1232 334768 1284
rect 337476 1232 337528 1284
rect 340512 1232 340564 1284
rect 343364 1232 343416 1284
rect 344008 1232 344060 1284
rect 346952 1232 347004 1284
rect 348608 1232 348660 1284
rect 351644 1232 351696 1284
rect 352104 1232 352156 1284
rect 355232 1232 355284 1284
rect 355600 1232 355652 1284
rect 358728 1232 358780 1284
rect 359096 1232 359148 1284
rect 362316 1232 362368 1284
rect 363696 1232 363748 1284
rect 367008 1232 367060 1284
rect 372988 1232 373040 1284
rect 376484 1232 376536 1284
rect 377588 1232 377640 1284
rect 381176 1232 381228 1284
rect 388076 1232 388128 1284
rect 391848 1232 391900 1284
rect 393872 1232 393924 1284
rect 397736 1232 397788 1284
rect 403164 1232 403216 1284
rect 407212 1232 407264 1284
rect 410064 1232 410116 1284
rect 414296 1232 414348 1284
rect 418252 1232 418304 1284
rect 422576 1232 422628 1284
rect 426348 1232 426400 1284
rect 430856 1232 430908 1284
rect 435640 1232 435692 1284
rect 439964 1232 440016 1284
rect 442632 1232 442684 1284
rect 447416 1232 447468 1284
rect 457628 1232 457680 1284
rect 462412 1232 462464 1284
rect 468116 1232 468168 1284
rect 473084 1232 473136 1284
rect 475108 1232 475160 1284
rect 480536 1232 480588 1284
rect 485504 1232 485556 1284
rect 490748 1232 490800 1284
rect 492496 1232 492548 1284
rect 498200 1232 498252 1284
rect 498292 1232 498344 1284
rect 503812 1232 503864 1284
rect 510988 1232 511040 1284
rect 517152 1232 517204 1284
rect 517980 1232 518032 1284
rect 523868 1232 523920 1284
rect 527272 1232 527324 1284
rect 533712 1232 533764 1284
rect 541164 1232 541216 1284
rect 547880 1232 547932 1284
rect 548156 1232 548208 1284
rect 554964 1232 555016 1284
rect 562048 1232 562100 1284
rect 569132 1232 569184 1284
rect 570144 1232 570196 1284
rect 577412 1232 577464 1284
rect 99840 1164 99892 1216
rect 101496 1164 101548 1216
rect 114008 1164 114060 1216
rect 115388 1164 115440 1216
rect 311532 1164 311584 1216
rect 313832 1164 313884 1216
rect 319628 1164 319680 1216
rect 322112 1164 322164 1216
rect 330024 1164 330076 1216
rect 332692 1164 332744 1216
rect 337016 1164 337068 1216
rect 339868 1164 339920 1216
rect 341708 1164 341760 1216
rect 344560 1164 344612 1216
rect 357900 1164 357952 1216
rect 361120 1164 361172 1216
rect 364892 1164 364944 1216
rect 368204 1164 368256 1216
rect 375288 1164 375340 1216
rect 378876 1164 378928 1216
rect 381084 1164 381136 1216
rect 384764 1164 384816 1216
rect 390376 1164 390428 1216
rect 394240 1164 394292 1216
rect 396172 1164 396224 1216
rect 400128 1164 400180 1216
rect 400864 1164 400916 1216
rect 404820 1164 404872 1216
rect 407764 1164 407816 1216
rect 411904 1164 411956 1216
rect 420552 1164 420604 1216
rect 424968 1164 425020 1216
rect 425152 1164 425204 1216
rect 429660 1164 429712 1216
rect 436744 1164 436796 1216
rect 441528 1164 441580 1216
rect 444932 1164 444984 1216
rect 449808 1164 449860 1216
rect 450728 1164 450780 1216
rect 455696 1164 455748 1216
rect 456524 1164 456576 1216
rect 461584 1164 461636 1216
rect 462228 1164 462280 1216
rect 467472 1164 467524 1216
rect 472716 1164 472768 1216
rect 478144 1164 478196 1216
rect 480904 1164 480956 1216
rect 486424 1164 486476 1216
rect 486700 1164 486752 1216
rect 492312 1164 492364 1216
rect 493600 1164 493652 1216
rect 499396 1164 499448 1216
rect 500592 1164 500644 1216
rect 506480 1164 506532 1216
rect 522672 1164 522724 1216
rect 529020 1164 529072 1216
rect 530768 1164 530820 1216
rect 537208 1164 537260 1216
rect 538864 1164 538916 1216
rect 545488 1164 545540 1216
rect 550456 1164 550508 1216
rect 557356 1164 557408 1216
rect 558460 1164 558512 1216
rect 565636 1164 565688 1216
rect 569040 1164 569092 1216
rect 576308 1164 576360 1216
rect 5632 1096 5684 1148
rect 8668 1096 8720 1148
rect 111616 1096 111668 1148
rect 113088 1096 113140 1148
rect 123484 1096 123536 1148
rect 124772 1096 124824 1148
rect 320824 1096 320876 1148
rect 323308 1096 323360 1148
rect 331128 1096 331180 1148
rect 333888 1096 333940 1148
rect 360108 1096 360160 1148
rect 363512 1096 363564 1148
rect 382188 1096 382240 1148
rect 385960 1096 386012 1148
rect 389272 1096 389324 1148
rect 393044 1096 393096 1148
rect 398472 1096 398524 1148
rect 402520 1096 402572 1148
rect 404268 1096 404320 1148
rect 408408 1096 408460 1148
rect 408960 1096 409012 1148
rect 413100 1096 413152 1148
rect 415952 1096 416004 1148
rect 420184 1096 420236 1148
rect 428648 1096 428700 1148
rect 433248 1096 433300 1148
rect 439136 1096 439188 1148
rect 443828 1096 443880 1148
rect 448428 1096 448480 1148
rect 453304 1096 453356 1148
rect 454224 1096 454276 1148
rect 459192 1096 459244 1148
rect 465816 1096 465868 1148
rect 470692 1096 470744 1148
rect 482008 1096 482060 1148
rect 487252 1096 487304 1148
rect 489000 1096 489052 1148
rect 494704 1096 494756 1148
rect 501788 1096 501840 1148
rect 507308 1096 507360 1148
rect 513288 1096 513340 1148
rect 519544 1096 519596 1148
rect 523776 1096 523828 1148
rect 530124 1096 530176 1148
rect 533068 1096 533120 1148
rect 539600 1096 539652 1148
rect 543464 1096 543516 1148
rect 550272 1096 550324 1148
rect 552756 1096 552808 1148
rect 559748 1096 559800 1148
rect 567844 1096 567896 1148
rect 575112 1096 575164 1148
rect 378784 1028 378836 1080
rect 382372 1028 382424 1080
rect 386880 1028 386932 1080
rect 390652 1028 390704 1080
rect 417056 1028 417108 1080
rect 421380 1028 421432 1080
rect 437940 1028 437992 1080
rect 442632 1028 442684 1080
rect 446036 1028 446088 1080
rect 450912 1028 450964 1080
rect 455328 1028 455380 1080
rect 460112 1028 460164 1080
rect 461124 1028 461176 1080
rect 466276 1028 466328 1080
rect 466920 1028 466972 1080
rect 472256 1028 472308 1080
rect 479708 1028 479760 1080
rect 484860 1028 484912 1080
rect 491208 1028 491260 1080
rect 497096 1028 497148 1080
rect 505192 1028 505244 1080
rect 511264 1028 511316 1080
rect 512184 1028 512236 1080
rect 517980 1028 518032 1080
rect 520188 1028 520240 1080
rect 526628 1028 526680 1080
rect 529572 1028 529624 1080
rect 536104 1028 536156 1080
rect 545856 1028 545908 1080
rect 552664 1028 552716 1080
rect 559656 1028 559708 1080
rect 566832 1028 566884 1080
rect 325424 960 325476 1012
rect 328000 960 328052 1012
rect 374184 960 374236 1012
rect 377680 960 377732 1012
rect 379888 960 379940 1012
rect 383568 960 383620 1012
rect 414756 960 414808 1012
rect 418988 960 419040 1012
rect 424048 960 424100 1012
rect 428464 960 428516 1012
rect 432144 960 432196 1012
rect 436744 960 436796 1012
rect 464620 960 464672 1012
rect 469864 960 469916 1012
rect 473912 960 473964 1012
rect 479340 960 479392 1012
rect 495992 960 496044 1012
rect 501788 960 501840 1012
rect 502892 960 502944 1012
rect 508872 960 508924 1012
rect 540060 960 540112 1012
rect 546684 960 546736 1012
rect 8760 892 8812 944
rect 12164 892 12216 944
rect 121092 892 121144 944
rect 122380 892 122432 944
rect 434352 892 434404 944
rect 439136 892 439188 944
rect 463424 892 463476 944
rect 468668 892 468720 944
rect 484308 892 484360 944
rect 489920 892 489972 944
rect 347504 824 347556 876
rect 350448 824 350500 876
rect 361396 824 361448 876
rect 364616 824 364668 876
rect 368388 824 368440 876
rect 371700 824 371752 876
rect 371792 824 371844 876
rect 375288 824 375340 876
rect 384580 824 384632 876
rect 388260 824 388312 876
rect 391572 824 391624 876
rect 395344 824 395396 876
rect 397368 824 397420 876
rect 401324 824 401376 876
rect 406660 824 406712 876
rect 410800 824 410852 876
rect 419356 824 419408 876
rect 423404 824 423456 876
rect 429844 824 429896 876
rect 434444 824 434496 876
rect 443736 824 443788 876
rect 448244 824 448296 876
rect 451832 824 451884 876
rect 456524 824 456576 876
rect 476212 824 476264 876
rect 481364 824 481416 876
rect 514484 824 514536 876
rect 520740 824 520792 876
rect 521476 824 521528 876
rect 527824 824 527876 876
rect 52552 688 52604 740
rect 55036 688 55088 740
rect 59636 688 59688 740
rect 61936 688 61988 740
rect 105728 688 105780 740
rect 107292 688 107344 740
rect 274364 688 274416 740
rect 276020 688 276072 740
rect 333520 688 333572 740
rect 336280 688 336332 740
rect 338212 688 338264 740
rect 340972 688 341024 740
rect 342812 688 342864 740
rect 345756 688 345808 740
rect 346308 688 346360 740
rect 349252 688 349304 740
rect 350908 688 350960 740
rect 354036 688 354088 740
rect 365996 688 366048 740
rect 369400 688 369452 740
rect 369492 688 369544 740
rect 372896 688 372948 740
rect 544660 688 544712 740
rect 551468 688 551520 740
rect 555148 688 555200 740
rect 562048 688 562100 740
rect 494796 620 494848 672
rect 500592 620 500644 672
rect 556252 620 556304 672
rect 563152 620 563204 672
rect 69112 552 69164 604
rect 71320 552 71372 604
rect 290648 552 290700 604
rect 292580 552 292632 604
rect 304540 552 304592 604
rect 306748 552 306800 604
rect 324228 552 324280 604
rect 326804 552 326856 604
rect 327724 552 327776 604
rect 330392 552 330444 604
rect 531872 552 531924 604
rect 538404 552 538456 604
rect 544384 552 544436 604
rect 549352 552 549404 604
rect 556160 552 556212 604
rect 563336 552 563388 604
rect 570328 552 570380 604
rect 537668 484 537720 536
rect 557540 484 557592 536
rect 564624 484 564676 536
rect 535368 416 535420 468
rect 542176 416 542228 468
rect 566648 416 566700 468
rect 573732 416 573784 468
rect 383384 280 383436 332
rect 386788 280 386840 332
rect 565452 280 565504 332
rect 572904 280 572956 332
rect 576124 280 576176 332
rect 583576 280 583628 332
rect 469312 212 469364 264
rect 474188 212 474240 264
rect 508688 212 508740 264
rect 514944 212 514996 264
rect 516784 212 516836 264
rect 523224 212 523276 264
rect 553952 212 554004 264
rect 560484 212 560536 264
rect 564256 212 564308 264
rect 571340 212 571392 264
rect 574836 212 574888 264
rect 581828 212 581880 264
rect 412456 144 412508 196
rect 416872 144 416924 196
rect 470416 144 470468 196
rect 475936 144 475988 196
rect 507492 144 507544 196
rect 513380 144 513432 196
rect 392676 76 392728 128
rect 396172 76 396224 128
rect 401968 76 402020 128
rect 406200 76 406252 128
rect 421748 76 421800 128
rect 425796 76 425848 128
rect 431040 76 431092 128
rect 435180 76 435232 128
rect 460020 76 460072 128
rect 464988 76 465040 128
rect 515680 76 515732 128
rect 521660 76 521712 128
rect 524972 76 525024 128
rect 531504 76 531556 128
rect 573640 76 573692 128
rect 581184 76 581236 128
rect 354404 8 354456 60
rect 357348 8 357400 60
rect 499212 8 499264 60
rect 505560 8 505612 60
rect 506296 8 506348 60
rect 512092 8 512144 60
rect 528468 8 528520 60
rect 534540 8 534592 60
rect 536564 8 536616 60
rect 542820 8 542872 60
rect 546960 8 547012 60
rect 553952 8 554004 60
rect 572536 8 572588 60
rect 579620 8 579672 60
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510632 703582 510844 703610
rect 8128 700806 8156 703520
rect 3884 700800 3936 700806
rect 3884 700742 3936 700748
rect 8116 700800 8168 700806
rect 8116 700742 8168 700748
rect 3514 697976 3570 697985
rect 3896 697966 3924 700742
rect 24320 700262 24348 703520
rect 40512 700262 40540 703520
rect 20352 700256 20404 700262
rect 20352 700198 20404 700204
rect 24308 700256 24360 700262
rect 24308 700198 24360 700204
rect 36728 700256 36780 700262
rect 36728 700198 36780 700204
rect 40500 700256 40552 700262
rect 40500 700198 40552 700204
rect 20364 698170 20392 700198
rect 36740 698170 36768 700198
rect 56796 700058 56824 703520
rect 72988 700262 73016 703520
rect 89180 700262 89208 703520
rect 105464 700806 105492 703520
rect 102048 700800 102100 700806
rect 102048 700742 102100 700748
rect 105452 700800 105504 700806
rect 105452 700742 105504 700748
rect 69388 700256 69440 700262
rect 69388 700198 69440 700204
rect 72976 700256 73028 700262
rect 72976 700198 73028 700204
rect 85764 700256 85816 700262
rect 85764 700198 85816 700204
rect 89168 700256 89220 700262
rect 89168 700198 89220 700204
rect 53012 700052 53064 700058
rect 53012 699994 53064 700000
rect 56784 700052 56836 700058
rect 56784 699994 56836 700000
rect 53024 698170 53052 699994
rect 69400 698170 69428 700198
rect 85776 698170 85804 700198
rect 102060 698170 102088 700742
rect 121656 700194 121684 703520
rect 137848 700262 137876 703520
rect 134708 700256 134760 700262
rect 134708 700198 134760 700204
rect 137836 700256 137888 700262
rect 137836 700198 137888 700204
rect 118424 700188 118476 700194
rect 118424 700130 118476 700136
rect 121644 700188 121696 700194
rect 121644 700130 121696 700136
rect 118436 698170 118464 700130
rect 134720 698170 134748 700198
rect 154132 700194 154160 703520
rect 170324 700262 170352 703520
rect 186516 700262 186544 703520
rect 202800 700806 202828 703520
rect 200028 700800 200080 700806
rect 200028 700742 200080 700748
rect 202788 700800 202840 700806
rect 202788 700742 202840 700748
rect 167368 700256 167420 700262
rect 167368 700198 167420 700204
rect 170312 700256 170364 700262
rect 170312 700198 170364 700204
rect 183744 700256 183796 700262
rect 183744 700198 183796 700204
rect 186504 700256 186556 700262
rect 186504 700198 186556 700204
rect 151084 700188 151136 700194
rect 151084 700130 151136 700136
rect 154120 700188 154172 700194
rect 154120 700130 154172 700136
rect 151096 698170 151124 700130
rect 167380 698170 167408 700198
rect 183756 698170 183784 700198
rect 20316 698142 20392 698170
rect 36692 698142 36768 698170
rect 52976 698142 53052 698170
rect 69352 698142 69428 698170
rect 85728 698142 85804 698170
rect 102012 698142 102088 698170
rect 118388 698142 118464 698170
rect 134672 698142 134748 698170
rect 151048 698142 151124 698170
rect 167332 698142 167408 698170
rect 183708 698142 183784 698170
rect 200040 698170 200068 700742
rect 218992 700194 219020 703520
rect 235184 700262 235212 703520
rect 251468 700262 251496 703520
rect 267660 700262 267688 703520
rect 283852 700262 283880 703520
rect 232780 700256 232832 700262
rect 232780 700198 232832 700204
rect 235172 700256 235224 700262
rect 235172 700198 235224 700204
rect 249064 700256 249116 700262
rect 249064 700198 249116 700204
rect 251456 700256 251508 700262
rect 251456 700198 251508 700204
rect 265440 700256 265492 700262
rect 265440 700198 265492 700204
rect 267648 700256 267700 700262
rect 267648 700198 267700 700204
rect 281816 700256 281868 700262
rect 281816 700198 281868 700204
rect 283840 700256 283892 700262
rect 283840 700198 283892 700204
rect 216404 700188 216456 700194
rect 216404 700130 216456 700136
rect 218980 700188 219032 700194
rect 218980 700130 219032 700136
rect 216416 698170 216444 700130
rect 232792 698170 232820 700198
rect 249076 698170 249104 700198
rect 265452 698170 265480 700198
rect 281828 698170 281856 700198
rect 300136 700194 300164 703520
rect 316328 700806 316356 703520
rect 314476 700800 314528 700806
rect 314476 700742 314528 700748
rect 316316 700800 316368 700806
rect 316316 700742 316368 700748
rect 298008 700188 298060 700194
rect 298008 700130 298060 700136
rect 300124 700188 300176 700194
rect 300124 700130 300176 700136
rect 200040 698142 200112 698170
rect 3896 697938 4046 697966
rect 20316 697959 20344 698142
rect 36692 697959 36720 698142
rect 52976 697959 53004 698142
rect 69352 697959 69380 698142
rect 85728 697959 85756 698142
rect 102012 697959 102040 698142
rect 118388 697959 118416 698142
rect 134672 697959 134700 698142
rect 151048 697959 151076 698142
rect 167332 697959 167360 698142
rect 183708 697959 183736 698142
rect 200084 697959 200112 698142
rect 216368 698142 216444 698170
rect 232744 698142 232820 698170
rect 249028 698142 249104 698170
rect 265404 698142 265480 698170
rect 281780 698142 281856 698170
rect 298020 698170 298048 700130
rect 314488 698170 314516 700742
rect 332520 700262 332548 703520
rect 348804 700262 348832 703520
rect 364996 700466 365024 703520
rect 363512 700460 363564 700466
rect 363512 700402 363564 700408
rect 364984 700460 365036 700466
rect 364984 700402 365036 700408
rect 330760 700256 330812 700262
rect 330760 700198 330812 700204
rect 332508 700256 332560 700262
rect 332508 700198 332560 700204
rect 347136 700256 347188 700262
rect 347136 700198 347188 700204
rect 348792 700256 348844 700262
rect 348792 700198 348844 700204
rect 330772 698170 330800 700198
rect 347148 698170 347176 700198
rect 363524 698170 363552 700402
rect 381188 699922 381216 703520
rect 397472 700262 397500 703520
rect 413664 700466 413692 703520
rect 412456 700460 412508 700466
rect 412456 700402 412508 700408
rect 413652 700460 413704 700466
rect 413652 700402 413704 700408
rect 396172 700256 396224 700262
rect 396172 700198 396224 700204
rect 397460 700256 397512 700262
rect 397460 700198 397512 700204
rect 379796 699916 379848 699922
rect 379796 699858 379848 699864
rect 381176 699916 381228 699922
rect 381176 699858 381228 699864
rect 379808 698170 379836 699858
rect 396184 698170 396212 700198
rect 412468 698170 412496 700402
rect 429856 700262 429884 703520
rect 446140 700262 446168 703520
rect 462332 700262 462360 703520
rect 428832 700256 428884 700262
rect 428832 700198 428884 700204
rect 429844 700256 429896 700262
rect 429844 700198 429896 700204
rect 445208 700256 445260 700262
rect 445208 700198 445260 700204
rect 446128 700256 446180 700262
rect 446128 700198 446180 700204
rect 461492 700256 461544 700262
rect 461492 700198 461544 700204
rect 462320 700256 462372 700262
rect 462320 700198 462372 700204
rect 428844 698170 428872 700198
rect 445220 698170 445248 700198
rect 461504 698170 461532 700198
rect 478524 700194 478552 703520
rect 494808 700194 494836 703520
rect 477868 700188 477920 700194
rect 477868 700130 477920 700136
rect 478512 700188 478564 700194
rect 478512 700130 478564 700136
rect 494244 700188 494296 700194
rect 494244 700130 494296 700136
rect 494796 700188 494848 700194
rect 494796 700130 494848 700136
rect 477880 698170 477908 700130
rect 494256 698170 494284 700130
rect 510632 699802 510660 703582
rect 510816 703474 510844 703582
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 511000 703474 511028 703520
rect 510816 703446 511028 703474
rect 527192 699802 527220 703520
rect 543476 702434 543504 703520
rect 559668 702434 559696 703520
rect 510540 699774 510660 699802
rect 526916 699774 527220 699802
rect 543200 702406 543504 702434
rect 559576 702406 559696 702434
rect 510540 698170 510568 699774
rect 526916 698170 526944 699774
rect 543200 698170 543228 702406
rect 559576 698170 559604 702406
rect 298020 698142 298092 698170
rect 216368 697959 216396 698142
rect 232744 697959 232772 698142
rect 249028 697959 249056 698142
rect 265404 697959 265432 698142
rect 281780 697959 281808 698142
rect 298064 697959 298092 698142
rect 314440 698142 314516 698170
rect 330724 698142 330800 698170
rect 347100 698142 347176 698170
rect 363476 698142 363552 698170
rect 379760 698142 379836 698170
rect 396136 698142 396212 698170
rect 412420 698142 412496 698170
rect 428796 698142 428872 698170
rect 445172 698142 445248 698170
rect 461456 698142 461532 698170
rect 477832 698142 477908 698170
rect 494208 698142 494284 698170
rect 510492 698142 510568 698170
rect 526868 698142 526944 698170
rect 543152 698142 543228 698170
rect 559528 698142 559604 698170
rect 575860 698170 575888 703520
rect 575860 698142 575932 698170
rect 314440 697959 314468 698142
rect 330724 697959 330752 698142
rect 347100 697959 347128 698142
rect 363476 697959 363504 698142
rect 379760 697959 379788 698142
rect 396136 697959 396164 698142
rect 412420 697959 412448 698142
rect 428796 697959 428824 698142
rect 445172 697959 445200 698142
rect 461456 697959 461484 698142
rect 477832 697959 477860 698142
rect 494208 697959 494236 698142
rect 510492 697959 510520 698142
rect 526868 697959 526896 698142
rect 543152 697959 543180 698142
rect 559528 697959 559556 698142
rect 575904 697959 575932 698142
rect 3514 697911 3570 697920
rect 3528 697377 3556 697911
rect 3514 697368 3570 697377
rect 3514 697303 3570 697312
rect 579526 684720 579582 684729
rect 579582 684678 579660 684706
rect 579526 684655 579582 684664
rect 579632 683913 579660 684678
rect 579618 683904 579674 683913
rect 579618 683839 579674 683848
rect 578330 644600 578386 644609
rect 578330 644535 578332 644544
rect 578384 644535 578386 644544
rect 580908 644564 580960 644570
rect 578332 644506 578384 644512
rect 580908 644506 580960 644512
rect 580920 644065 580948 644506
rect 580906 644056 580962 644065
rect 580906 643991 580962 644000
rect 3422 436656 3478 436665
rect 3422 436591 3478 436600
rect 3436 436051 3464 436591
rect 3422 436042 3478 436051
rect 3422 435977 3478 435986
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3436 422997 3464 423535
rect 3422 422988 3478 422997
rect 3422 422923 3478 422932
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 3436 409943 3464 410479
rect 3422 409934 3478 409943
rect 3422 409869 3478 409878
rect 3422 397488 3478 397497
rect 3422 397423 3478 397432
rect 3436 396889 3464 397423
rect 3422 396880 3478 396889
rect 3422 396815 3478 396824
rect 3422 384432 3478 384441
rect 3422 384367 3478 384376
rect 3436 383713 3464 384367
rect 3422 383704 3478 383713
rect 3422 383639 3478 383648
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 3436 370659 3464 371311
rect 3422 370650 3478 370659
rect 3422 370585 3478 370594
rect 3422 358456 3478 358465
rect 3422 358391 3478 358400
rect 3436 357605 3464 358391
rect 3422 357596 3478 357605
rect 3422 357531 3478 357540
rect 579526 351928 579582 351937
rect 579526 351863 579582 351872
rect 579540 351121 579568 351863
rect 579526 351112 579582 351121
rect 579526 351047 579582 351056
rect 3422 345400 3478 345409
rect 3422 345335 3478 345344
rect 3436 344429 3464 345335
rect 3422 344420 3478 344429
rect 3422 344355 3478 344364
rect 579618 338600 579674 338609
rect 579618 338535 579674 338544
rect 579526 337920 579582 337929
rect 579632 337906 579660 338535
rect 579582 337878 579660 337906
rect 579526 337855 579582 337864
rect 3422 332344 3478 332353
rect 3422 332279 3478 332288
rect 3436 331375 3464 332279
rect 3422 331366 3478 331375
rect 3422 331301 3478 331310
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324465 580212 325207
rect 580170 324456 580226 324465
rect 580170 324391 580226 324400
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 318321 3464 319223
rect 3422 318312 3478 318321
rect 3422 318247 3478 318256
rect 579618 312080 579674 312089
rect 579618 312015 579674 312024
rect 579526 311128 579582 311137
rect 579632 311114 579660 312015
rect 579582 311086 579660 311114
rect 579526 311063 579582 311072
rect 3422 306232 3478 306241
rect 3422 306167 3478 306176
rect 3436 305145 3464 306167
rect 3422 305136 3478 305145
rect 3422 305071 3478 305080
rect 579618 298752 579674 298761
rect 579618 298687 579674 298696
rect 579526 297800 579582 297809
rect 579632 297786 579660 298687
rect 579582 297758 579660 297786
rect 579526 297735 579582 297744
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 3436 292091 3464 293111
rect 3422 292082 3478 292091
rect 3422 292017 3478 292026
rect 580170 285424 580226 285433
rect 580170 285359 580226 285368
rect 580184 284481 580212 285359
rect 580170 284472 580226 284481
rect 580170 284407 580226 284416
rect 3422 280120 3478 280129
rect 3422 280055 3478 280064
rect 3436 279037 3464 280055
rect 3422 279028 3478 279037
rect 3422 278963 3478 278972
rect 579618 272232 579674 272241
rect 579618 272167 579674 272176
rect 579526 271144 579582 271153
rect 579632 271130 579660 272167
rect 579582 271102 579660 271130
rect 579526 271079 579582 271088
rect 3422 267200 3478 267209
rect 3422 267135 3478 267144
rect 3436 265983 3464 267135
rect 3422 265974 3478 265983
rect 3422 265909 3478 265918
rect 580906 258904 580962 258913
rect 580906 258839 580962 258848
rect 580920 257854 580948 258839
rect 578884 257848 578936 257854
rect 578884 257790 578936 257796
rect 580908 257848 580960 257854
rect 580908 257790 580960 257796
rect 578896 257689 578924 257790
rect 578882 257680 578938 257689
rect 578882 257615 578938 257624
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3436 252807 3464 254079
rect 3422 252798 3478 252807
rect 3422 252733 3478 252742
rect 580170 245576 580226 245585
rect 580170 245511 580226 245520
rect 580184 244497 580212 245511
rect 580170 244488 580226 244497
rect 580170 244423 580226 244432
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 3436 239753 3464 241023
rect 3422 239744 3478 239753
rect 3422 239679 3478 239688
rect 579618 232384 579674 232393
rect 579618 232319 579674 232328
rect 579526 231160 579582 231169
rect 579632 231146 579660 232319
rect 579582 231118 579660 231146
rect 579526 231095 579582 231104
rect 3422 228032 3478 228041
rect 3422 227967 3478 227976
rect 3436 226699 3464 227967
rect 3422 226690 3478 226699
rect 3422 226625 3478 226634
rect 579618 219056 579674 219065
rect 579618 218991 579674 219000
rect 579526 217696 579582 217705
rect 579632 217682 579660 218991
rect 579582 217654 579660 217682
rect 579526 217631 579582 217640
rect 3422 214976 3478 214985
rect 3422 214911 3478 214920
rect 3436 213523 3464 214911
rect 3422 213514 3478 213523
rect 3422 213449 3478 213458
rect 579618 205728 579674 205737
rect 579618 205663 579674 205672
rect 579526 204368 579582 204377
rect 579632 204354 579660 205663
rect 579582 204326 579660 204354
rect 579526 204303 579582 204312
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 3436 200469 3464 201855
rect 3422 200460 3478 200469
rect 3422 200395 3478 200404
rect 579618 192536 579674 192545
rect 579618 192471 579674 192480
rect 579526 191040 579582 191049
rect 579632 191026 579660 192471
rect 579582 190998 579660 191026
rect 579526 190975 579582 190984
rect 3606 188864 3662 188873
rect 3606 188799 3662 188808
rect 3620 187415 3648 188799
rect 3606 187406 3662 187415
rect 3606 187341 3662 187350
rect 579618 179208 579674 179217
rect 579618 179143 579674 179152
rect 579526 177712 579582 177721
rect 579632 177698 579660 179143
rect 579582 177670 579660 177698
rect 579526 177647 579582 177656
rect 3422 175944 3478 175953
rect 3422 175879 3478 175888
rect 3436 174239 3464 175879
rect 3422 174230 3478 174239
rect 3422 174165 3478 174174
rect 579618 165880 579674 165889
rect 579618 165815 579674 165824
rect 579526 164384 579582 164393
rect 579632 164370 579660 165815
rect 579582 164342 579660 164370
rect 579526 164319 579582 164328
rect 2134 162888 2190 162897
rect 2134 162823 2190 162832
rect 2148 161129 2176 162823
rect 2134 161120 2190 161129
rect 2134 161055 2190 161064
rect 580906 152688 580962 152697
rect 580906 152623 580962 152632
rect 580920 151502 580948 152623
rect 578516 151496 578568 151502
rect 578516 151438 578568 151444
rect 580908 151496 580960 151502
rect 580908 151438 580960 151444
rect 578528 151065 578556 151438
rect 578514 151056 578570 151065
rect 578514 150991 578570 151000
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3436 148131 3464 149767
rect 3422 148122 3478 148131
rect 3422 148057 3478 148066
rect 579618 139360 579674 139369
rect 579618 139295 579674 139304
rect 579526 137592 579582 137601
rect 579632 137578 579660 139295
rect 579582 137550 579660 137578
rect 579526 137527 579582 137536
rect 2134 136776 2190 136785
rect 2134 136711 2190 136720
rect 2148 135017 2176 136711
rect 2134 135008 2190 135017
rect 2134 134943 2190 134952
rect 579618 126032 579674 126041
rect 579618 125967 579674 125976
rect 579526 124400 579582 124409
rect 579632 124386 579660 125967
rect 579582 124358 579660 124386
rect 579526 124335 579582 124344
rect 3422 123720 3478 123729
rect 3422 123655 3478 123664
rect 3436 121901 3464 123655
rect 3422 121892 3478 121901
rect 3422 121827 3478 121836
rect 579618 112840 579674 112849
rect 579618 112775 579674 112784
rect 579526 110936 579582 110945
rect 579632 110922 579660 112775
rect 579582 110894 579660 110922
rect 579526 110871 579582 110880
rect 2134 110664 2190 110673
rect 2134 110599 2190 110608
rect 2148 108905 2176 110599
rect 2134 108896 2190 108905
rect 2134 108831 2190 108840
rect 579618 99512 579674 99521
rect 579618 99447 579674 99456
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 579526 97608 579582 97617
rect 579632 97594 579660 99447
rect 579582 97566 579660 97594
rect 579526 97543 579582 97552
rect 3436 95793 3464 97543
rect 3422 95784 3478 95793
rect 3422 95719 3478 95728
rect 579618 86184 579674 86193
rect 579618 86119 579674 86128
rect 2134 84688 2190 84697
rect 2134 84623 2190 84632
rect 2148 82657 2176 84623
rect 579526 84280 579582 84289
rect 579632 84266 579660 86119
rect 579582 84238 579660 84266
rect 579526 84215 579582 84224
rect 2134 82648 2190 82657
rect 2134 82583 2190 82592
rect 579618 72992 579674 73001
rect 579618 72927 579674 72936
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3436 69563 3464 71567
rect 579526 70952 579582 70961
rect 579632 70938 579660 72927
rect 579582 70910 579660 70938
rect 579526 70887 579582 70896
rect 3422 69554 3478 69563
rect 3422 69489 3478 69498
rect 579618 59664 579674 59673
rect 579618 59599 579674 59608
rect 2134 58576 2190 58585
rect 2134 58511 2190 58520
rect 2148 56545 2176 58511
rect 579526 57624 579582 57633
rect 579632 57610 579660 59599
rect 579582 57582 579660 57610
rect 579526 57559 579582 57568
rect 2134 56536 2190 56545
rect 2134 56471 2190 56480
rect 579986 46336 580042 46345
rect 579986 46271 580042 46280
rect 3422 45520 3478 45529
rect 3422 45455 3478 45464
rect 3436 43333 3464 45455
rect 580000 45014 580028 46271
rect 578332 45008 578384 45014
rect 578332 44950 578384 44956
rect 579988 45008 580040 45014
rect 579988 44950 580040 44956
rect 578344 44305 578372 44950
rect 578330 44296 578386 44305
rect 578330 44231 578386 44240
rect 3422 43324 3478 43333
rect 3422 43259 3478 43268
rect 579618 33144 579674 33153
rect 579618 33079 579674 33088
rect 2134 32464 2190 32473
rect 2134 32399 2190 32408
rect 2148 30297 2176 32399
rect 579526 30968 579582 30977
rect 579632 30954 579660 33079
rect 579582 30926 579660 30954
rect 579526 30903 579582 30912
rect 2134 30288 2190 30297
rect 2134 30223 2190 30232
rect 579618 19816 579674 19825
rect 579618 19751 579674 19760
rect 2042 19408 2098 19417
rect 2042 19343 2098 19352
rect 2056 17241 2084 19343
rect 579526 17640 579582 17649
rect 579632 17626 579660 19751
rect 579582 17598 579660 17626
rect 579526 17575 579582 17584
rect 2042 17232 2098 17241
rect 2042 17167 2098 17176
rect 579618 6624 579674 6633
rect 579618 6559 579674 6568
rect 2778 6488 2834 6497
rect 2778 6423 2834 6432
rect 2792 4185 2820 6423
rect 2778 4176 2834 4185
rect 2778 4111 2834 4120
rect 579526 4176 579582 4185
rect 579632 4162 579660 6559
rect 579582 4134 579660 4162
rect 579526 4111 579582 4120
rect 1676 3868 1728 3874
rect 1676 3810 1728 3816
rect 572 3800 624 3806
rect 572 3742 624 3748
rect 584 480 612 3742
rect 1688 480 1716 3810
rect 4124 3806 4152 4012
rect 5228 3874 5256 4012
rect 5216 3868 5268 3874
rect 5216 3810 5268 3816
rect 4112 3800 4164 3806
rect 6424 3754 6452 4012
rect 7528 3754 7556 4012
rect 4112 3742 4164 3748
rect 6380 3726 6452 3754
rect 7484 3726 7556 3754
rect 7656 3800 7708 3806
rect 8724 3754 8752 4012
rect 9920 3754 9948 4012
rect 11024 3806 11052 4012
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 7656 3742 7708 3748
rect 4068 2916 4120 2922
rect 4068 2858 4120 2864
rect 3240 1352 3292 1358
rect 3240 1294 3292 1300
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 354 2954 480
rect 3252 354 3280 1294
rect 4080 480 4108 2858
rect 6380 1358 6408 3726
rect 7484 2922 7512 3726
rect 7472 2916 7524 2922
rect 7472 2858 7524 2864
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 6368 1352 6420 1358
rect 6368 1294 6420 1300
rect 5632 1148 5684 1154
rect 5632 1090 5684 1096
rect 2842 326 3280 354
rect 2842 -960 2954 326
rect 4038 -960 4150 480
rect 5234 354 5346 480
rect 5644 354 5672 1090
rect 6472 480 6500 2790
rect 7668 480 7696 3742
rect 8680 3726 8752 3754
rect 9876 3726 9948 3754
rect 11012 3800 11064 3806
rect 11012 3742 11064 3748
rect 8680 1154 8708 3726
rect 9876 2854 9904 3726
rect 9864 2848 9916 2854
rect 9864 2790 9916 2796
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 8668 1148 8720 1154
rect 8668 1090 8720 1096
rect 8760 944 8812 950
rect 8760 886 8812 892
rect 8772 480 8800 886
rect 9968 480 9996 2790
rect 11164 480 11192 3878
rect 12220 3754 12248 4012
rect 12176 3726 12248 3754
rect 12348 3800 12400 3806
rect 13324 3754 13352 4012
rect 14520 3942 14548 4012
rect 14508 3936 14560 3942
rect 14508 3878 14560 3884
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 13544 3868 13596 3874
rect 13544 3810 13596 3816
rect 12348 3742 12400 3748
rect 12176 950 12204 3726
rect 12164 944 12216 950
rect 12164 886 12216 892
rect 12360 480 12388 3742
rect 13280 3726 13352 3754
rect 13280 2854 13308 3726
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 13556 480 13584 3810
rect 14752 480 14780 3878
rect 15716 3806 15744 4012
rect 16820 3874 16848 4012
rect 18016 3942 18044 4012
rect 18004 3936 18056 3942
rect 18004 3878 18056 3884
rect 16808 3868 16860 3874
rect 16808 3810 16860 3816
rect 19120 3806 19148 4012
rect 19432 3868 19484 3874
rect 19432 3810 19484 3816
rect 15704 3800 15756 3806
rect 15704 3742 15756 3748
rect 15936 3800 15988 3806
rect 15936 3742 15988 3748
rect 19108 3800 19160 3806
rect 19108 3742 19160 3748
rect 15948 480 15976 3742
rect 18236 2916 18288 2922
rect 18236 2858 18288 2864
rect 17040 2848 17092 2854
rect 17040 2790 17092 2796
rect 17052 480 17080 2790
rect 18248 480 18276 2858
rect 19444 480 19472 3810
rect 20316 3754 20344 4012
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 20272 3726 20344 3754
rect 20272 2854 20300 3726
rect 20260 2848 20312 2854
rect 20260 2790 20312 2796
rect 20640 480 20668 3878
rect 21512 3754 21540 4012
rect 22616 3874 22644 4012
rect 23812 3942 23840 4012
rect 23800 3936 23852 3942
rect 23800 3878 23852 3884
rect 24216 3936 24268 3942
rect 24216 3878 24268 3884
rect 22604 3868 22656 3874
rect 22604 3810 22656 3816
rect 23020 3868 23072 3874
rect 23020 3810 23072 3816
rect 21468 3726 21540 3754
rect 21824 3800 21876 3806
rect 21824 3742 21876 3748
rect 21468 2922 21496 3726
rect 21456 2916 21508 2922
rect 21456 2858 21508 2864
rect 21836 480 21864 3742
rect 23032 480 23060 3810
rect 24228 480 24256 3878
rect 24916 3806 24944 4012
rect 26112 3874 26140 4012
rect 27308 3942 27336 4012
rect 27296 3936 27348 3942
rect 27296 3878 27348 3884
rect 27712 3936 27764 3942
rect 27712 3878 27764 3884
rect 26100 3868 26152 3874
rect 26100 3810 26152 3816
rect 26516 3868 26568 3874
rect 26516 3810 26568 3816
rect 24904 3800 24956 3806
rect 24904 3742 24956 3748
rect 25320 3800 25372 3806
rect 25320 3742 25372 3748
rect 25332 480 25360 3742
rect 26528 480 26556 3810
rect 27724 480 27752 3878
rect 28412 3806 28440 4012
rect 29608 3874 29636 4012
rect 30712 3942 30740 4012
rect 30700 3936 30752 3942
rect 30700 3878 30752 3884
rect 29596 3868 29648 3874
rect 29596 3810 29648 3816
rect 30104 3868 30156 3874
rect 30104 3810 30156 3816
rect 28400 3800 28452 3806
rect 28400 3742 28452 3748
rect 28908 2848 28960 2854
rect 28908 2790 28960 2796
rect 28920 480 28948 2790
rect 30116 480 30144 3810
rect 31300 3800 31352 3806
rect 31908 3754 31936 4012
rect 32404 3936 32456 3942
rect 32404 3878 32456 3884
rect 31300 3742 31352 3748
rect 31312 480 31340 3742
rect 31864 3726 31936 3754
rect 31864 2854 31892 3726
rect 31852 2848 31904 2854
rect 31852 2790 31904 2796
rect 32416 480 32444 3878
rect 33104 3874 33132 4012
rect 33092 3868 33144 3874
rect 33092 3810 33144 3816
rect 33600 3868 33652 3874
rect 33600 3810 33652 3816
rect 33612 480 33640 3810
rect 34208 3806 34236 4012
rect 35404 3942 35432 4012
rect 35392 3936 35444 3942
rect 35392 3878 35444 3884
rect 36600 3874 36628 4012
rect 36588 3868 36640 3874
rect 36588 3810 36640 3816
rect 37188 3868 37240 3874
rect 37188 3810 37240 3816
rect 34196 3800 34248 3806
rect 34196 3742 34248 3748
rect 34796 3800 34848 3806
rect 34796 3742 34848 3748
rect 34808 480 34836 3742
rect 35992 2848 36044 2854
rect 35992 2790 36044 2796
rect 36004 480 36032 2790
rect 37200 480 37228 3810
rect 37704 3806 37732 4012
rect 38384 3936 38436 3942
rect 38384 3878 38436 3884
rect 37692 3800 37744 3806
rect 37692 3742 37744 3748
rect 38396 480 38424 3878
rect 38900 3754 38928 4012
rect 40004 3874 40032 4012
rect 41200 3942 41228 4012
rect 41188 3936 41240 3942
rect 41188 3878 41240 3884
rect 39992 3868 40044 3874
rect 39992 3810 40044 3816
rect 41880 3868 41932 3874
rect 41880 3810 41932 3816
rect 38856 3726 38928 3754
rect 40684 3800 40736 3806
rect 40684 3742 40736 3748
rect 38856 2854 38884 3726
rect 38844 2848 38896 2854
rect 38844 2790 38896 2796
rect 39580 2848 39632 2854
rect 39580 2790 39632 2796
rect 39592 480 39620 2790
rect 40696 480 40724 3742
rect 41892 480 41920 3810
rect 42396 3754 42424 4012
rect 43076 3936 43128 3942
rect 43076 3878 43128 3884
rect 42352 3726 42424 3754
rect 42352 2854 42380 3726
rect 42340 2848 42392 2854
rect 42340 2790 42392 2796
rect 43088 480 43116 3878
rect 43500 3806 43528 4012
rect 44696 3874 44724 4012
rect 45800 3942 45828 4012
rect 45788 3936 45840 3942
rect 45788 3878 45840 3884
rect 46664 3936 46716 3942
rect 46664 3878 46716 3884
rect 44684 3868 44736 3874
rect 44684 3810 44736 3816
rect 45468 3868 45520 3874
rect 45468 3810 45520 3816
rect 43488 3800 43540 3806
rect 43488 3742 43540 3748
rect 44272 3800 44324 3806
rect 44272 3742 44324 3748
rect 44284 480 44312 3742
rect 45480 480 45508 3810
rect 46676 480 46704 3878
rect 46996 3806 47024 4012
rect 48192 3874 48220 4012
rect 49296 3942 49324 4012
rect 49284 3936 49336 3942
rect 49284 3878 49336 3884
rect 50160 3936 50212 3942
rect 50160 3878 50212 3884
rect 48180 3868 48232 3874
rect 48180 3810 48232 3816
rect 48964 3868 49016 3874
rect 48964 3810 49016 3816
rect 46984 3800 47036 3806
rect 46984 3742 47036 3748
rect 47860 3800 47912 3806
rect 47860 3742 47912 3748
rect 47872 480 47900 3742
rect 48976 480 49004 3810
rect 50172 480 50200 3878
rect 50492 3806 50520 4012
rect 51596 3874 51624 4012
rect 52792 3942 52820 4012
rect 52780 3936 52832 3942
rect 52780 3878 52832 3884
rect 51584 3868 51636 3874
rect 51584 3810 51636 3816
rect 53748 3868 53800 3874
rect 53748 3810 53800 3816
rect 50480 3800 50532 3806
rect 50480 3742 50532 3748
rect 51356 3800 51408 3806
rect 51356 3742 51408 3748
rect 51368 480 51396 3742
rect 52552 740 52604 746
rect 52552 682 52604 688
rect 52564 480 52592 682
rect 53760 480 53788 3810
rect 53988 3806 54016 4012
rect 53976 3800 54028 3806
rect 53976 3742 54028 3748
rect 54944 3800 54996 3806
rect 55092 3754 55120 4012
rect 56048 3936 56100 3942
rect 56048 3878 56100 3884
rect 54944 3742 54996 3748
rect 54956 480 54984 3742
rect 55048 3726 55120 3754
rect 55048 746 55076 3726
rect 55036 740 55088 746
rect 55036 682 55088 688
rect 56060 480 56088 3878
rect 56288 3874 56316 4012
rect 56276 3868 56328 3874
rect 56276 3810 56328 3816
rect 57244 3868 57296 3874
rect 57244 3810 57296 3816
rect 57256 480 57284 3810
rect 57392 3806 57420 4012
rect 58588 3942 58616 4012
rect 58576 3936 58628 3942
rect 58576 3878 58628 3884
rect 59784 3874 59812 4012
rect 59772 3868 59824 3874
rect 59772 3810 59824 3816
rect 60888 3806 60916 4012
rect 62084 3890 62112 4012
rect 61948 3862 62112 3890
rect 57380 3800 57432 3806
rect 57380 3742 57432 3748
rect 58440 3800 58492 3806
rect 58440 3742 58492 3748
rect 60876 3800 60928 3806
rect 60876 3742 60928 3748
rect 58452 480 58480 3742
rect 60832 1352 60884 1358
rect 60832 1294 60884 1300
rect 59636 740 59688 746
rect 59636 682 59688 688
rect 59648 480 59676 682
rect 60844 480 60872 1294
rect 61948 746 61976 3862
rect 63280 3754 63308 4012
rect 64384 3890 64412 4012
rect 64384 3862 64460 3890
rect 64328 3800 64380 3806
rect 63280 3726 63356 3754
rect 64328 3742 64380 3748
rect 63224 3052 63276 3058
rect 63224 2994 63276 3000
rect 62028 2848 62080 2854
rect 62028 2790 62080 2796
rect 61936 740 61988 746
rect 61936 682 61988 688
rect 62040 480 62068 2790
rect 63236 480 63264 2994
rect 63328 1358 63356 3726
rect 63316 1352 63368 1358
rect 63316 1294 63368 1300
rect 64340 480 64368 3742
rect 64432 2854 64460 3862
rect 65580 3754 65608 4012
rect 66684 3806 66712 4012
rect 65536 3726 65608 3754
rect 66672 3800 66724 3806
rect 66672 3742 66724 3748
rect 67088 3800 67140 3806
rect 67880 3754 67908 4012
rect 69076 3806 69104 4012
rect 67088 3742 67140 3748
rect 65536 3058 65564 3726
rect 65524 3052 65576 3058
rect 65524 2994 65576 3000
rect 64420 2848 64472 2854
rect 64420 2790 64472 2796
rect 65524 2848 65576 2854
rect 65524 2790 65576 2796
rect 65536 480 65564 2790
rect 5234 326 5672 354
rect 5234 -960 5346 326
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 218 66802 480
rect 67100 218 67128 3742
rect 67836 3726 67908 3754
rect 69064 3800 69116 3806
rect 70180 3754 70208 4012
rect 69064 3742 69116 3748
rect 70136 3726 70208 3754
rect 70308 3800 70360 3806
rect 71376 3754 71404 4012
rect 71504 3868 71556 3874
rect 71504 3810 71556 3816
rect 70308 3742 70360 3748
rect 67836 2854 67864 3726
rect 67824 2848 67876 2854
rect 67824 2790 67876 2796
rect 70136 1358 70164 3726
rect 67916 1352 67968 1358
rect 67916 1294 67968 1300
rect 70124 1352 70176 1358
rect 70124 1294 70176 1300
rect 67928 480 67956 1294
rect 69112 604 69164 610
rect 69112 546 69164 552
rect 69124 480 69152 546
rect 70320 480 70348 3742
rect 71332 3726 71404 3754
rect 71332 610 71360 3726
rect 71320 604 71372 610
rect 71320 546 71372 552
rect 71516 480 71544 3810
rect 72480 3806 72508 4012
rect 72608 3936 72660 3942
rect 72608 3878 72660 3884
rect 72468 3800 72520 3806
rect 72468 3742 72520 3748
rect 72620 480 72648 3878
rect 73676 3874 73704 4012
rect 74872 3942 74900 4012
rect 74860 3936 74912 3942
rect 74860 3878 74912 3884
rect 73664 3868 73716 3874
rect 73664 3810 73716 3816
rect 75976 3806 76004 4012
rect 73804 3800 73856 3806
rect 73804 3742 73856 3748
rect 75964 3800 76016 3806
rect 77172 3754 77200 4012
rect 78276 3754 78304 4012
rect 78588 3868 78640 3874
rect 78588 3810 78640 3816
rect 75964 3742 76016 3748
rect 73816 480 73844 3742
rect 77128 3726 77200 3754
rect 78232 3726 78304 3754
rect 76196 1352 76248 1358
rect 76196 1294 76248 1300
rect 75000 1284 75052 1290
rect 75000 1226 75052 1232
rect 75012 480 75040 1226
rect 76208 480 76236 1294
rect 77128 1290 77156 3726
rect 78232 1358 78260 3726
rect 78220 1352 78272 1358
rect 78220 1294 78272 1300
rect 77116 1284 77168 1290
rect 77116 1226 77168 1232
rect 77392 1284 77444 1290
rect 77392 1226 77444 1232
rect 77404 480 77432 1226
rect 78600 480 78628 3810
rect 79472 3754 79500 4012
rect 80668 3874 80696 4012
rect 80656 3868 80708 3874
rect 80656 3810 80708 3816
rect 80888 3868 80940 3874
rect 80888 3810 80940 3816
rect 79428 3726 79500 3754
rect 79692 3800 79744 3806
rect 79692 3742 79744 3748
rect 79428 1290 79456 3726
rect 79416 1284 79468 1290
rect 79416 1226 79468 1232
rect 79704 480 79732 3742
rect 80900 480 80928 3810
rect 81772 3806 81800 4012
rect 82968 3874 82996 4012
rect 82956 3868 83008 3874
rect 82956 3810 83008 3816
rect 81760 3800 81812 3806
rect 84072 3754 84100 4012
rect 85268 3754 85296 4012
rect 86464 3754 86492 4012
rect 81760 3742 81812 3748
rect 84028 3726 84100 3754
rect 85224 3726 85296 3754
rect 86420 3726 86492 3754
rect 86868 3800 86920 3806
rect 87568 3754 87596 4012
rect 87972 3868 88024 3874
rect 87972 3810 88024 3816
rect 86868 3742 86920 3748
rect 83280 1352 83332 1358
rect 83280 1294 83332 1300
rect 82084 1284 82136 1290
rect 82084 1226 82136 1232
rect 82096 480 82124 1226
rect 83292 480 83320 1294
rect 84028 1290 84056 3726
rect 85224 1358 85252 3726
rect 85212 1352 85264 1358
rect 85212 1294 85264 1300
rect 85672 1352 85724 1358
rect 85672 1294 85724 1300
rect 84016 1284 84068 1290
rect 84016 1226 84068 1232
rect 84476 1284 84528 1290
rect 84476 1226 84528 1232
rect 84488 480 84516 1226
rect 85684 480 85712 1294
rect 86420 1290 86448 3726
rect 86408 1284 86460 1290
rect 86408 1226 86460 1232
rect 86880 480 86908 3742
rect 87524 3726 87596 3754
rect 87524 1358 87552 3726
rect 87512 1352 87564 1358
rect 87512 1294 87564 1300
rect 87984 480 88012 3810
rect 88764 3806 88792 4012
rect 89960 3874 89988 4012
rect 89948 3868 90000 3874
rect 89948 3810 90000 3816
rect 88752 3800 88804 3806
rect 91064 3754 91092 4012
rect 92260 3754 92288 4012
rect 93364 3754 93392 4012
rect 94560 3754 94588 4012
rect 88752 3742 88804 3748
rect 91020 3726 91092 3754
rect 92216 3726 92288 3754
rect 93320 3726 93392 3754
rect 94516 3726 94588 3754
rect 95148 3800 95200 3806
rect 95756 3754 95784 4012
rect 96252 3868 96304 3874
rect 96252 3810 96304 3816
rect 95148 3742 95200 3748
rect 91020 1358 91048 3726
rect 89168 1352 89220 1358
rect 89168 1294 89220 1300
rect 91008 1352 91060 1358
rect 91008 1294 91060 1300
rect 91560 1352 91612 1358
rect 91560 1294 91612 1300
rect 89180 480 89208 1294
rect 90364 1284 90416 1290
rect 90364 1226 90416 1232
rect 90376 480 90404 1226
rect 91572 480 91600 1294
rect 92216 1290 92244 3726
rect 93320 1358 93348 3726
rect 93308 1352 93360 1358
rect 93308 1294 93360 1300
rect 93952 1352 94004 1358
rect 93952 1294 94004 1300
rect 92204 1284 92256 1290
rect 92204 1226 92256 1232
rect 92756 1284 92808 1290
rect 92756 1226 92808 1232
rect 92768 480 92796 1226
rect 93964 480 93992 1294
rect 94516 1290 94544 3726
rect 94504 1284 94556 1290
rect 94504 1226 94556 1232
rect 95160 480 95188 3742
rect 95712 3726 95784 3754
rect 95712 1358 95740 3726
rect 95700 1352 95752 1358
rect 95700 1294 95752 1300
rect 96264 480 96292 3810
rect 96860 3806 96888 4012
rect 98056 3874 98084 4012
rect 98044 3868 98096 3874
rect 98044 3810 98096 3816
rect 96848 3800 96900 3806
rect 99160 3754 99188 4012
rect 100356 3754 100384 4012
rect 101552 3754 101580 4012
rect 102656 3754 102684 4012
rect 96848 3742 96900 3748
rect 99116 3726 99188 3754
rect 100312 3726 100384 3754
rect 101508 3726 101580 3754
rect 102612 3726 102684 3754
rect 103336 3800 103388 3806
rect 103852 3754 103880 4012
rect 104956 3806 104984 4012
rect 103336 3742 103388 3748
rect 99116 1358 99144 3726
rect 97448 1352 97500 1358
rect 97448 1294 97500 1300
rect 99104 1352 99156 1358
rect 99104 1294 99156 1300
rect 97460 480 97488 1294
rect 100312 1290 100340 3726
rect 101036 1352 101088 1358
rect 101036 1294 101088 1300
rect 98644 1284 98696 1290
rect 98644 1226 98696 1232
rect 100300 1284 100352 1290
rect 100300 1226 100352 1232
rect 98656 480 98684 1226
rect 99840 1216 99892 1222
rect 99840 1158 99892 1164
rect 99852 480 99880 1158
rect 101048 480 101076 1294
rect 101508 1222 101536 3726
rect 102612 1358 102640 3726
rect 102600 1352 102652 1358
rect 102600 1294 102652 1300
rect 102232 1284 102284 1290
rect 102232 1226 102284 1232
rect 101496 1216 101548 1222
rect 101496 1158 101548 1164
rect 102244 480 102272 1226
rect 103348 480 103376 3742
rect 103808 3726 103880 3754
rect 104944 3800 104996 3806
rect 106152 3754 106180 4012
rect 107348 3754 107376 4012
rect 108452 3754 108480 4012
rect 109648 3754 109676 4012
rect 110752 3754 110780 4012
rect 111948 3754 111976 4012
rect 113144 3754 113172 4012
rect 114248 3754 114276 4012
rect 115444 3754 115472 4012
rect 116640 3754 116668 4012
rect 117744 3754 117772 4012
rect 118940 3754 118968 4012
rect 120044 3754 120072 4012
rect 121240 3754 121268 4012
rect 122436 3754 122464 4012
rect 123540 3754 123568 4012
rect 104944 3742 104996 3748
rect 106108 3726 106180 3754
rect 107304 3726 107376 3754
rect 108408 3726 108480 3754
rect 109604 3726 109676 3754
rect 110708 3726 110780 3754
rect 111904 3726 111976 3754
rect 113100 3726 113172 3754
rect 114204 3726 114276 3754
rect 115400 3726 115472 3754
rect 116596 3726 116668 3754
rect 117700 3726 117772 3754
rect 118896 3726 118968 3754
rect 119264 3726 120072 3754
rect 121196 3726 121268 3754
rect 122392 3726 122464 3754
rect 123496 3726 123568 3754
rect 124736 3754 124764 4012
rect 125840 3754 125868 4012
rect 127036 3754 127064 4012
rect 128232 3754 128260 4012
rect 129336 3754 129364 4012
rect 130532 3754 130560 4012
rect 131636 3754 131664 4012
rect 132832 3754 132860 4012
rect 134028 3754 134056 4012
rect 135132 3754 135160 4012
rect 136328 3754 136356 4012
rect 137432 3754 137460 4012
rect 138628 3754 138656 4012
rect 139824 3754 139852 4012
rect 140928 3754 140956 4012
rect 142124 3754 142152 4012
rect 143320 3754 143348 4012
rect 144424 3754 144452 4012
rect 145620 3754 145648 4012
rect 146724 3754 146752 4012
rect 147920 3754 147948 4012
rect 149116 3754 149144 4012
rect 150220 3754 150248 4012
rect 151416 3754 151444 4012
rect 152520 3754 152548 4012
rect 153716 3754 153744 4012
rect 154912 3754 154940 4012
rect 156016 3754 156044 4012
rect 157212 3754 157240 4012
rect 158316 3754 158344 4012
rect 159512 3754 159540 4012
rect 160708 3754 160736 4012
rect 161812 3754 161840 4012
rect 163008 3754 163036 4012
rect 164112 3754 164140 4012
rect 165308 3754 165336 4012
rect 166504 3754 166532 4012
rect 167608 3754 167636 4012
rect 168804 3754 168832 4012
rect 170000 3754 170028 4012
rect 171104 3754 171132 4012
rect 172300 3754 172328 4012
rect 173404 3754 173432 4012
rect 174600 3754 174628 4012
rect 175796 3754 175824 4012
rect 176900 3754 176928 4012
rect 178096 3754 178124 4012
rect 179200 3754 179228 4012
rect 124736 3726 124812 3754
rect 103808 1290 103836 3726
rect 106108 1358 106136 3726
rect 104532 1352 104584 1358
rect 104532 1294 104584 1300
rect 106096 1352 106148 1358
rect 106096 1294 106148 1300
rect 106924 1352 106976 1358
rect 106924 1294 106976 1300
rect 103796 1284 103848 1290
rect 103796 1226 103848 1232
rect 104544 480 104572 1294
rect 105728 740 105780 746
rect 105728 682 105780 688
rect 105740 480 105768 682
rect 106936 480 106964 1294
rect 107304 746 107332 3726
rect 108408 1358 108436 3726
rect 108396 1352 108448 1358
rect 108396 1294 108448 1300
rect 109316 1352 109368 1358
rect 109316 1294 109368 1300
rect 108120 1284 108172 1290
rect 108120 1226 108172 1232
rect 107292 740 107344 746
rect 107292 682 107344 688
rect 108132 480 108160 1226
rect 109328 480 109356 1294
rect 109604 1290 109632 3726
rect 110708 1358 110736 3726
rect 110696 1352 110748 1358
rect 110696 1294 110748 1300
rect 111904 1290 111932 3726
rect 112812 1352 112864 1358
rect 112812 1294 112864 1300
rect 109592 1284 109644 1290
rect 109592 1226 109644 1232
rect 110512 1284 110564 1290
rect 110512 1226 110564 1232
rect 111892 1284 111944 1290
rect 111892 1226 111944 1232
rect 110524 480 110552 1226
rect 111616 1148 111668 1154
rect 111616 1090 111668 1096
rect 111628 480 111656 1090
rect 112824 480 112852 1294
rect 113100 1154 113128 3726
rect 114204 1358 114232 3726
rect 114192 1352 114244 1358
rect 114192 1294 114244 1300
rect 115204 1284 115256 1290
rect 115204 1226 115256 1232
rect 114008 1216 114060 1222
rect 114008 1158 114060 1164
rect 113088 1148 113140 1154
rect 113088 1090 113140 1096
rect 114020 480 114048 1158
rect 115216 480 115244 1226
rect 115400 1222 115428 3726
rect 116400 1352 116452 1358
rect 116400 1294 116452 1300
rect 115388 1216 115440 1222
rect 115388 1158 115440 1164
rect 116412 480 116440 1294
rect 116596 1290 116624 3726
rect 117700 1358 117728 3726
rect 117688 1352 117740 1358
rect 117688 1294 117740 1300
rect 118896 1290 118924 3726
rect 116584 1284 116636 1290
rect 116584 1226 116636 1232
rect 117596 1284 117648 1290
rect 117596 1226 117648 1232
rect 118884 1284 118936 1290
rect 118884 1226 118936 1232
rect 117608 480 117636 1226
rect 66690 190 67128 218
rect 66690 -960 66802 190
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 354 118874 480
rect 119264 354 119292 3726
rect 121196 1358 121224 3726
rect 119896 1352 119948 1358
rect 119896 1294 119948 1300
rect 121184 1352 121236 1358
rect 121184 1294 121236 1300
rect 119908 480 119936 1294
rect 122288 1284 122340 1290
rect 122288 1226 122340 1232
rect 121092 944 121144 950
rect 121092 886 121144 892
rect 121104 480 121132 886
rect 122300 480 122328 1226
rect 122392 950 122420 3726
rect 123496 1290 123524 3726
rect 123484 1284 123536 1290
rect 123484 1226 123536 1232
rect 124680 1284 124732 1290
rect 124680 1226 124732 1232
rect 123484 1148 123536 1154
rect 123484 1090 123536 1096
rect 122380 944 122432 950
rect 122380 886 122432 892
rect 123496 480 123524 1090
rect 124692 480 124720 1226
rect 124784 1154 124812 3726
rect 125796 3726 125868 3754
rect 126992 3726 127064 3754
rect 127176 3726 128260 3754
rect 129292 3726 129364 3754
rect 130488 3726 130560 3754
rect 131592 3726 131664 3754
rect 132788 3726 132860 3754
rect 133984 3726 134056 3754
rect 134168 3726 135160 3754
rect 135272 3726 136356 3754
rect 137388 3726 137460 3754
rect 138584 3726 138656 3754
rect 139780 3726 139852 3754
rect 140884 3726 140956 3754
rect 141712 3726 142152 3754
rect 142448 3726 143348 3754
rect 143552 3726 144452 3754
rect 145576 3726 145648 3754
rect 146680 3726 146752 3754
rect 147600 3726 147948 3754
rect 149072 3726 149144 3754
rect 149992 3726 150248 3754
rect 151096 3726 151444 3754
rect 151832 3726 152548 3754
rect 153488 3726 153744 3754
rect 154868 3726 154940 3754
rect 155880 3726 156044 3754
rect 156616 3726 157240 3754
rect 158272 3726 158344 3754
rect 159376 3726 159540 3754
rect 160112 3726 160736 3754
rect 161584 3726 161840 3754
rect 162964 3726 163036 3754
rect 164068 3726 164140 3754
rect 164896 3726 165336 3754
rect 166460 3726 166532 3754
rect 167564 3726 167636 3754
rect 168392 3726 168832 3754
rect 169956 3726 170028 3754
rect 170784 3726 171132 3754
rect 172256 3726 172328 3754
rect 173176 3726 173432 3754
rect 174280 3726 174628 3754
rect 175752 3726 175824 3754
rect 176672 3726 176928 3754
rect 178052 3726 178124 3754
rect 179064 3726 179228 3754
rect 180396 3754 180424 4012
rect 181592 3754 181620 4012
rect 182696 3754 182724 4012
rect 180396 3726 180472 3754
rect 125796 1290 125824 3726
rect 126992 1358 127020 3726
rect 125876 1352 125928 1358
rect 125876 1294 125928 1300
rect 126980 1352 127032 1358
rect 126980 1294 127032 1300
rect 125784 1284 125836 1290
rect 125784 1226 125836 1232
rect 124772 1148 124824 1154
rect 124772 1090 124824 1096
rect 125888 480 125916 1294
rect 127176 1170 127204 3726
rect 129292 1290 129320 3726
rect 130488 1358 130516 3726
rect 131592 1358 131620 3726
rect 132788 1358 132816 3726
rect 133984 1358 134012 3726
rect 129372 1352 129424 1358
rect 129372 1294 129424 1300
rect 130476 1352 130528 1358
rect 130476 1294 130528 1300
rect 130568 1352 130620 1358
rect 130568 1294 130620 1300
rect 131580 1352 131632 1358
rect 131580 1294 131632 1300
rect 131764 1352 131816 1358
rect 131764 1294 131816 1300
rect 132776 1352 132828 1358
rect 132776 1294 132828 1300
rect 132960 1352 133012 1358
rect 132960 1294 133012 1300
rect 133972 1352 134024 1358
rect 133972 1294 134024 1300
rect 128176 1284 128228 1290
rect 128176 1226 128228 1232
rect 129280 1284 129332 1290
rect 129280 1226 129332 1232
rect 126992 1142 127204 1170
rect 126992 480 127020 1142
rect 128188 480 128216 1226
rect 129384 480 129412 1294
rect 130580 480 130608 1294
rect 131776 480 131804 1294
rect 132972 480 133000 1294
rect 134168 480 134196 3726
rect 135272 480 135300 3726
rect 137388 1290 137416 3726
rect 138584 1358 138612 3726
rect 137652 1352 137704 1358
rect 137652 1294 137704 1300
rect 138572 1352 138624 1358
rect 138572 1294 138624 1300
rect 136456 1284 136508 1290
rect 136456 1226 136508 1232
rect 137376 1284 137428 1290
rect 137376 1226 137428 1232
rect 136468 480 136496 1226
rect 137664 480 137692 1294
rect 139780 1290 139808 3726
rect 140884 1290 140912 3726
rect 138848 1284 138900 1290
rect 138848 1226 138900 1232
rect 139768 1284 139820 1290
rect 139768 1226 139820 1232
rect 140044 1284 140096 1290
rect 140044 1226 140096 1232
rect 140872 1284 140924 1290
rect 140872 1226 140924 1232
rect 138860 480 138888 1226
rect 140056 480 140084 1226
rect 118762 326 119292 354
rect 118762 -960 118874 326
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 354 141322 480
rect 141712 354 141740 3726
rect 142448 480 142476 3726
rect 143552 480 143580 3726
rect 145576 1358 145604 3726
rect 146680 1358 146708 3726
rect 144736 1352 144788 1358
rect 144736 1294 144788 1300
rect 145564 1352 145616 1358
rect 145564 1294 145616 1300
rect 145932 1352 145984 1358
rect 145932 1294 145984 1300
rect 146668 1352 146720 1358
rect 146668 1294 146720 1300
rect 144748 480 144776 1294
rect 145944 480 145972 1294
rect 141210 326 141740 354
rect 141210 -960 141322 326
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 354 147210 480
rect 147600 354 147628 3726
rect 149072 1358 149100 3726
rect 148324 1352 148376 1358
rect 148324 1294 148376 1300
rect 149060 1352 149112 1358
rect 149060 1294 149112 1300
rect 148336 480 148364 1294
rect 147098 326 147628 354
rect 147098 -960 147210 326
rect 148294 -960 148406 480
rect 149490 354 149602 480
rect 149992 354 150020 3726
rect 149490 326 150020 354
rect 150594 354 150706 480
rect 151096 354 151124 3726
rect 151832 480 151860 3726
rect 150594 326 151124 354
rect 149490 -960 149602 326
rect 150594 -960 150706 326
rect 151790 -960 151902 480
rect 152986 354 153098 480
rect 153488 354 153516 3726
rect 154868 1358 154896 3726
rect 154212 1352 154264 1358
rect 154212 1294 154264 1300
rect 154856 1352 154908 1358
rect 154856 1294 154908 1300
rect 154224 480 154252 1294
rect 152986 326 153516 354
rect 152986 -960 153098 326
rect 154182 -960 154294 480
rect 155378 354 155490 480
rect 155880 354 155908 3726
rect 156616 480 156644 3726
rect 155378 326 155908 354
rect 155378 -960 155490 326
rect 156574 -960 156686 480
rect 157770 354 157882 480
rect 158272 354 158300 3726
rect 157770 326 158300 354
rect 158874 354 158986 480
rect 159376 354 159404 3726
rect 160112 480 160140 3726
rect 158874 326 159404 354
rect 157770 -960 157882 326
rect 158874 -960 158986 326
rect 160070 -960 160182 480
rect 161266 354 161378 480
rect 161584 354 161612 3726
rect 162964 1358 162992 3726
rect 162492 1352 162544 1358
rect 162492 1294 162544 1300
rect 162952 1352 163004 1358
rect 162952 1294 163004 1300
rect 162504 480 162532 1294
rect 161266 326 161612 354
rect 161266 -960 161378 326
rect 162462 -960 162574 480
rect 163658 354 163770 480
rect 164068 354 164096 3726
rect 164896 480 164924 3726
rect 163658 326 164096 354
rect 163658 -960 163770 326
rect 164854 -960 164966 480
rect 166050 354 166162 480
rect 166460 354 166488 3726
rect 166050 326 166488 354
rect 167154 354 167266 480
rect 167564 354 167592 3726
rect 168392 480 168420 3726
rect 167154 326 167592 354
rect 166050 -960 166162 326
rect 167154 -960 167266 326
rect 168350 -960 168462 480
rect 169546 354 169658 480
rect 169956 354 169984 3726
rect 170784 480 170812 3726
rect 169546 326 169984 354
rect 169546 -960 169658 326
rect 170742 -960 170854 480
rect 171938 354 172050 480
rect 172256 354 172284 3726
rect 173176 480 173204 3726
rect 174280 480 174308 3726
rect 171938 326 172284 354
rect 171938 -960 172050 326
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 354 175546 480
rect 175752 354 175780 3726
rect 176672 480 176700 3726
rect 175434 326 175780 354
rect 175434 -960 175546 326
rect 176630 -960 176742 480
rect 177826 354 177938 480
rect 178052 354 178080 3726
rect 179064 480 179092 3726
rect 177826 326 178080 354
rect 177826 -960 177938 326
rect 179022 -960 179134 480
rect 180218 218 180330 480
rect 180444 218 180472 3726
rect 181456 3726 181620 3754
rect 182560 3726 182724 3754
rect 183892 3754 183920 4012
rect 184996 3754 185024 4012
rect 186192 3754 186220 4012
rect 187388 3754 187416 4012
rect 183892 3726 183968 3754
rect 181456 480 181484 3726
rect 182560 480 182588 3726
rect 180218 190 180472 218
rect 180218 -960 180330 190
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 218 183826 480
rect 183940 218 183968 3726
rect 184952 3726 185024 3754
rect 186148 3726 186220 3754
rect 187344 3726 187416 3754
rect 188492 3754 188520 4012
rect 189688 3754 189716 4012
rect 190792 3754 190820 4012
rect 191988 3754 192016 4012
rect 193184 3754 193212 4012
rect 194288 3754 194316 4012
rect 195484 3754 195512 4012
rect 188492 3726 188568 3754
rect 189688 3726 189764 3754
rect 190792 3726 190868 3754
rect 191988 3726 192064 3754
rect 193184 3726 193260 3754
rect 194288 3726 194456 3754
rect 184952 480 184980 3726
rect 186148 480 186176 3726
rect 187344 480 187372 3726
rect 188540 480 188568 3726
rect 189736 480 189764 3726
rect 190840 480 190868 3726
rect 192036 480 192064 3726
rect 193232 480 193260 3726
rect 194428 480 194456 3726
rect 195440 3726 195512 3754
rect 196680 3754 196708 4012
rect 197784 3754 197812 4012
rect 198980 3754 199008 4012
rect 196680 3726 196848 3754
rect 197784 3726 197952 3754
rect 183714 190 183968 218
rect 183714 -960 183826 190
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195440 218 195468 3726
rect 196820 480 196848 3726
rect 197924 480 197952 3726
rect 198936 3726 199008 3754
rect 200084 3754 200112 4012
rect 201280 3754 201308 4012
rect 202476 3754 202504 4012
rect 203580 3754 203608 4012
rect 204776 3754 204804 4012
rect 205880 3754 205908 4012
rect 207076 3754 207104 4012
rect 208272 3754 208300 4012
rect 209376 3754 209404 4012
rect 210572 3754 210600 4012
rect 211676 3754 211704 4012
rect 212872 3754 212900 4012
rect 214068 3754 214096 4012
rect 215172 3754 215200 4012
rect 216368 3806 216396 4012
rect 216356 3800 216408 3806
rect 200084 3726 200344 3754
rect 201280 3726 201356 3754
rect 202476 3726 202736 3754
rect 203580 3726 203656 3754
rect 204776 3726 205128 3754
rect 205880 3726 206232 3754
rect 207076 3726 207152 3754
rect 208272 3726 208624 3754
rect 209376 3726 209728 3754
rect 210572 3726 211016 3754
rect 211676 3726 211752 3754
rect 212872 3726 213408 3754
rect 214068 3726 214512 3754
rect 215172 3726 215248 3754
rect 216356 3742 216408 3748
rect 216864 3800 216916 3806
rect 216864 3742 216916 3748
rect 217472 3754 217500 4012
rect 218668 3754 218696 4012
rect 219864 3754 219892 4012
rect 220968 3754 220996 4012
rect 222164 3806 222192 4012
rect 222152 3800 222204 3806
rect 195582 218 195694 480
rect 195440 190 195694 218
rect 195582 -960 195694 190
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198936 218 198964 3726
rect 200316 480 200344 3726
rect 199078 218 199190 480
rect 198936 190 199190 218
rect 199078 -960 199190 190
rect 200274 -960 200386 480
rect 201328 354 201356 3726
rect 202708 480 202736 3726
rect 201470 354 201582 480
rect 201328 326 201582 354
rect 201470 -960 201582 326
rect 202666 -960 202778 480
rect 203628 354 203656 3726
rect 205100 480 205128 3726
rect 206204 480 206232 3726
rect 203862 354 203974 480
rect 203628 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207124 354 207152 3726
rect 208596 480 208624 3726
rect 209700 626 209728 3726
rect 209700 598 209774 626
rect 209746 480 209774 598
rect 210988 480 211016 3726
rect 207358 354 207470 480
rect 207124 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209746 326 209862 480
rect 209750 -960 209862 326
rect 210946 -960 211058 480
rect 211724 354 211752 3726
rect 213380 480 213408 3726
rect 214484 480 214512 3726
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215220 354 215248 3726
rect 216876 480 216904 3742
rect 217472 3726 217640 3754
rect 218668 3726 219296 3754
rect 219864 3726 220032 3754
rect 220968 3726 221136 3754
rect 222152 3742 222204 3748
rect 222752 3800 222804 3806
rect 222752 3742 222804 3748
rect 223360 3754 223388 4012
rect 224464 3806 224492 4012
rect 224452 3800 224504 3806
rect 215638 354 215750 480
rect 215220 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 217612 354 217640 3726
rect 219268 480 219296 3726
rect 218030 354 218142 480
rect 217612 326 218142 354
rect 218030 -960 218142 326
rect 219226 -960 219338 480
rect 220004 354 220032 3726
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 3726
rect 222764 480 222792 3742
rect 223360 3726 223528 3754
rect 224452 3742 224504 3748
rect 225144 3800 225196 3806
rect 225144 3742 225196 3748
rect 225660 3754 225688 4012
rect 226764 3754 226792 4012
rect 227960 3754 227988 4012
rect 229156 3754 229184 4012
rect 230260 3806 230288 4012
rect 231456 3806 231484 4012
rect 232560 3806 232588 4012
rect 233756 3806 233784 4012
rect 230248 3800 230300 3806
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223500 354 223528 3726
rect 225156 480 225184 3742
rect 225660 3726 225920 3754
rect 226764 3726 227576 3754
rect 227960 3726 228312 3754
rect 229156 3726 229416 3754
rect 230248 3742 230300 3748
rect 231032 3800 231084 3806
rect 231032 3742 231084 3748
rect 231444 3800 231496 3806
rect 231444 3742 231496 3748
rect 232228 3800 232280 3806
rect 232228 3742 232280 3748
rect 232548 3800 232600 3806
rect 232548 3742 232600 3748
rect 233424 3800 233476 3806
rect 233424 3742 233476 3748
rect 233744 3800 233796 3806
rect 233744 3742 233796 3748
rect 234620 3800 234672 3806
rect 234620 3742 234672 3748
rect 234952 3754 234980 4012
rect 236056 3754 236084 4012
rect 237252 3806 237280 4012
rect 238356 3806 238384 4012
rect 239552 3806 239580 4012
rect 240748 3806 240776 4012
rect 241852 3806 241880 4012
rect 237240 3800 237292 3806
rect 223918 354 224030 480
rect 223500 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 225892 354 225920 3726
rect 227548 480 227576 3726
rect 226310 354 226422 480
rect 225892 326 226422 354
rect 226310 -960 226422 326
rect 227506 -960 227618 480
rect 228284 354 228312 3726
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 3726
rect 231044 480 231072 3742
rect 232240 480 232268 3742
rect 233436 480 233464 3742
rect 234632 480 234660 3742
rect 234952 3726 235856 3754
rect 236056 3726 236592 3754
rect 237240 3742 237292 3748
rect 238116 3800 238168 3806
rect 238116 3742 238168 3748
rect 238344 3800 238396 3806
rect 238344 3742 238396 3748
rect 239312 3800 239364 3806
rect 239312 3742 239364 3748
rect 239540 3800 239592 3806
rect 239540 3742 239592 3748
rect 240508 3800 240560 3806
rect 240508 3742 240560 3748
rect 240736 3800 240788 3806
rect 240736 3742 240788 3748
rect 241704 3800 241756 3806
rect 241704 3742 241756 3748
rect 241840 3800 241892 3806
rect 241840 3742 241892 3748
rect 242900 3800 242952 3806
rect 242900 3742 242952 3748
rect 243048 3754 243076 4012
rect 244152 3874 244180 4012
rect 244140 3868 244192 3874
rect 244140 3810 244192 3816
rect 245200 3868 245252 3874
rect 245200 3810 245252 3816
rect 235828 480 235856 3726
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 3726
rect 238128 480 238156 3742
rect 239324 480 239352 3742
rect 240520 480 240548 3742
rect 241716 480 241744 3742
rect 242912 480 242940 3742
rect 243048 3726 244136 3754
rect 244108 480 244136 3726
rect 245212 480 245240 3810
rect 245348 3806 245376 4012
rect 246544 3806 246572 4012
rect 247648 3942 247676 4012
rect 247636 3936 247688 3942
rect 247636 3878 247688 3884
rect 248604 3936 248656 3942
rect 248604 3878 248656 3884
rect 248844 3890 248872 4012
rect 245336 3800 245388 3806
rect 245336 3742 245388 3748
rect 246396 3800 246448 3806
rect 246396 3742 246448 3748
rect 246532 3800 246584 3806
rect 246532 3742 246584 3748
rect 247592 3800 247644 3806
rect 247592 3742 247644 3748
rect 246408 480 246436 3742
rect 247604 480 247632 3742
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 236982 -960 237094 326
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248616 354 248644 3878
rect 248844 3862 248920 3890
rect 248892 2854 248920 3862
rect 250040 3806 250068 4012
rect 251144 3890 251172 4012
rect 251100 3862 251172 3890
rect 250028 3800 250080 3806
rect 250028 3742 250080 3748
rect 251100 2854 251128 3862
rect 252340 3806 252368 4012
rect 253444 3890 253472 4012
rect 254640 3890 254668 4012
rect 253400 3862 253472 3890
rect 254596 3862 254668 3890
rect 251180 3800 251232 3806
rect 251180 3742 251232 3748
rect 252328 3800 252380 3806
rect 252328 3742 252380 3748
rect 248880 2848 248932 2854
rect 248880 2790 248932 2796
rect 249984 2848 250036 2854
rect 249984 2790 250036 2796
rect 251088 2848 251140 2854
rect 251088 2790 251140 2796
rect 249996 480 250024 2790
rect 251192 480 251220 3742
rect 253400 2922 253428 3862
rect 253480 3800 253532 3806
rect 253480 3742 253532 3748
rect 253388 2916 253440 2922
rect 253388 2858 253440 2864
rect 252376 2848 252428 2854
rect 252376 2790 252428 2796
rect 252388 480 252416 2790
rect 253492 480 253520 3742
rect 254596 2854 254624 3862
rect 255836 3806 255864 4012
rect 256940 3874 256968 4012
rect 256928 3868 256980 3874
rect 256928 3810 256980 3816
rect 258136 3806 258164 4012
rect 259240 3874 259268 4012
rect 258264 3868 258316 3874
rect 258264 3810 258316 3816
rect 259228 3868 259280 3874
rect 259228 3810 259280 3816
rect 255824 3800 255876 3806
rect 255824 3742 255876 3748
rect 257068 3800 257120 3806
rect 257068 3742 257120 3748
rect 258124 3800 258176 3806
rect 258124 3742 258176 3748
rect 254676 2916 254728 2922
rect 254676 2858 254728 2864
rect 254584 2848 254636 2854
rect 254584 2790 254636 2796
rect 254688 480 254716 2858
rect 255872 2848 255924 2854
rect 255872 2790 255924 2796
rect 255884 480 255912 2790
rect 257080 480 257108 3742
rect 258276 480 258304 3810
rect 260436 3806 260464 4012
rect 261632 3874 261660 4012
rect 260656 3868 260708 3874
rect 260656 3810 260708 3816
rect 261620 3868 261672 3874
rect 261620 3810 261672 3816
rect 259460 3800 259512 3806
rect 259460 3742 259512 3748
rect 260424 3800 260476 3806
rect 260424 3742 260476 3748
rect 259472 480 259500 3742
rect 260668 480 260696 3810
rect 262736 3806 262764 4012
rect 263932 3874 263960 4012
rect 262956 3868 263008 3874
rect 262956 3810 263008 3816
rect 263920 3868 263972 3874
rect 263920 3810 263972 3816
rect 261760 3800 261812 3806
rect 261760 3742 261812 3748
rect 262724 3800 262776 3806
rect 262724 3742 262776 3748
rect 261772 480 261800 3742
rect 262968 480 262996 3810
rect 265036 3806 265064 4012
rect 265348 3868 265400 3874
rect 265348 3810 265400 3816
rect 264152 3800 264204 3806
rect 264152 3742 264204 3748
rect 265024 3800 265076 3806
rect 265024 3742 265076 3748
rect 264164 480 264192 3742
rect 265360 480 265388 3810
rect 266232 3754 266260 4012
rect 267428 3806 267456 4012
rect 268532 3874 268560 4012
rect 268520 3868 268572 3874
rect 268520 3810 268572 3816
rect 269728 3806 269756 4012
rect 270832 3874 270860 4012
rect 270040 3868 270092 3874
rect 270040 3810 270092 3816
rect 270820 3868 270872 3874
rect 270820 3810 270872 3816
rect 266544 3800 266596 3806
rect 266232 3726 266308 3754
rect 266544 3742 266596 3748
rect 267416 3800 267468 3806
rect 267416 3742 267468 3748
rect 268844 3800 268896 3806
rect 268844 3742 268896 3748
rect 269716 3800 269768 3806
rect 269716 3742 269768 3748
rect 266280 1358 266308 3726
rect 266268 1352 266320 1358
rect 266268 1294 266320 1300
rect 266556 480 266584 3742
rect 267740 1352 267792 1358
rect 267740 1294 267792 1300
rect 267752 480 267780 1294
rect 268856 480 268884 3742
rect 270052 480 270080 3810
rect 272028 3806 272056 4012
rect 272432 3868 272484 3874
rect 272432 3810 272484 3816
rect 271236 3800 271288 3806
rect 271236 3742 271288 3748
rect 272016 3800 272068 3806
rect 272016 3742 272068 3748
rect 271248 480 271276 3742
rect 272444 480 272472 3810
rect 273224 3754 273252 4012
rect 273180 3726 273252 3754
rect 273628 3800 273680 3806
rect 273628 3742 273680 3748
rect 274328 3754 274356 4012
rect 275524 3874 275552 4012
rect 275512 3868 275564 3874
rect 275512 3810 275564 3816
rect 276720 3806 276748 4012
rect 277824 3874 277852 4012
rect 277124 3868 277176 3874
rect 277124 3810 277176 3816
rect 277812 3868 277864 3874
rect 277812 3810 277864 3816
rect 276708 3800 276760 3806
rect 273180 1358 273208 3726
rect 273168 1352 273220 1358
rect 273168 1294 273220 1300
rect 273640 480 273668 3742
rect 274328 3726 274404 3754
rect 276708 3742 276760 3748
rect 274376 746 274404 3726
rect 274824 1352 274876 1358
rect 274824 1294 274876 1300
rect 274364 740 274416 746
rect 274364 682 274416 688
rect 274836 480 274864 1294
rect 276020 740 276072 746
rect 276020 682 276072 688
rect 276032 480 276060 682
rect 277136 480 277164 3810
rect 279020 3806 279048 4012
rect 279516 3868 279568 3874
rect 279516 3810 279568 3816
rect 278320 3800 278372 3806
rect 278320 3742 278372 3748
rect 279008 3800 279060 3806
rect 279008 3742 279060 3748
rect 278332 480 278360 3742
rect 279528 480 279556 3810
rect 280124 3754 280152 4012
rect 280080 3726 280152 3754
rect 280712 3800 280764 3806
rect 280712 3742 280764 3748
rect 281320 3754 281348 4012
rect 282516 3754 282544 4012
rect 283620 3806 283648 4012
rect 284816 3874 284844 4012
rect 285920 3942 285948 4012
rect 285908 3936 285960 3942
rect 285908 3878 285960 3884
rect 284804 3868 284856 3874
rect 284804 3810 284856 3816
rect 286600 3868 286652 3874
rect 286600 3810 286652 3816
rect 283608 3800 283660 3806
rect 280080 1358 280108 3726
rect 280068 1352 280120 1358
rect 280068 1294 280120 1300
rect 280724 480 280752 3742
rect 281320 3726 281396 3754
rect 282516 3726 282592 3754
rect 283608 3742 283660 3748
rect 285404 3800 285456 3806
rect 285404 3742 285456 3748
rect 281368 1290 281396 3726
rect 282564 1358 282592 3726
rect 281908 1352 281960 1358
rect 281908 1294 281960 1300
rect 282552 1352 282604 1358
rect 282552 1294 282604 1300
rect 284300 1352 284352 1358
rect 284300 1294 284352 1300
rect 281356 1284 281408 1290
rect 281356 1226 281408 1232
rect 281920 480 281948 1294
rect 283104 1284 283156 1290
rect 283104 1226 283156 1232
rect 283116 480 283144 1226
rect 284312 480 284340 1294
rect 285416 480 285444 3742
rect 286612 480 286640 3810
rect 287116 3806 287144 4012
rect 287796 3936 287848 3942
rect 287796 3878 287848 3884
rect 287104 3800 287156 3806
rect 287104 3742 287156 3748
rect 287808 480 287836 3878
rect 288312 3754 288340 4012
rect 288992 3800 289044 3806
rect 288312 3726 288388 3754
rect 288992 3742 289044 3748
rect 289416 3754 289444 4012
rect 290612 3754 290640 4012
rect 291716 3806 291744 4012
rect 292912 3874 292940 4012
rect 292900 3868 292952 3874
rect 292900 3810 292952 3816
rect 294108 3806 294136 4012
rect 294880 3868 294932 3874
rect 294880 3810 294932 3816
rect 291704 3800 291756 3806
rect 288360 1358 288388 3726
rect 288348 1352 288400 1358
rect 288348 1294 288400 1300
rect 289004 480 289032 3742
rect 289416 3726 289492 3754
rect 290612 3726 290688 3754
rect 291704 3742 291756 3748
rect 293684 3800 293736 3806
rect 293684 3742 293736 3748
rect 294096 3800 294148 3806
rect 294096 3742 294148 3748
rect 289464 1290 289492 3726
rect 290188 1352 290240 1358
rect 290188 1294 290240 1300
rect 289452 1284 289504 1290
rect 289452 1226 289504 1232
rect 290200 480 290228 1294
rect 290660 610 290688 3726
rect 291384 1284 291436 1290
rect 291384 1226 291436 1232
rect 290648 604 290700 610
rect 290648 546 290700 552
rect 291396 480 291424 1226
rect 292580 604 292632 610
rect 292580 546 292632 552
rect 292592 480 292620 546
rect 293696 480 293724 3742
rect 294892 480 294920 3810
rect 295212 3754 295240 4012
rect 296076 3800 296128 3806
rect 295212 3726 295288 3754
rect 296076 3742 296128 3748
rect 296408 3754 296436 4012
rect 297512 3754 297540 4012
rect 298708 3806 298736 4012
rect 299904 3874 299932 4012
rect 299892 3868 299944 3874
rect 299892 3810 299944 3816
rect 301008 3806 301036 4012
rect 301964 3868 302016 3874
rect 301964 3810 302016 3816
rect 298696 3800 298748 3806
rect 295260 1358 295288 3726
rect 295248 1352 295300 1358
rect 295248 1294 295300 1300
rect 296088 480 296116 3742
rect 296408 3726 296484 3754
rect 297512 3726 297588 3754
rect 298696 3742 298748 3748
rect 300768 3800 300820 3806
rect 300768 3742 300820 3748
rect 300996 3800 301048 3806
rect 300996 3742 301048 3748
rect 296456 1290 296484 3726
rect 297560 1358 297588 3726
rect 297272 1352 297324 1358
rect 297272 1294 297324 1300
rect 297548 1352 297600 1358
rect 297548 1294 297600 1300
rect 299664 1352 299716 1358
rect 299664 1294 299716 1300
rect 296444 1284 296496 1290
rect 296444 1226 296496 1232
rect 297284 480 297312 1294
rect 298468 1284 298520 1290
rect 298468 1226 298520 1232
rect 298480 480 298508 1226
rect 299676 480 299704 1294
rect 300780 480 300808 3742
rect 301976 480 302004 3810
rect 302204 3754 302232 4012
rect 302160 3726 302232 3754
rect 303160 3800 303212 3806
rect 303160 3742 303212 3748
rect 303308 3754 303336 4012
rect 304504 3754 304532 4012
rect 305700 3754 305728 4012
rect 306804 3874 306832 4012
rect 306792 3868 306844 3874
rect 306792 3810 306844 3816
rect 308000 3806 308028 4012
rect 309048 3868 309100 3874
rect 309048 3810 309100 3816
rect 307988 3800 308040 3806
rect 302160 1358 302188 3726
rect 302148 1352 302200 1358
rect 302148 1294 302200 1300
rect 303172 480 303200 3742
rect 303308 3726 303384 3754
rect 304504 3726 304580 3754
rect 305700 3726 305776 3754
rect 307988 3742 308040 3748
rect 303356 1290 303384 3726
rect 304356 1352 304408 1358
rect 304356 1294 304408 1300
rect 303344 1284 303396 1290
rect 303344 1226 303396 1232
rect 304368 480 304396 1294
rect 304552 610 304580 3726
rect 305748 1358 305776 3726
rect 305736 1352 305788 1358
rect 305736 1294 305788 1300
rect 307944 1352 307996 1358
rect 307944 1294 307996 1300
rect 305552 1284 305604 1290
rect 305552 1226 305604 1232
rect 304540 604 304592 610
rect 304540 546 304592 552
rect 305564 480 305592 1226
rect 306748 604 306800 610
rect 306748 546 306800 552
rect 306760 480 306788 546
rect 307956 480 307984 1294
rect 309060 480 309088 3810
rect 309196 3754 309224 4012
rect 310300 3890 310328 4012
rect 311496 3890 311524 4012
rect 310300 3862 310376 3890
rect 311496 3862 311572 3890
rect 310244 3800 310296 3806
rect 309196 3726 309272 3754
rect 310244 3742 310296 3748
rect 309244 2854 309272 3726
rect 309232 2848 309284 2854
rect 309232 2790 309284 2796
rect 310256 480 310284 3742
rect 310348 1358 310376 3862
rect 311440 2848 311492 2854
rect 311440 2790 311492 2796
rect 310336 1352 310388 1358
rect 310336 1294 310388 1300
rect 311452 480 311480 2790
rect 311544 1222 311572 3862
rect 312600 3754 312628 4012
rect 312556 3726 312628 3754
rect 313796 3754 313824 4012
rect 314992 3754 315020 4012
rect 316096 3806 316124 4012
rect 316084 3800 316136 3806
rect 313796 3726 313872 3754
rect 314992 3726 315068 3754
rect 317292 3754 317320 4012
rect 316084 3742 316136 3748
rect 312556 1290 312584 3726
rect 313844 1358 313872 3726
rect 315040 2854 315068 3726
rect 317248 3726 317320 3754
rect 318396 3754 318424 4012
rect 318524 3800 318576 3806
rect 318396 3726 318472 3754
rect 318524 3742 318576 3748
rect 319592 3754 319620 4012
rect 320788 3754 320816 4012
rect 321892 3754 321920 4012
rect 323088 3806 323116 4012
rect 323076 3800 323128 3806
rect 315028 2848 315080 2854
rect 315028 2790 315080 2796
rect 317248 1358 317276 3726
rect 317328 2848 317380 2854
rect 317328 2790 317380 2796
rect 312636 1352 312688 1358
rect 312636 1294 312688 1300
rect 313832 1352 313884 1358
rect 313832 1294 313884 1300
rect 316224 1352 316276 1358
rect 316224 1294 316276 1300
rect 317236 1352 317288 1358
rect 317236 1294 317288 1300
rect 312544 1284 312596 1290
rect 312544 1226 312596 1232
rect 311532 1216 311584 1222
rect 311532 1158 311584 1164
rect 312648 480 312676 1294
rect 315028 1284 315080 1290
rect 315028 1226 315080 1232
rect 313832 1216 313884 1222
rect 313832 1158 313884 1164
rect 313844 480 313872 1158
rect 315040 480 315068 1226
rect 316236 480 316264 1294
rect 317340 480 317368 2790
rect 318444 1290 318472 3726
rect 318432 1284 318484 1290
rect 318432 1226 318484 1232
rect 318536 480 318564 3742
rect 319592 3726 319668 3754
rect 320788 3726 320864 3754
rect 321892 3726 321968 3754
rect 323076 3742 323128 3748
rect 324192 3754 324220 4012
rect 325388 3754 325416 4012
rect 325608 3800 325660 3806
rect 324192 3726 324268 3754
rect 325388 3726 325464 3754
rect 325608 3742 325660 3748
rect 326584 3754 326612 4012
rect 327688 3754 327716 4012
rect 328884 3754 328912 4012
rect 329988 3754 330016 4012
rect 331184 3754 331212 4012
rect 319640 1222 319668 3726
rect 319720 1352 319772 1358
rect 319720 1294 319772 1300
rect 319628 1216 319680 1222
rect 319628 1158 319680 1164
rect 319732 480 319760 1294
rect 320836 1154 320864 3726
rect 321940 1358 321968 3726
rect 321928 1352 321980 1358
rect 321928 1294 321980 1300
rect 320916 1284 320968 1290
rect 320916 1226 320968 1232
rect 320824 1148 320876 1154
rect 320824 1090 320876 1096
rect 320928 480 320956 1226
rect 322112 1216 322164 1222
rect 322112 1158 322164 1164
rect 322124 480 322152 1158
rect 323308 1148 323360 1154
rect 323308 1090 323360 1096
rect 323320 480 323348 1090
rect 324240 610 324268 3726
rect 324412 1352 324464 1358
rect 324412 1294 324464 1300
rect 324228 604 324280 610
rect 324228 546 324280 552
rect 324424 480 324452 1294
rect 325436 1018 325464 3726
rect 325424 1012 325476 1018
rect 325424 954 325476 960
rect 325620 480 325648 3742
rect 326584 3726 326660 3754
rect 327688 3726 327764 3754
rect 328884 3726 328960 3754
rect 329988 3726 330064 3754
rect 326632 1358 326660 3726
rect 326620 1352 326672 1358
rect 326620 1294 326672 1300
rect 327736 610 327764 3726
rect 328932 1290 328960 3726
rect 329196 1352 329248 1358
rect 329196 1294 329248 1300
rect 328920 1284 328972 1290
rect 328920 1226 328972 1232
rect 328000 1012 328052 1018
rect 328000 954 328052 960
rect 326804 604 326856 610
rect 326804 546 326856 552
rect 327724 604 327776 610
rect 327724 546 327776 552
rect 326816 480 326844 546
rect 328012 480 328040 954
rect 329208 480 329236 1294
rect 330036 1222 330064 3726
rect 331140 3726 331212 3754
rect 332380 3754 332408 4012
rect 333484 3754 333512 4012
rect 334680 3754 334708 4012
rect 335876 3754 335904 4012
rect 336980 3754 337008 4012
rect 338176 3754 338204 4012
rect 339280 3754 339308 4012
rect 340476 3754 340504 4012
rect 341672 3754 341700 4012
rect 342776 3754 342804 4012
rect 343972 3754 344000 4012
rect 345076 3754 345104 4012
rect 346272 3754 346300 4012
rect 347468 3754 347496 4012
rect 348572 3754 348600 4012
rect 349768 3754 349796 4012
rect 350872 3754 350900 4012
rect 352068 3754 352096 4012
rect 353264 3754 353292 4012
rect 332380 3726 332456 3754
rect 333484 3726 333560 3754
rect 334680 3726 334756 3754
rect 335876 3726 335952 3754
rect 336980 3726 337056 3754
rect 338176 3726 338252 3754
rect 339280 3726 339356 3754
rect 340476 3726 340552 3754
rect 341672 3726 341748 3754
rect 342776 3726 342852 3754
rect 343972 3726 344048 3754
rect 345076 3726 345152 3754
rect 346272 3726 346348 3754
rect 347468 3726 347544 3754
rect 348572 3726 348648 3754
rect 349768 3726 349844 3754
rect 350872 3726 350948 3754
rect 352068 3726 352144 3754
rect 330024 1216 330076 1222
rect 330024 1158 330076 1164
rect 331140 1154 331168 3726
rect 332428 1358 332456 3726
rect 332416 1352 332468 1358
rect 332416 1294 332468 1300
rect 331588 1284 331640 1290
rect 331588 1226 331640 1232
rect 331128 1148 331180 1154
rect 331128 1090 331180 1096
rect 330392 604 330444 610
rect 330392 546 330444 552
rect 330404 480 330432 546
rect 331600 480 331628 1226
rect 332692 1216 332744 1222
rect 332692 1158 332744 1164
rect 332704 480 332732 1158
rect 333532 746 333560 3726
rect 334728 1290 334756 3726
rect 335924 1358 335952 3726
rect 335084 1352 335136 1358
rect 335084 1294 335136 1300
rect 335912 1352 335964 1358
rect 335912 1294 335964 1300
rect 334716 1284 334768 1290
rect 334716 1226 334768 1232
rect 333888 1148 333940 1154
rect 333888 1090 333940 1096
rect 333520 740 333572 746
rect 333520 682 333572 688
rect 333900 480 333928 1090
rect 335096 480 335124 1294
rect 337028 1222 337056 3726
rect 337476 1284 337528 1290
rect 337476 1226 337528 1232
rect 337016 1216 337068 1222
rect 337016 1158 337068 1164
rect 336280 740 336332 746
rect 336280 682 336332 688
rect 336292 480 336320 682
rect 337488 480 337516 1226
rect 338224 746 338252 3726
rect 339328 1358 339356 3726
rect 338672 1352 338724 1358
rect 338672 1294 338724 1300
rect 339316 1352 339368 1358
rect 339316 1294 339368 1300
rect 338212 740 338264 746
rect 338212 682 338264 688
rect 338684 480 338712 1294
rect 340524 1290 340552 3726
rect 340512 1284 340564 1290
rect 340512 1226 340564 1232
rect 341720 1222 341748 3726
rect 342168 1352 342220 1358
rect 342168 1294 342220 1300
rect 339868 1216 339920 1222
rect 339868 1158 339920 1164
rect 341708 1216 341760 1222
rect 341708 1158 341760 1164
rect 339880 480 339908 1158
rect 340972 740 341024 746
rect 340972 682 341024 688
rect 340984 480 341012 682
rect 342180 480 342208 1294
rect 342824 746 342852 3726
rect 344020 1290 344048 3726
rect 345124 1358 345152 3726
rect 345112 1352 345164 1358
rect 345112 1294 345164 1300
rect 343364 1284 343416 1290
rect 343364 1226 343416 1232
rect 344008 1284 344060 1290
rect 344008 1226 344060 1232
rect 342812 740 342864 746
rect 342812 682 342864 688
rect 343376 480 343404 1226
rect 344560 1216 344612 1222
rect 344560 1158 344612 1164
rect 344572 480 344600 1158
rect 346320 746 346348 3726
rect 346952 1284 347004 1290
rect 346952 1226 347004 1232
rect 345756 740 345808 746
rect 345756 682 345808 688
rect 346308 740 346360 746
rect 346308 682 346360 688
rect 345768 480 345796 682
rect 346964 480 346992 1226
rect 347516 882 347544 3726
rect 348056 1352 348108 1358
rect 348056 1294 348108 1300
rect 347504 876 347556 882
rect 347504 818 347556 824
rect 348068 480 348096 1294
rect 348620 1290 348648 3726
rect 349816 1358 349844 3726
rect 349804 1352 349856 1358
rect 349804 1294 349856 1300
rect 348608 1284 348660 1290
rect 348608 1226 348660 1232
rect 350448 876 350500 882
rect 350448 818 350500 824
rect 349252 740 349304 746
rect 349252 682 349304 688
rect 349264 480 349292 682
rect 350460 480 350488 818
rect 350920 746 350948 3726
rect 352116 1290 352144 3726
rect 353220 3726 353292 3754
rect 354368 3754 354396 4012
rect 355564 3754 355592 4012
rect 356668 3754 356696 4012
rect 357864 3754 357892 4012
rect 359060 3754 359088 4012
rect 360164 3754 360192 4012
rect 354368 3726 354444 3754
rect 355564 3726 355640 3754
rect 356668 3726 356744 3754
rect 357864 3726 357940 3754
rect 359060 3726 359136 3754
rect 353220 1358 353248 3726
rect 352840 1352 352892 1358
rect 352840 1294 352892 1300
rect 353208 1352 353260 1358
rect 353208 1294 353260 1300
rect 351644 1284 351696 1290
rect 351644 1226 351696 1232
rect 352104 1284 352156 1290
rect 352104 1226 352156 1232
rect 350908 740 350960 746
rect 350908 682 350960 688
rect 351656 480 351684 1226
rect 352852 480 352880 1294
rect 354036 740 354088 746
rect 354036 682 354088 688
rect 354048 480 354076 682
rect 248758 354 248870 480
rect 248616 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 354416 66 354444 3726
rect 355612 1290 355640 3726
rect 356716 1358 356744 3726
rect 356336 1352 356388 1358
rect 356336 1294 356388 1300
rect 356704 1352 356756 1358
rect 356704 1294 356756 1300
rect 355232 1284 355284 1290
rect 355232 1226 355284 1232
rect 355600 1284 355652 1290
rect 355600 1226 355652 1232
rect 355244 480 355272 1226
rect 356348 480 356376 1294
rect 357912 1222 357940 3726
rect 359108 1290 359136 3726
rect 360120 3726 360192 3754
rect 361360 3754 361388 4012
rect 362556 3754 362584 4012
rect 363660 3754 363688 4012
rect 364856 3754 364884 4012
rect 365960 3754 365988 4012
rect 367156 3754 367184 4012
rect 368352 3754 368380 4012
rect 369456 3754 369484 4012
rect 370652 3754 370680 4012
rect 371756 3754 371784 4012
rect 372952 3754 372980 4012
rect 374148 3754 374176 4012
rect 375252 3754 375280 4012
rect 376448 3754 376476 4012
rect 361360 3726 361436 3754
rect 362556 3726 362632 3754
rect 363660 3726 363736 3754
rect 364856 3726 364932 3754
rect 365960 3726 366036 3754
rect 367156 3726 367232 3754
rect 368352 3726 368428 3754
rect 369456 3726 369532 3754
rect 370652 3726 370728 3754
rect 371756 3726 371832 3754
rect 372952 3726 373028 3754
rect 374148 3726 374224 3754
rect 375252 3726 375328 3754
rect 359924 1352 359976 1358
rect 359924 1294 359976 1300
rect 358728 1284 358780 1290
rect 358728 1226 358780 1232
rect 359096 1284 359148 1290
rect 359096 1226 359148 1232
rect 357900 1216 357952 1222
rect 357900 1158 357952 1164
rect 358740 480 358768 1226
rect 359936 480 359964 1294
rect 360120 1154 360148 3726
rect 361120 1216 361172 1222
rect 361120 1158 361172 1164
rect 360108 1148 360160 1154
rect 360108 1090 360160 1096
rect 361132 480 361160 1158
rect 361408 882 361436 3726
rect 362604 1358 362632 3726
rect 362592 1352 362644 1358
rect 362592 1294 362644 1300
rect 363708 1290 363736 3726
rect 362316 1284 362368 1290
rect 362316 1226 362368 1232
rect 363696 1284 363748 1290
rect 363696 1226 363748 1232
rect 361396 876 361448 882
rect 361396 818 361448 824
rect 362328 480 362356 1226
rect 364904 1222 364932 3726
rect 365812 1352 365864 1358
rect 365812 1294 365864 1300
rect 364892 1216 364944 1222
rect 364892 1158 364944 1164
rect 363512 1148 363564 1154
rect 363512 1090 363564 1096
rect 363524 480 363552 1090
rect 364616 876 364668 882
rect 364616 818 364668 824
rect 364628 480 364656 818
rect 365824 480 365852 1294
rect 366008 746 366036 3726
rect 367204 1358 367232 3726
rect 367192 1352 367244 1358
rect 367192 1294 367244 1300
rect 367008 1284 367060 1290
rect 367008 1226 367060 1232
rect 365996 740 366048 746
rect 365996 682 366048 688
rect 367020 480 367048 1226
rect 368204 1216 368256 1222
rect 368204 1158 368256 1164
rect 368216 480 368244 1158
rect 368400 882 368428 3726
rect 368388 876 368440 882
rect 368388 818 368440 824
rect 369504 746 369532 3726
rect 370700 1358 370728 3726
rect 370596 1352 370648 1358
rect 370596 1294 370648 1300
rect 370688 1352 370740 1358
rect 370688 1294 370740 1300
rect 369400 740 369452 746
rect 369400 682 369452 688
rect 369492 740 369544 746
rect 369492 682 369544 688
rect 369412 480 369440 682
rect 370608 480 370636 1294
rect 371804 882 371832 3726
rect 373000 1290 373028 3726
rect 374092 1352 374144 1358
rect 374092 1294 374144 1300
rect 372988 1284 373040 1290
rect 372988 1226 373040 1232
rect 371700 876 371752 882
rect 371700 818 371752 824
rect 371792 876 371844 882
rect 371792 818 371844 824
rect 371712 480 371740 818
rect 372896 740 372948 746
rect 372896 682 372948 688
rect 372908 480 372936 682
rect 374104 480 374132 1294
rect 374196 1018 374224 3726
rect 375300 1222 375328 3726
rect 376404 3726 376476 3754
rect 377552 3754 377580 4012
rect 378748 3754 378776 4012
rect 379944 3754 379972 4012
rect 377552 3726 377628 3754
rect 378748 3726 378824 3754
rect 376404 1358 376432 3726
rect 376392 1352 376444 1358
rect 376392 1294 376444 1300
rect 377600 1290 377628 3726
rect 376484 1284 376536 1290
rect 376484 1226 376536 1232
rect 377588 1284 377640 1290
rect 377588 1226 377640 1232
rect 375288 1216 375340 1222
rect 375288 1158 375340 1164
rect 374184 1012 374236 1018
rect 374184 954 374236 960
rect 375288 876 375340 882
rect 375288 818 375340 824
rect 375300 480 375328 818
rect 376496 480 376524 1226
rect 378796 1086 378824 3726
rect 379900 3726 379972 3754
rect 381048 3754 381076 4012
rect 382244 3754 382272 4012
rect 381048 3726 381124 3754
rect 378876 1216 378928 1222
rect 378876 1158 378928 1164
rect 378784 1080 378836 1086
rect 378784 1022 378836 1028
rect 377680 1012 377732 1018
rect 377680 954 377732 960
rect 377692 480 377720 954
rect 378888 480 378916 1158
rect 379900 1018 379928 3726
rect 379980 1352 380032 1358
rect 379980 1294 380032 1300
rect 379888 1012 379940 1018
rect 379888 954 379940 960
rect 379992 480 380020 1294
rect 381096 1222 381124 3726
rect 382200 3726 382272 3754
rect 383348 3754 383376 4012
rect 384544 3754 384572 4012
rect 385740 3754 385768 4012
rect 386844 3754 386872 4012
rect 388040 3754 388068 4012
rect 389236 3754 389264 4012
rect 390340 3754 390368 4012
rect 391536 3754 391564 4012
rect 392640 3754 392668 4012
rect 393836 3754 393864 4012
rect 395032 3754 395060 4012
rect 396136 3754 396164 4012
rect 397332 3754 397360 4012
rect 398436 3754 398464 4012
rect 399632 3754 399660 4012
rect 400828 3754 400856 4012
rect 401932 3754 401960 4012
rect 403128 3754 403156 4012
rect 404232 3754 404260 4012
rect 405428 3754 405456 4012
rect 406624 3754 406652 4012
rect 407728 3754 407756 4012
rect 408924 3754 408952 4012
rect 410028 3754 410056 4012
rect 411224 3754 411252 4012
rect 383348 3726 383424 3754
rect 384544 3726 384620 3754
rect 385740 3726 385816 3754
rect 386844 3726 386920 3754
rect 388040 3726 388116 3754
rect 389236 3726 389312 3754
rect 390340 3726 390416 3754
rect 391536 3726 391612 3754
rect 392640 3726 392716 3754
rect 393836 3726 393912 3754
rect 395032 3726 395108 3754
rect 396136 3726 396212 3754
rect 397332 3726 397408 3754
rect 398436 3726 398512 3754
rect 399632 3726 399708 3754
rect 400828 3726 400904 3754
rect 401932 3726 402008 3754
rect 403128 3726 403204 3754
rect 404232 3726 404308 3754
rect 405428 3726 405504 3754
rect 406624 3726 406700 3754
rect 407728 3726 407804 3754
rect 408924 3726 409000 3754
rect 410028 3726 410104 3754
rect 381176 1284 381228 1290
rect 381176 1226 381228 1232
rect 381084 1216 381136 1222
rect 381084 1158 381136 1164
rect 381188 480 381216 1226
rect 382200 1154 382228 3726
rect 382188 1148 382240 1154
rect 382188 1090 382240 1096
rect 382372 1080 382424 1086
rect 382372 1022 382424 1028
rect 382384 480 382412 1022
rect 354404 60 354456 66
rect 354404 2 354456 8
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 82 357614 480
rect 357360 66 357614 82
rect 357348 60 357614 66
rect 357400 54 357614 60
rect 357348 2 357400 8
rect 357502 -960 357614 54
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383396 338 383424 3726
rect 383568 1012 383620 1018
rect 383568 954 383620 960
rect 383580 480 383608 954
rect 384592 882 384620 3726
rect 385788 1358 385816 3726
rect 385776 1352 385828 1358
rect 385776 1294 385828 1300
rect 384764 1216 384816 1222
rect 384764 1158 384816 1164
rect 384580 876 384632 882
rect 384580 818 384632 824
rect 384776 480 384804 1158
rect 385960 1148 386012 1154
rect 385960 1090 386012 1096
rect 385972 480 386000 1090
rect 386892 1086 386920 3726
rect 388088 1290 388116 3726
rect 388076 1284 388128 1290
rect 388076 1226 388128 1232
rect 389284 1154 389312 3726
rect 389456 1352 389508 1358
rect 389456 1294 389508 1300
rect 389272 1148 389324 1154
rect 389272 1090 389324 1096
rect 386880 1080 386932 1086
rect 386880 1022 386932 1028
rect 388260 876 388312 882
rect 388260 818 388312 824
rect 388272 480 388300 818
rect 389468 480 389496 1294
rect 390388 1222 390416 3726
rect 390376 1216 390428 1222
rect 390376 1158 390428 1164
rect 390652 1080 390704 1086
rect 390652 1022 390704 1028
rect 390664 480 390692 1022
rect 391584 882 391612 3726
rect 391848 1284 391900 1290
rect 391848 1226 391900 1232
rect 391572 876 391624 882
rect 391572 818 391624 824
rect 391860 480 391888 1226
rect 383384 332 383436 338
rect 383384 274 383436 280
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 354 387238 480
rect 386800 338 387238 354
rect 386788 332 387238 338
rect 386840 326 387238 332
rect 386788 274 386840 280
rect 387126 -960 387238 326
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392688 134 392716 3726
rect 393884 1290 393912 3726
rect 395080 1358 395108 3726
rect 395068 1352 395120 1358
rect 395068 1294 395120 1300
rect 393872 1284 393924 1290
rect 393872 1226 393924 1232
rect 396184 1222 396212 3726
rect 394240 1216 394292 1222
rect 394240 1158 394292 1164
rect 396172 1216 396224 1222
rect 396172 1158 396224 1164
rect 393044 1148 393096 1154
rect 393044 1090 393096 1096
rect 393056 480 393084 1090
rect 394252 480 394280 1158
rect 397380 882 397408 3726
rect 397736 1284 397788 1290
rect 397736 1226 397788 1232
rect 395344 876 395396 882
rect 395344 818 395396 824
rect 397368 876 397420 882
rect 397368 818 397420 824
rect 395356 480 395384 818
rect 397748 480 397776 1226
rect 398484 1154 398512 3726
rect 399680 1358 399708 3726
rect 398932 1352 398984 1358
rect 398932 1294 398984 1300
rect 399668 1352 399720 1358
rect 399668 1294 399720 1300
rect 398472 1148 398524 1154
rect 398472 1090 398524 1096
rect 398944 480 398972 1294
rect 400876 1222 400904 3726
rect 400128 1216 400180 1222
rect 400128 1158 400180 1164
rect 400864 1216 400916 1222
rect 400864 1158 400916 1164
rect 400140 480 400168 1158
rect 401324 876 401376 882
rect 401324 818 401376 824
rect 401336 480 401364 818
rect 392676 128 392728 134
rect 392676 70 392728 76
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396172 128 396224 134
rect 396510 82 396622 480
rect 396224 76 396622 82
rect 396172 70 396622 76
rect 396184 54 396622 70
rect 396510 -960 396622 54
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 401980 134 402008 3726
rect 403176 1290 403204 3726
rect 403624 1352 403676 1358
rect 403624 1294 403676 1300
rect 403164 1284 403216 1290
rect 403164 1226 403216 1232
rect 402520 1148 402572 1154
rect 402520 1090 402572 1096
rect 402532 480 402560 1090
rect 403636 480 403664 1294
rect 404280 1154 404308 3726
rect 405476 1358 405504 3726
rect 405464 1352 405516 1358
rect 405464 1294 405516 1300
rect 404820 1216 404872 1222
rect 404820 1158 404872 1164
rect 404268 1148 404320 1154
rect 404268 1090 404320 1096
rect 404832 480 404860 1158
rect 406672 882 406700 3726
rect 407212 1284 407264 1290
rect 407212 1226 407264 1232
rect 406660 876 406712 882
rect 406660 818 406712 824
rect 407224 480 407252 1226
rect 407776 1222 407804 3726
rect 407764 1216 407816 1222
rect 407764 1158 407816 1164
rect 408972 1154 409000 3726
rect 409604 1352 409656 1358
rect 409604 1294 409656 1300
rect 408408 1148 408460 1154
rect 408408 1090 408460 1096
rect 408960 1148 409012 1154
rect 408960 1090 409012 1096
rect 408420 480 408448 1090
rect 409616 480 409644 1294
rect 410076 1290 410104 3726
rect 411180 3726 411252 3754
rect 412420 3754 412448 4012
rect 413524 3754 413552 4012
rect 414720 3754 414748 4012
rect 415916 3754 415944 4012
rect 417020 3754 417048 4012
rect 418216 3754 418244 4012
rect 419320 3754 419348 4012
rect 420516 3754 420544 4012
rect 421712 3754 421740 4012
rect 422816 3754 422844 4012
rect 424012 3754 424040 4012
rect 425116 3754 425144 4012
rect 426312 3754 426340 4012
rect 427508 3754 427536 4012
rect 428612 3754 428640 4012
rect 429808 3754 429836 4012
rect 430912 3754 430940 4012
rect 432108 3754 432136 4012
rect 433304 3754 433332 4012
rect 434408 3754 434436 4012
rect 412420 3726 412496 3754
rect 413524 3726 413600 3754
rect 414720 3726 414796 3754
rect 415916 3726 415992 3754
rect 417020 3726 417096 3754
rect 418216 3726 418292 3754
rect 419320 3726 419396 3754
rect 420516 3726 420592 3754
rect 421712 3726 421788 3754
rect 422816 3726 422892 3754
rect 424012 3726 424088 3754
rect 425116 3726 425192 3754
rect 426312 3726 426388 3754
rect 427508 3726 427584 3754
rect 428612 3726 428688 3754
rect 429808 3726 429884 3754
rect 430912 3726 431080 3754
rect 432108 3726 432184 3754
rect 411180 2854 411208 3726
rect 411168 2848 411220 2854
rect 411168 2790 411220 2796
rect 410064 1284 410116 1290
rect 410064 1226 410116 1232
rect 411904 1216 411956 1222
rect 411904 1158 411956 1164
rect 410800 876 410852 882
rect 410800 818 410852 824
rect 410812 480 410840 818
rect 411916 480 411944 1158
rect 401968 128 402020 134
rect 401968 70 402020 76
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 82 406098 480
rect 406200 128 406252 134
rect 405986 76 406200 82
rect 405986 70 406252 76
rect 405986 54 406240 70
rect 405986 -960 406098 54
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412468 202 412496 3726
rect 413572 1358 413600 3726
rect 413560 1352 413612 1358
rect 413560 1294 413612 1300
rect 414296 1284 414348 1290
rect 414296 1226 414348 1232
rect 413100 1148 413152 1154
rect 413100 1090 413152 1096
rect 413112 480 413140 1090
rect 414308 480 414336 1226
rect 414768 1018 414796 3726
rect 415492 2848 415544 2854
rect 415492 2790 415544 2796
rect 414756 1012 414808 1018
rect 414756 954 414808 960
rect 415504 480 415532 2790
rect 415964 1154 415992 3726
rect 415952 1148 416004 1154
rect 415952 1090 416004 1096
rect 417068 1086 417096 3726
rect 417884 1352 417936 1358
rect 417884 1294 417936 1300
rect 417056 1080 417108 1086
rect 417056 1022 417108 1028
rect 417896 480 417924 1294
rect 418264 1290 418292 3726
rect 418252 1284 418304 1290
rect 418252 1226 418304 1232
rect 418988 1012 419040 1018
rect 418988 954 419040 960
rect 419000 480 419028 954
rect 419368 882 419396 3726
rect 420564 1222 420592 3726
rect 420552 1216 420604 1222
rect 420552 1158 420604 1164
rect 420184 1148 420236 1154
rect 420184 1090 420236 1096
rect 419356 876 419408 882
rect 419356 818 419408 824
rect 420196 480 420224 1090
rect 421380 1080 421432 1086
rect 421380 1022 421432 1028
rect 421392 480 421420 1022
rect 412456 196 412508 202
rect 412456 138 412508 144
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 218 416770 480
rect 416658 202 416912 218
rect 416658 196 416924 202
rect 416658 190 416872 196
rect 416658 -960 416770 190
rect 416872 138 416924 144
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 421760 134 421788 3726
rect 422864 1358 422892 3726
rect 422852 1352 422904 1358
rect 422852 1294 422904 1300
rect 422576 1284 422628 1290
rect 422576 1226 422628 1232
rect 422588 480 422616 1226
rect 424060 1018 424088 3726
rect 425164 1222 425192 3726
rect 426360 1290 426388 3726
rect 427556 1358 427584 3726
rect 427268 1352 427320 1358
rect 427268 1294 427320 1300
rect 427544 1352 427596 1358
rect 427544 1294 427596 1300
rect 426348 1284 426400 1290
rect 426348 1226 426400 1232
rect 424968 1216 425020 1222
rect 424968 1158 425020 1164
rect 425152 1216 425204 1222
rect 425152 1158 425204 1164
rect 424048 1012 424100 1018
rect 424048 954 424100 960
rect 423404 876 423456 882
rect 423404 818 423456 824
rect 421748 128 421800 134
rect 421748 70 421800 76
rect 422546 -960 422658 480
rect 423416 354 423444 818
rect 424980 480 425008 1158
rect 427280 480 427308 1294
rect 428660 1154 428688 3726
rect 429660 1216 429712 1222
rect 429660 1158 429712 1164
rect 428648 1148 428700 1154
rect 428648 1090 428700 1096
rect 428464 1012 428516 1018
rect 428464 954 428516 960
rect 428476 480 428504 954
rect 429672 480 429700 1158
rect 429856 882 429884 3726
rect 430856 1284 430908 1290
rect 430856 1226 430908 1232
rect 429844 876 429896 882
rect 429844 818 429896 824
rect 430868 480 430896 1226
rect 423742 354 423854 480
rect 423416 326 423854 354
rect 423742 -960 423854 326
rect 424938 -960 425050 480
rect 425796 128 425848 134
rect 426134 82 426246 480
rect 425848 76 426246 82
rect 425796 70 426246 76
rect 425808 54 426246 70
rect 426134 -960 426246 54
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 431052 134 431080 3726
rect 431868 1352 431920 1358
rect 431868 1294 431920 1300
rect 431880 354 431908 1294
rect 432156 1018 432184 3726
rect 433260 3726 433332 3754
rect 434364 3726 434436 3754
rect 435604 3754 435632 4012
rect 436708 3754 436736 4012
rect 437904 3754 437932 4012
rect 439100 3754 439128 4012
rect 440204 3754 440232 4012
rect 435604 3726 435680 3754
rect 436708 3726 436784 3754
rect 437904 3726 437980 3754
rect 439100 3726 439176 3754
rect 433260 1358 433288 3726
rect 433248 1352 433300 1358
rect 433248 1294 433300 1300
rect 433248 1148 433300 1154
rect 433248 1090 433300 1096
rect 432144 1012 432196 1018
rect 432144 954 432196 960
rect 433260 480 433288 1090
rect 434364 950 434392 3726
rect 435652 1290 435680 3726
rect 435640 1284 435692 1290
rect 435640 1226 435692 1232
rect 436756 1222 436784 3726
rect 437848 1352 437900 1358
rect 437848 1294 437900 1300
rect 436744 1216 436796 1222
rect 436744 1158 436796 1164
rect 436744 1012 436796 1018
rect 436744 954 436796 960
rect 434352 944 434404 950
rect 434352 886 434404 892
rect 434444 876 434496 882
rect 434444 818 434496 824
rect 434456 480 434484 818
rect 436756 480 436784 954
rect 437860 898 437888 1294
rect 437952 1086 437980 3726
rect 439148 1154 439176 3726
rect 440160 3726 440232 3754
rect 441400 3754 441428 4012
rect 442596 3754 442624 4012
rect 443700 3754 443728 4012
rect 444896 3754 444924 4012
rect 446000 3754 446028 4012
rect 447196 3754 447224 4012
rect 448392 3754 448420 4012
rect 449496 3754 449524 4012
rect 450692 3754 450720 4012
rect 451796 3754 451824 4012
rect 452992 3754 453020 4012
rect 454188 3754 454216 4012
rect 455292 3754 455320 4012
rect 456488 3754 456516 4012
rect 457592 3754 457620 4012
rect 458788 3754 458816 4012
rect 459984 3754 460012 4012
rect 461088 3754 461116 4012
rect 462284 3754 462312 4012
rect 441400 3726 441476 3754
rect 442596 3726 442672 3754
rect 443700 3726 443776 3754
rect 444896 3726 444972 3754
rect 446000 3726 446076 3754
rect 447196 3726 447272 3754
rect 448392 3726 448468 3754
rect 449496 3726 449572 3754
rect 450692 3726 450768 3754
rect 451796 3726 451872 3754
rect 452992 3726 453068 3754
rect 454188 3726 454264 3754
rect 455292 3726 455368 3754
rect 456488 3726 456564 3754
rect 457592 3726 457668 3754
rect 458788 3726 458864 3754
rect 459984 3726 460060 3754
rect 461088 3726 461164 3754
rect 440160 2854 440188 3726
rect 440148 2848 440200 2854
rect 440148 2790 440200 2796
rect 441448 1358 441476 3726
rect 441436 1352 441488 1358
rect 441436 1294 441488 1300
rect 442644 1290 442672 3726
rect 439964 1284 440016 1290
rect 439964 1226 440016 1232
rect 442632 1284 442684 1290
rect 442632 1226 442684 1232
rect 439136 1148 439188 1154
rect 439136 1090 439188 1096
rect 437940 1080 437992 1086
rect 437940 1022 437992 1028
rect 439136 944 439188 950
rect 437860 870 437980 898
rect 439136 886 439188 892
rect 437952 480 437980 870
rect 439148 480 439176 886
rect 432022 354 432134 480
rect 431880 326 432134 354
rect 431040 128 431092 134
rect 431040 70 431092 76
rect 432022 -960 432134 326
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435180 128 435232 134
rect 435518 82 435630 480
rect 435232 76 435630 82
rect 435180 70 435630 76
rect 435192 54 435630 70
rect 435518 -960 435630 54
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 439976 354 440004 1226
rect 441528 1216 441580 1222
rect 441528 1158 441580 1164
rect 441540 480 441568 1158
rect 442632 1080 442684 1086
rect 442632 1022 442684 1028
rect 442644 480 442672 1022
rect 443748 882 443776 3726
rect 444944 1222 444972 3726
rect 445024 2848 445076 2854
rect 445024 2790 445076 2796
rect 444932 1216 444984 1222
rect 444932 1158 444984 1164
rect 443828 1148 443880 1154
rect 443828 1090 443880 1096
rect 443736 876 443788 882
rect 443736 818 443788 824
rect 443840 480 443868 1090
rect 445036 480 445064 2790
rect 445852 1352 445904 1358
rect 445852 1294 445904 1300
rect 440302 354 440414 480
rect 439976 326 440414 354
rect 440302 -960 440414 326
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445864 354 445892 1294
rect 446048 1086 446076 3726
rect 447244 1358 447272 3726
rect 447232 1352 447284 1358
rect 447232 1294 447284 1300
rect 447416 1284 447468 1290
rect 447416 1226 447468 1232
rect 446036 1080 446088 1086
rect 446036 1022 446088 1028
rect 447428 480 447456 1226
rect 448440 1154 448468 3726
rect 449544 2854 449572 3726
rect 449532 2848 449584 2854
rect 449532 2790 449584 2796
rect 450740 1222 450768 3726
rect 449808 1216 449860 1222
rect 449808 1158 449860 1164
rect 450728 1216 450780 1222
rect 450728 1158 450780 1164
rect 448428 1148 448480 1154
rect 448428 1090 448480 1096
rect 448244 876 448296 882
rect 448244 818 448296 824
rect 446190 354 446302 480
rect 445864 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448256 354 448284 818
rect 449820 480 449848 1158
rect 450912 1080 450964 1086
rect 450912 1022 450964 1028
rect 450924 480 450952 1022
rect 451844 882 451872 3726
rect 453040 1358 453068 3726
rect 452108 1352 452160 1358
rect 452108 1294 452160 1300
rect 453028 1352 453080 1358
rect 453028 1294 453080 1300
rect 451832 876 451884 882
rect 451832 818 451884 824
rect 452120 480 452148 1294
rect 454236 1154 454264 3726
rect 454500 2848 454552 2854
rect 454500 2790 454552 2796
rect 453304 1148 453356 1154
rect 453304 1090 453356 1096
rect 454224 1148 454276 1154
rect 454224 1090 454276 1096
rect 453316 480 453344 1090
rect 454512 480 454540 2790
rect 455340 1086 455368 3726
rect 456536 1222 456564 3726
rect 457640 1290 457668 3726
rect 458836 1358 458864 3726
rect 458088 1352 458140 1358
rect 458088 1294 458140 1300
rect 458824 1352 458876 1358
rect 458824 1294 458876 1300
rect 457628 1284 457680 1290
rect 457628 1226 457680 1232
rect 455696 1216 455748 1222
rect 455696 1158 455748 1164
rect 456524 1216 456576 1222
rect 456524 1158 456576 1164
rect 455328 1080 455380 1086
rect 455328 1022 455380 1028
rect 455708 480 455736 1158
rect 456524 876 456576 882
rect 456524 818 456576 824
rect 448582 354 448694 480
rect 448256 326 448694 354
rect 448582 -960 448694 326
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456536 354 456564 818
rect 458100 480 458128 1294
rect 459192 1148 459244 1154
rect 459192 1090 459244 1096
rect 459204 480 459232 1090
rect 456862 354 456974 480
rect 456536 326 456974 354
rect 456862 -960 456974 326
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460032 134 460060 3726
rect 461136 1086 461164 3726
rect 462240 3726 462312 3754
rect 463388 3754 463416 4012
rect 464584 3754 464612 4012
rect 465780 3754 465808 4012
rect 466884 3754 466912 4012
rect 468080 3754 468108 4012
rect 469276 3754 469304 4012
rect 470380 3754 470408 4012
rect 471576 3754 471604 4012
rect 472680 3754 472708 4012
rect 473876 3754 473904 4012
rect 475072 3754 475100 4012
rect 476176 3754 476204 4012
rect 477372 3754 477400 4012
rect 478476 3754 478504 4012
rect 479672 3754 479700 4012
rect 480868 3754 480896 4012
rect 481972 3754 482000 4012
rect 483168 3754 483196 4012
rect 484272 3754 484300 4012
rect 485468 3754 485496 4012
rect 486664 3754 486692 4012
rect 487768 3754 487796 4012
rect 488964 3754 488992 4012
rect 490068 3754 490096 4012
rect 491264 3754 491292 4012
rect 463388 3726 463464 3754
rect 464584 3726 464660 3754
rect 465780 3726 465856 3754
rect 466884 3726 466960 3754
rect 468080 3726 468156 3754
rect 469276 3726 469352 3754
rect 470380 3726 470456 3754
rect 471576 3726 471652 3754
rect 472680 3726 472756 3754
rect 473876 3726 473952 3754
rect 475072 3726 475148 3754
rect 476176 3726 476252 3754
rect 477372 3726 477448 3754
rect 478476 3726 478552 3754
rect 479672 3726 479748 3754
rect 480868 3726 480944 3754
rect 481972 3726 482048 3754
rect 483168 3726 483244 3754
rect 484272 3726 484348 3754
rect 485468 3726 485544 3754
rect 486664 3726 486740 3754
rect 487768 3726 487844 3754
rect 488964 3726 489040 3754
rect 490068 3726 490144 3754
rect 462240 1222 462268 3726
rect 462412 1284 462464 1290
rect 462412 1226 462464 1232
rect 461584 1216 461636 1222
rect 461584 1158 461636 1164
rect 462228 1216 462280 1222
rect 462228 1158 462280 1164
rect 460112 1080 460164 1086
rect 460112 1022 460164 1028
rect 461124 1080 461176 1086
rect 461124 1022 461176 1028
rect 460124 354 460152 1022
rect 461596 480 461624 1158
rect 460358 354 460470 480
rect 460124 326 460470 354
rect 460020 128 460072 134
rect 460020 70 460072 76
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462424 354 462452 1226
rect 463436 950 463464 3726
rect 463976 1352 464028 1358
rect 463976 1294 464028 1300
rect 463424 944 463476 950
rect 463424 886 463476 892
rect 463988 480 464016 1294
rect 464632 1018 464660 3726
rect 465828 1154 465856 3726
rect 465816 1148 465868 1154
rect 465816 1090 465868 1096
rect 466932 1086 466960 3726
rect 468128 1290 468156 3726
rect 468116 1284 468168 1290
rect 468116 1226 468168 1232
rect 467472 1216 467524 1222
rect 467472 1158 467524 1164
rect 466276 1080 466328 1086
rect 466276 1022 466328 1028
rect 466920 1080 466972 1086
rect 466920 1022 466972 1028
rect 464620 1012 464672 1018
rect 464620 954 464672 960
rect 466288 480 466316 1022
rect 467484 480 467512 1158
rect 468668 944 468720 950
rect 468668 886 468720 892
rect 468680 480 468708 886
rect 462750 354 462862 480
rect 462424 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 464988 128 465040 134
rect 465142 82 465254 480
rect 465040 76 465254 82
rect 464988 70 465254 76
rect 465000 54 465254 70
rect 465142 -960 465254 54
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469324 270 469352 3726
rect 469864 1012 469916 1018
rect 469864 954 469916 960
rect 469876 480 469904 954
rect 469312 264 469364 270
rect 469312 206 469364 212
rect 469834 -960 469946 480
rect 470428 202 470456 3726
rect 471624 1358 471652 3726
rect 471612 1352 471664 1358
rect 471612 1294 471664 1300
rect 472728 1222 472756 3726
rect 473084 1284 473136 1290
rect 473084 1226 473136 1232
rect 472716 1216 472768 1222
rect 472716 1158 472768 1164
rect 470692 1148 470744 1154
rect 470692 1090 470744 1096
rect 470704 354 470732 1090
rect 472256 1080 472308 1086
rect 472256 1022 472308 1028
rect 472268 480 472296 1022
rect 471030 354 471142 480
rect 470704 326 471142 354
rect 470416 196 470468 202
rect 470416 138 470468 144
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473096 354 473124 1226
rect 473924 1018 473952 3726
rect 475120 1290 475148 3726
rect 475108 1284 475160 1290
rect 475108 1226 475160 1232
rect 473912 1012 473964 1018
rect 473912 954 473964 960
rect 476224 882 476252 3726
rect 477420 1358 477448 3726
rect 478524 2854 478552 3726
rect 478512 2848 478564 2854
rect 478512 2790 478564 2796
rect 476580 1352 476632 1358
rect 476580 1294 476632 1300
rect 477408 1352 477460 1358
rect 477408 1294 477460 1300
rect 476212 876 476264 882
rect 476212 818 476264 824
rect 473422 354 473534 480
rect 473096 326 473534 354
rect 473422 -960 473534 326
rect 474188 264 474240 270
rect 474526 218 474638 480
rect 474240 212 474638 218
rect 474188 206 474638 212
rect 474200 190 474638 206
rect 474526 -960 474638 190
rect 475722 218 475834 480
rect 476592 354 476620 1294
rect 478144 1216 478196 1222
rect 478144 1158 478196 1164
rect 478156 480 478184 1158
rect 479720 1086 479748 3726
rect 480536 1284 480588 1290
rect 480536 1226 480588 1232
rect 479708 1080 479760 1086
rect 479708 1022 479760 1028
rect 479340 1012 479392 1018
rect 479340 954 479392 960
rect 479352 480 479380 954
rect 480548 480 480576 1226
rect 480916 1222 480944 3726
rect 480904 1216 480956 1222
rect 480904 1158 480956 1164
rect 482020 1154 482048 3726
rect 483216 1358 483244 3726
rect 484032 2848 484084 2854
rect 484032 2790 484084 2796
rect 482468 1352 482520 1358
rect 482468 1294 482520 1300
rect 483204 1352 483256 1358
rect 483204 1294 483256 1300
rect 482008 1148 482060 1154
rect 482008 1090 482060 1096
rect 481364 876 481416 882
rect 481364 818 481416 824
rect 476918 354 477030 480
rect 476592 326 477030 354
rect 475722 202 475976 218
rect 475722 196 475988 202
rect 475722 190 475936 196
rect 475722 -960 475834 190
rect 475936 138 475988 144
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481376 354 481404 818
rect 481702 354 481814 480
rect 481376 326 481814 354
rect 482480 354 482508 1294
rect 484044 480 484072 2790
rect 484320 950 484348 3726
rect 485516 1290 485544 3726
rect 485504 1284 485556 1290
rect 485504 1226 485556 1232
rect 486712 1222 486740 3726
rect 487816 2854 487844 3726
rect 487804 2848 487856 2854
rect 487804 2790 487856 2796
rect 488816 1352 488868 1358
rect 488816 1294 488868 1300
rect 486424 1216 486476 1222
rect 486424 1158 486476 1164
rect 486700 1216 486752 1222
rect 486700 1158 486752 1164
rect 484860 1080 484912 1086
rect 484860 1022 484912 1028
rect 484308 944 484360 950
rect 484308 886 484360 892
rect 482806 354 482918 480
rect 482480 326 482918 354
rect 481702 -960 481814 326
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484872 354 484900 1022
rect 486436 480 486464 1158
rect 487252 1148 487304 1154
rect 487252 1090 487304 1096
rect 485198 354 485310 480
rect 484872 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487264 354 487292 1090
rect 488828 480 488856 1294
rect 489012 1154 489040 3726
rect 490116 1358 490144 3726
rect 491220 3726 491292 3754
rect 492460 3754 492488 4012
rect 493564 3754 493592 4012
rect 494760 3754 494788 4012
rect 495956 3754 495984 4012
rect 497060 3754 497088 4012
rect 498256 3754 498284 4012
rect 499360 3754 499388 4012
rect 492460 3726 492536 3754
rect 493564 3726 493640 3754
rect 494760 3726 494836 3754
rect 495956 3726 496032 3754
rect 497060 3726 497136 3754
rect 498256 3726 498332 3754
rect 490104 1352 490156 1358
rect 490104 1294 490156 1300
rect 490748 1284 490800 1290
rect 490748 1226 490800 1232
rect 489000 1148 489052 1154
rect 489000 1090 489052 1096
rect 489920 944 489972 950
rect 489920 886 489972 892
rect 489932 480 489960 886
rect 487590 354 487702 480
rect 487264 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 1226
rect 491220 1086 491248 3726
rect 492508 1290 492536 3726
rect 493508 2848 493560 2854
rect 493508 2790 493560 2796
rect 492496 1284 492548 1290
rect 492496 1226 492548 1232
rect 492312 1216 492364 1222
rect 492312 1158 492364 1164
rect 491208 1080 491260 1086
rect 491208 1022 491260 1028
rect 492324 480 492352 1158
rect 493520 480 493548 2790
rect 493612 1222 493640 3726
rect 493600 1216 493652 1222
rect 493600 1158 493652 1164
rect 494704 1148 494756 1154
rect 494704 1090 494756 1096
rect 494716 480 494744 1090
rect 494808 678 494836 3726
rect 495532 1352 495584 1358
rect 495532 1294 495584 1300
rect 494796 672 494848 678
rect 494796 614 494848 620
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495544 354 495572 1294
rect 496004 1018 496032 3726
rect 497108 1358 497136 3726
rect 497096 1352 497148 1358
rect 497096 1294 497148 1300
rect 498304 1290 498332 3726
rect 499224 3726 499388 3754
rect 500556 3754 500584 4012
rect 501752 3754 501780 4012
rect 502856 3754 502884 4012
rect 504052 3754 504080 4012
rect 505156 3754 505184 4012
rect 506352 3754 506380 4012
rect 507548 3754 507576 4012
rect 500556 3726 500632 3754
rect 501752 3726 501828 3754
rect 502856 3726 502932 3754
rect 504052 3726 504128 3754
rect 505156 3726 505232 3754
rect 498200 1284 498252 1290
rect 498200 1226 498252 1232
rect 498292 1284 498344 1290
rect 498292 1226 498344 1232
rect 497096 1080 497148 1086
rect 497096 1022 497148 1028
rect 495992 1012 496044 1018
rect 495992 954 496044 960
rect 497108 480 497136 1022
rect 498212 480 498240 1226
rect 495870 354 495982 480
rect 495544 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499224 66 499252 3726
rect 500604 1222 500632 3726
rect 499396 1216 499448 1222
rect 499396 1158 499448 1164
rect 500592 1216 500644 1222
rect 500592 1158 500644 1164
rect 499408 480 499436 1158
rect 501800 1154 501828 3726
rect 501788 1148 501840 1154
rect 501788 1090 501840 1096
rect 502904 1018 502932 3726
rect 504100 1358 504128 3726
rect 502984 1352 503036 1358
rect 502984 1294 503036 1300
rect 504088 1352 504140 1358
rect 504088 1294 504140 1300
rect 501788 1012 501840 1018
rect 501788 954 501840 960
rect 502892 1012 502944 1018
rect 502892 954 502944 960
rect 500592 672 500644 678
rect 500592 614 500644 620
rect 500604 480 500632 614
rect 501800 480 501828 954
rect 502996 480 503024 1294
rect 503812 1284 503864 1290
rect 503812 1226 503864 1232
rect 499212 60 499264 66
rect 499212 2 499264 8
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503824 354 503852 1226
rect 505204 1086 505232 3726
rect 506308 3726 506380 3754
rect 507504 3726 507576 3754
rect 508652 3754 508680 4012
rect 509848 3754 509876 4012
rect 510952 3754 510980 4012
rect 512148 3754 512176 4012
rect 513344 3754 513372 4012
rect 508652 3726 508728 3754
rect 509848 3726 509924 3754
rect 510952 3726 511028 3754
rect 512148 3726 512224 3754
rect 505192 1080 505244 1086
rect 505192 1022 505244 1028
rect 504150 354 504262 480
rect 503824 326 504262 354
rect 504150 -960 504262 326
rect 505346 82 505458 480
rect 505346 66 505600 82
rect 506308 66 506336 3726
rect 506480 1216 506532 1222
rect 506480 1158 506532 1164
rect 506492 480 506520 1158
rect 507308 1148 507360 1154
rect 507308 1090 507360 1096
rect 505346 60 505612 66
rect 505346 54 505560 60
rect 505346 -960 505458 54
rect 505560 2 505612 8
rect 506296 60 506348 66
rect 506296 2 506348 8
rect 506450 -960 506562 480
rect 507320 82 507348 1090
rect 507504 202 507532 3726
rect 507492 196 507544 202
rect 507492 138 507544 144
rect 507646 82 507758 480
rect 508700 270 508728 3726
rect 509896 1358 509924 3726
rect 509700 1352 509752 1358
rect 509700 1294 509752 1300
rect 509884 1352 509936 1358
rect 509884 1294 509936 1300
rect 508872 1012 508924 1018
rect 508872 954 508924 960
rect 508884 480 508912 954
rect 508688 264 508740 270
rect 508688 206 508740 212
rect 507320 54 507758 82
rect 507646 -960 507758 54
rect 508842 -960 508954 480
rect 509712 354 509740 1294
rect 511000 1290 511028 3726
rect 510988 1284 511040 1290
rect 510988 1226 511040 1232
rect 512196 1086 512224 3726
rect 513300 3726 513372 3754
rect 514448 3754 514476 4012
rect 515644 3754 515672 4012
rect 516748 3754 516776 4012
rect 517944 3754 517972 4012
rect 519140 3754 519168 4012
rect 520244 3754 520272 4012
rect 514448 3726 514524 3754
rect 515644 3726 515720 3754
rect 516748 3726 516824 3754
rect 517944 3726 518020 3754
rect 519140 3726 519216 3754
rect 513300 1154 513328 3726
rect 513288 1148 513340 1154
rect 513288 1090 513340 1096
rect 511264 1080 511316 1086
rect 511264 1022 511316 1028
rect 512184 1080 512236 1086
rect 512184 1022 512236 1028
rect 511276 480 511304 1022
rect 514496 882 514524 3726
rect 514484 876 514536 882
rect 514484 818 514536 824
rect 510038 354 510150 480
rect 509712 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512430 82 512542 480
rect 513534 218 513646 480
rect 513392 202 513646 218
rect 513380 196 513646 202
rect 513432 190 513646 196
rect 513380 138 513432 144
rect 512104 66 512542 82
rect 512092 60 512542 66
rect 512144 54 512542 60
rect 512092 2 512144 8
rect 512430 -960 512542 54
rect 513534 -960 513646 190
rect 514730 218 514842 480
rect 514944 264 514996 270
rect 514730 212 514944 218
rect 514730 206 514996 212
rect 514730 190 514984 206
rect 514730 -960 514842 190
rect 515692 134 515720 3726
rect 515772 1352 515824 1358
rect 515772 1294 515824 1300
rect 515784 354 515812 1294
rect 515926 354 516038 480
rect 515784 326 516038 354
rect 515680 128 515732 134
rect 515680 70 515732 76
rect 515926 -960 516038 326
rect 516796 270 516824 3726
rect 517992 1290 518020 3726
rect 519188 1358 519216 3726
rect 520200 3726 520272 3754
rect 521440 3754 521468 4012
rect 522636 3754 522664 4012
rect 523740 3754 523768 4012
rect 524936 3754 524964 4012
rect 526040 3754 526068 4012
rect 527236 3754 527264 4012
rect 528432 3754 528460 4012
rect 529536 3754 529564 4012
rect 530732 3754 530760 4012
rect 531836 3754 531864 4012
rect 533032 3754 533060 4012
rect 534228 3754 534256 4012
rect 535332 3754 535360 4012
rect 536528 3754 536556 4012
rect 537632 3754 537660 4012
rect 538828 3754 538856 4012
rect 540024 3754 540052 4012
rect 541128 3754 541156 4012
rect 542324 3754 542352 4012
rect 521440 3726 521516 3754
rect 522636 3726 522712 3754
rect 523740 3726 523816 3754
rect 524936 3726 525012 3754
rect 526040 3726 526116 3754
rect 527236 3726 527312 3754
rect 528432 3726 528508 3754
rect 529536 3726 529612 3754
rect 530732 3726 530808 3754
rect 531836 3726 531912 3754
rect 533032 3726 533108 3754
rect 534228 3726 534304 3754
rect 535332 3726 535408 3754
rect 536528 3726 536604 3754
rect 537632 3726 537708 3754
rect 538828 3726 538904 3754
rect 540024 3726 540100 3754
rect 541128 3726 541204 3754
rect 519176 1352 519228 1358
rect 519176 1294 519228 1300
rect 517152 1284 517204 1290
rect 517152 1226 517204 1232
rect 517980 1284 518032 1290
rect 517980 1226 518032 1232
rect 517164 480 517192 1226
rect 519544 1148 519596 1154
rect 519544 1090 519596 1096
rect 517980 1080 518032 1086
rect 517980 1022 518032 1028
rect 516784 264 516836 270
rect 516784 206 516836 212
rect 517122 -960 517234 480
rect 517992 354 518020 1022
rect 519556 480 519584 1090
rect 520200 1086 520228 3726
rect 520188 1080 520240 1086
rect 520188 1022 520240 1028
rect 521488 882 521516 3726
rect 522684 1222 522712 3726
rect 522672 1216 522724 1222
rect 522672 1158 522724 1164
rect 523788 1154 523816 3726
rect 523868 1284 523920 1290
rect 523868 1226 523920 1232
rect 523776 1148 523828 1154
rect 523776 1090 523828 1096
rect 520740 876 520792 882
rect 520740 818 520792 824
rect 521476 876 521528 882
rect 521476 818 521528 824
rect 520752 480 520780 818
rect 518318 354 518430 480
rect 517992 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521660 128 521712 134
rect 521814 82 521926 480
rect 521712 76 521926 82
rect 521660 70 521926 76
rect 521672 54 521926 70
rect 521814 -960 521926 54
rect 523010 218 523122 480
rect 523880 354 523908 1226
rect 524206 354 524318 480
rect 523880 326 524318 354
rect 523224 264 523276 270
rect 523010 212 523224 218
rect 523010 206 523276 212
rect 523010 190 523264 206
rect 523010 -960 523122 190
rect 524206 -960 524318 326
rect 524984 134 525012 3726
rect 526088 1358 526116 3726
rect 525432 1352 525484 1358
rect 525432 1294 525484 1300
rect 526076 1352 526128 1358
rect 526076 1294 526128 1300
rect 525444 480 525472 1294
rect 527284 1290 527312 3726
rect 527272 1284 527324 1290
rect 527272 1226 527324 1232
rect 526628 1080 526680 1086
rect 526628 1022 526680 1028
rect 526640 480 526668 1022
rect 527824 876 527876 882
rect 527824 818 527876 824
rect 527836 480 527864 818
rect 524972 128 525024 134
rect 524972 70 525024 76
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528480 66 528508 3726
rect 529020 1216 529072 1222
rect 529020 1158 529072 1164
rect 529032 480 529060 1158
rect 529584 1086 529612 3726
rect 530780 1222 530808 3726
rect 530768 1216 530820 1222
rect 530768 1158 530820 1164
rect 530124 1148 530176 1154
rect 530124 1090 530176 1096
rect 529572 1080 529624 1086
rect 529572 1022 529624 1028
rect 530136 480 530164 1090
rect 531884 610 531912 3726
rect 532148 1352 532200 1358
rect 532148 1294 532200 1300
rect 531872 604 531924 610
rect 531872 546 531924 552
rect 528468 60 528520 66
rect 528468 2 528520 8
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 82 531402 480
rect 532160 354 532188 1294
rect 533080 1154 533108 3726
rect 534276 1358 534304 3726
rect 534264 1352 534316 1358
rect 534264 1294 534316 1300
rect 533712 1284 533764 1290
rect 533712 1226 533764 1232
rect 533068 1148 533120 1154
rect 533068 1090 533120 1096
rect 533724 480 533752 1226
rect 532486 354 532598 480
rect 532160 326 532598 354
rect 531504 128 531556 134
rect 531290 76 531504 82
rect 531290 70 531556 76
rect 531290 54 531544 70
rect 531290 -960 531402 54
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534878 82 534990 480
rect 535380 474 535408 3726
rect 536104 1080 536156 1086
rect 536104 1022 536156 1028
rect 536116 480 536144 1022
rect 535368 468 535420 474
rect 535368 410 535420 416
rect 534552 66 534990 82
rect 534540 60 534990 66
rect 534592 54 534990 60
rect 534540 2 534592 8
rect 534878 -960 534990 54
rect 536074 -960 536186 480
rect 536576 66 536604 3726
rect 537208 1216 537260 1222
rect 537208 1158 537260 1164
rect 537220 480 537248 1158
rect 537680 542 537708 3726
rect 538876 1222 538904 3726
rect 538864 1216 538916 1222
rect 538864 1158 538916 1164
rect 539600 1148 539652 1154
rect 539600 1090 539652 1096
rect 538404 604 538456 610
rect 538404 546 538456 552
rect 537668 536 537720 542
rect 536564 60 536616 66
rect 536564 2 536616 8
rect 537178 -960 537290 480
rect 537668 478 537720 484
rect 538416 480 538444 546
rect 539612 480 539640 1090
rect 540072 1018 540100 3726
rect 540428 1352 540480 1358
rect 540428 1294 540480 1300
rect 540060 1012 540112 1018
rect 540060 954 540112 960
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540440 354 540468 1294
rect 541176 1290 541204 3726
rect 542280 3726 542352 3754
rect 543428 3754 543456 4012
rect 544624 3754 544652 4012
rect 545820 3754 545848 4012
rect 546924 3754 546952 4012
rect 548120 3754 548148 4012
rect 549316 3754 549344 4012
rect 550420 3754 550448 4012
rect 551616 3754 551644 4012
rect 552720 3754 552748 4012
rect 553916 3754 553944 4012
rect 555112 3754 555140 4012
rect 556216 3754 556244 4012
rect 557412 3754 557440 4012
rect 558516 3754 558544 4012
rect 559712 3754 559740 4012
rect 543428 3726 543504 3754
rect 544624 3726 544700 3754
rect 545820 3726 545896 3754
rect 546924 3726 547000 3754
rect 548120 3726 548196 3754
rect 549316 3726 549392 3754
rect 550420 3726 550496 3754
rect 551616 3726 551692 3754
rect 552720 3726 552796 3754
rect 553916 3726 553992 3754
rect 555112 3726 555188 3754
rect 556216 3726 556292 3754
rect 557412 3726 557488 3754
rect 542280 1358 542308 3726
rect 542268 1352 542320 1358
rect 542268 1294 542320 1300
rect 541164 1284 541216 1290
rect 541164 1226 541216 1232
rect 543476 1154 543504 3726
rect 543464 1148 543516 1154
rect 543464 1090 543516 1096
rect 544672 746 544700 3726
rect 545488 1216 545540 1222
rect 545488 1158 545540 1164
rect 544660 740 544712 746
rect 544660 682 544712 688
rect 544384 604 544436 610
rect 544384 546 544436 552
rect 544396 480 544424 546
rect 545500 480 545528 1158
rect 545868 1086 545896 3726
rect 545856 1080 545908 1086
rect 545856 1022 545908 1028
rect 546684 1012 546736 1018
rect 546684 954 546736 960
rect 546696 480 546724 954
rect 540766 354 540878 480
rect 540440 326 540878 354
rect 540766 -960 540878 326
rect 541962 354 542074 480
rect 542176 468 542228 474
rect 542176 410 542228 416
rect 542188 354 542216 410
rect 541962 326 542216 354
rect 541962 -960 542074 326
rect 543158 82 543270 480
rect 542832 66 543270 82
rect 542820 60 543270 66
rect 542872 54 543270 60
rect 542820 2 542872 8
rect 543158 -960 543270 54
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 546972 66 547000 3726
rect 548168 1290 548196 3726
rect 549076 1352 549128 1358
rect 549076 1294 549128 1300
rect 547880 1284 547932 1290
rect 547880 1226 547932 1232
rect 548156 1284 548208 1290
rect 548156 1226 548208 1232
rect 547892 480 547920 1226
rect 549088 480 549116 1294
rect 549364 610 549392 3726
rect 550468 1222 550496 3726
rect 551664 1358 551692 3726
rect 551652 1352 551704 1358
rect 551652 1294 551704 1300
rect 550456 1216 550508 1222
rect 550456 1158 550508 1164
rect 552768 1154 552796 3726
rect 550272 1148 550324 1154
rect 550272 1090 550324 1096
rect 552756 1148 552808 1154
rect 552756 1090 552808 1096
rect 549352 604 549404 610
rect 549352 546 549404 552
rect 550284 480 550312 1090
rect 552664 1080 552716 1086
rect 552664 1022 552716 1028
rect 551468 740 551520 746
rect 551468 682 551520 688
rect 551480 480 551508 682
rect 552676 480 552704 1022
rect 546960 60 547012 66
rect 546960 2 547012 8
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 82 553850 480
rect 553964 270 553992 3726
rect 554964 1284 555016 1290
rect 554964 1226 555016 1232
rect 554976 480 555004 1226
rect 555160 746 555188 3726
rect 555148 740 555200 746
rect 555148 682 555200 688
rect 556264 678 556292 3726
rect 557356 1216 557408 1222
rect 557356 1158 557408 1164
rect 556252 672 556304 678
rect 556252 614 556304 620
rect 556160 604 556212 610
rect 556160 546 556212 552
rect 556172 480 556200 546
rect 557368 480 557396 1158
rect 557460 626 557488 3726
rect 558472 3726 558544 3754
rect 559668 3726 559740 3754
rect 560908 3754 560936 4012
rect 562012 3754 562040 4012
rect 563208 3754 563236 4012
rect 564312 3754 564340 4012
rect 565508 3754 565536 4012
rect 566704 3754 566732 4012
rect 560908 3726 560984 3754
rect 562012 3726 562088 3754
rect 563208 3726 563376 3754
rect 558472 1222 558500 3726
rect 558552 1352 558604 1358
rect 558552 1294 558604 1300
rect 558460 1216 558512 1222
rect 558460 1158 558512 1164
rect 557460 598 557580 626
rect 557552 542 557580 598
rect 557540 536 557592 542
rect 553952 264 554004 270
rect 553952 206 554004 212
rect 553738 66 553992 82
rect 553738 60 554004 66
rect 553738 54 553952 60
rect 553738 -960 553850 54
rect 553952 2 554004 8
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 557540 478 557592 484
rect 558564 480 558592 1294
rect 559668 1086 559696 3726
rect 560956 1358 560984 3726
rect 560944 1352 560996 1358
rect 560944 1294 560996 1300
rect 562060 1290 562088 3726
rect 562048 1284 562100 1290
rect 562048 1226 562100 1232
rect 559748 1148 559800 1154
rect 559748 1090 559800 1096
rect 559656 1080 559708 1086
rect 559656 1022 559708 1028
rect 559760 480 559788 1090
rect 562048 740 562100 746
rect 562048 682 562100 688
rect 562060 480 562088 682
rect 563152 672 563204 678
rect 563204 620 563284 626
rect 563152 614 563284 620
rect 563164 598 563284 614
rect 563348 610 563376 3726
rect 564268 3726 564340 3754
rect 565464 3726 565536 3754
rect 566660 3726 566732 3754
rect 567808 3754 567836 4012
rect 569004 3754 569032 4012
rect 570108 3754 570136 4012
rect 571304 3754 571332 4012
rect 567808 3726 567884 3754
rect 569004 3726 569080 3754
rect 570108 3726 570184 3754
rect 563256 480 563284 598
rect 563336 604 563388 610
rect 563336 546 563388 552
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560484 264 560536 270
rect 560822 218 560934 480
rect 560536 212 560934 218
rect 560484 206 560934 212
rect 560496 190 560934 206
rect 560822 -960 560934 190
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564268 270 564296 3726
rect 564624 536 564676 542
rect 564410 354 564522 480
rect 564624 478 564676 484
rect 564636 354 564664 478
rect 564410 326 564664 354
rect 565464 338 565492 3726
rect 565636 1216 565688 1222
rect 565636 1158 565688 1164
rect 565648 480 565676 1158
rect 565452 332 565504 338
rect 564256 264 564308 270
rect 564256 206 564308 212
rect 564410 -960 564522 326
rect 565452 274 565504 280
rect 565606 -960 565718 480
rect 566660 474 566688 3726
rect 567856 1154 567884 3726
rect 568028 1352 568080 1358
rect 568028 1294 568080 1300
rect 567844 1148 567896 1154
rect 567844 1090 567896 1096
rect 566832 1080 566884 1086
rect 566832 1022 566884 1028
rect 566844 480 566872 1022
rect 568040 480 568068 1294
rect 569052 1222 569080 3726
rect 570156 1290 570184 3726
rect 571260 3726 571332 3754
rect 572500 3754 572528 4012
rect 573604 3754 573632 4012
rect 574800 3754 574828 4012
rect 575918 3998 576164 4026
rect 572500 3726 572576 3754
rect 573604 3726 573680 3754
rect 574800 3726 574876 3754
rect 571260 1358 571288 3726
rect 571248 1352 571300 1358
rect 571248 1294 571300 1300
rect 569132 1284 569184 1290
rect 569132 1226 569184 1232
rect 570144 1284 570196 1290
rect 570144 1226 570196 1232
rect 569040 1216 569092 1222
rect 569040 1158 569092 1164
rect 569144 480 569172 1226
rect 570328 604 570380 610
rect 570328 546 570380 552
rect 570340 480 570368 546
rect 566648 468 566700 474
rect 566648 410 566700 416
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571340 264 571392 270
rect 571494 218 571606 480
rect 571392 212 571606 218
rect 571340 206 571606 212
rect 571352 190 571606 206
rect 571494 -960 571606 190
rect 572548 66 572576 3726
rect 572690 354 572802 480
rect 572690 338 572944 354
rect 572690 332 572956 338
rect 572690 326 572904 332
rect 572536 60 572588 66
rect 572536 2 572588 8
rect 572690 -960 572802 326
rect 572904 274 572956 280
rect 573652 134 573680 3726
rect 573732 468 573784 474
rect 573732 410 573784 416
rect 573744 354 573772 410
rect 573886 354 573998 480
rect 573744 326 573998 354
rect 573640 128 573692 134
rect 573640 70 573692 76
rect 573886 -960 573998 326
rect 574848 270 574876 3726
rect 575112 1148 575164 1154
rect 575112 1090 575164 1096
rect 575124 480 575152 1090
rect 574836 264 574888 270
rect 574836 206 574888 212
rect 575082 -960 575194 480
rect 576136 338 576164 3998
rect 578608 1352 578660 1358
rect 578608 1294 578660 1300
rect 577412 1284 577464 1290
rect 577412 1226 577464 1232
rect 576308 1216 576360 1222
rect 576308 1158 576360 1164
rect 576320 480 576348 1158
rect 577424 480 577452 1226
rect 578620 480 578648 1294
rect 576124 332 576176 338
rect 576124 274 576176 280
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 82 579886 480
rect 579632 66 579886 82
rect 579620 60 579886 66
rect 579672 54 579886 60
rect 579620 2 579672 8
rect 579774 -960 579886 54
rect 580970 82 581082 480
rect 581828 264 581880 270
rect 582166 218 582278 480
rect 581880 212 582278 218
rect 581828 206 582278 212
rect 581840 190 582278 206
rect 581184 128 581236 134
rect 580970 76 581184 82
rect 580970 70 581236 76
rect 580970 54 581224 70
rect 580970 -960 581082 54
rect 582166 -960 582278 190
rect 583362 354 583474 480
rect 583362 338 583616 354
rect 583362 332 583628 338
rect 583362 326 583576 332
rect 583362 -960 583474 326
rect 583576 274 583628 280
<< via2 >>
rect 3514 697920 3570 697976
rect 3514 697312 3570 697368
rect 579526 684664 579582 684720
rect 579618 683848 579674 683904
rect 578330 644564 578386 644600
rect 578330 644544 578332 644564
rect 578332 644544 578384 644564
rect 578384 644544 578386 644564
rect 580906 644000 580962 644056
rect 3422 436600 3478 436656
rect 3422 435986 3478 436042
rect 3422 423544 3478 423600
rect 3422 422932 3478 422988
rect 3422 410488 3478 410544
rect 3422 409878 3478 409934
rect 3422 397432 3478 397488
rect 3422 396824 3478 396880
rect 3422 384376 3478 384432
rect 3422 383648 3478 383704
rect 3422 371320 3478 371376
rect 3422 370594 3478 370650
rect 3422 358400 3478 358456
rect 3422 357540 3478 357596
rect 579526 351872 579582 351928
rect 579526 351056 579582 351112
rect 3422 345344 3478 345400
rect 3422 344364 3478 344420
rect 579618 338544 579674 338600
rect 579526 337864 579582 337920
rect 3422 332288 3478 332344
rect 3422 331310 3478 331366
rect 580170 325216 580226 325272
rect 580170 324400 580226 324456
rect 3422 319232 3478 319288
rect 3422 318256 3478 318312
rect 579618 312024 579674 312080
rect 579526 311072 579582 311128
rect 3422 306176 3478 306232
rect 3422 305080 3478 305136
rect 579618 298696 579674 298752
rect 579526 297744 579582 297800
rect 3422 293120 3478 293176
rect 3422 292026 3478 292082
rect 580170 285368 580226 285424
rect 580170 284416 580226 284472
rect 3422 280064 3478 280120
rect 3422 278972 3478 279028
rect 579618 272176 579674 272232
rect 579526 271088 579582 271144
rect 3422 267144 3478 267200
rect 3422 265918 3478 265974
rect 580906 258848 580962 258904
rect 578882 257624 578938 257680
rect 3422 254088 3478 254144
rect 3422 252742 3478 252798
rect 580170 245520 580226 245576
rect 580170 244432 580226 244488
rect 3422 241032 3478 241088
rect 3422 239688 3478 239744
rect 579618 232328 579674 232384
rect 579526 231104 579582 231160
rect 3422 227976 3478 228032
rect 3422 226634 3478 226690
rect 579618 219000 579674 219056
rect 579526 217640 579582 217696
rect 3422 214920 3478 214976
rect 3422 213458 3478 213514
rect 579618 205672 579674 205728
rect 579526 204312 579582 204368
rect 3422 201864 3478 201920
rect 3422 200404 3478 200460
rect 579618 192480 579674 192536
rect 579526 190984 579582 191040
rect 3606 188808 3662 188864
rect 3606 187350 3662 187406
rect 579618 179152 579674 179208
rect 579526 177656 579582 177712
rect 3422 175888 3478 175944
rect 3422 174174 3478 174230
rect 579618 165824 579674 165880
rect 579526 164328 579582 164384
rect 2134 162832 2190 162888
rect 2134 161064 2190 161120
rect 580906 152632 580962 152688
rect 578514 151000 578570 151056
rect 3422 149776 3478 149832
rect 3422 148066 3478 148122
rect 579618 139304 579674 139360
rect 579526 137536 579582 137592
rect 2134 136720 2190 136776
rect 2134 134952 2190 135008
rect 579618 125976 579674 126032
rect 579526 124344 579582 124400
rect 3422 123664 3478 123720
rect 3422 121836 3478 121892
rect 579618 112784 579674 112840
rect 579526 110880 579582 110936
rect 2134 110608 2190 110664
rect 2134 108840 2190 108896
rect 579618 99456 579674 99512
rect 3422 97552 3478 97608
rect 579526 97552 579582 97608
rect 3422 95728 3478 95784
rect 579618 86128 579674 86184
rect 2134 84632 2190 84688
rect 579526 84224 579582 84280
rect 2134 82592 2190 82648
rect 579618 72936 579674 72992
rect 3422 71576 3478 71632
rect 579526 70896 579582 70952
rect 3422 69498 3478 69554
rect 579618 59608 579674 59664
rect 2134 58520 2190 58576
rect 579526 57568 579582 57624
rect 2134 56480 2190 56536
rect 579986 46280 580042 46336
rect 3422 45464 3478 45520
rect 578330 44240 578386 44296
rect 3422 43268 3478 43324
rect 579618 33088 579674 33144
rect 2134 32408 2190 32464
rect 579526 30912 579582 30968
rect 2134 30232 2190 30288
rect 579618 19760 579674 19816
rect 2042 19352 2098 19408
rect 579526 17584 579582 17640
rect 2042 17176 2098 17232
rect 579618 6568 579674 6624
rect 2778 6432 2834 6488
rect 2778 4120 2834 4176
rect 579526 4120 579582 4176
<< metal3 >>
rect 3509 697978 3575 697981
rect 3509 697976 4048 697978
rect 3509 697920 3514 697976
rect 3570 697920 4048 697976
rect 3509 697918 4048 697920
rect 575920 697918 576410 697978
rect 3509 697915 3575 697918
rect 576350 697914 576410 697918
rect 576350 697854 583586 697914
rect -960 697370 480 697460
rect 3509 697370 3575 697373
rect 583526 697370 583586 697854
rect -960 697368 3575 697370
rect -960 697312 3514 697368
rect 3570 697312 3575 697368
rect -960 697310 3575 697312
rect -960 697220 480 697310
rect 3509 697307 3575 697310
rect 583342 697324 583586 697370
rect 583342 697310 584960 697324
rect 583342 697234 583402 697310
rect 583520 697234 584960 697310
rect 583342 697174 584960 697234
rect 583520 697084 584960 697174
rect 3374 684742 4048 684802
rect -960 684314 480 684404
rect 3374 684314 3434 684742
rect 579521 684722 579587 684725
rect 576350 684720 579587 684722
rect 576350 684680 579526 684720
rect 575920 684664 579526 684680
rect 579582 684664 579587 684720
rect 575920 684662 579587 684664
rect 575920 684620 576410 684662
rect 579521 684659 579587 684662
rect -960 684254 3434 684314
rect -960 684164 480 684254
rect 579613 683906 579679 683909
rect 583520 683906 584960 683996
rect 579613 683904 584960 683906
rect 579613 683848 579618 683904
rect 579674 683848 584960 683904
rect 579613 683846 584960 683848
rect 579613 683843 579679 683846
rect 583520 683756 584960 683846
rect 3374 671688 4048 671748
rect -960 671258 480 671348
rect 3374 671258 3434 671688
rect 576350 671382 583586 671394
rect 575920 671334 583586 671382
rect 575920 671322 576410 671334
rect -960 671198 3434 671258
rect -960 671108 480 671198
rect 583526 670850 583586 671334
rect 583342 670804 583586 670850
rect 583342 670790 584960 670804
rect 583342 670714 583402 670790
rect 583520 670714 584960 670790
rect 583342 670654 584960 670714
rect 583520 670564 584960 670654
rect 3374 658634 4048 658694
rect -960 658202 480 658292
rect 3374 658202 3434 658634
rect -960 658142 3434 658202
rect -960 658052 480 658142
rect 575920 657930 576410 657962
rect 575920 657902 583586 657930
rect 576350 657870 583586 657902
rect 583526 657522 583586 657870
rect 583342 657476 583586 657522
rect 583342 657462 584960 657476
rect 583342 657386 583402 657462
rect 583520 657386 584960 657462
rect 583342 657326 584960 657386
rect 583520 657236 584960 657326
rect 3374 645458 4048 645518
rect -960 645146 480 645236
rect 3374 645146 3434 645458
rect -960 645086 3434 645146
rect -960 644996 480 645086
rect 575920 644604 576410 644664
rect 576350 644602 576410 644604
rect 578325 644602 578391 644605
rect 576350 644600 578391 644602
rect 576350 644544 578330 644600
rect 578386 644544 578391 644600
rect 576350 644542 578391 644544
rect 578325 644539 578391 644542
rect 580901 644058 580967 644061
rect 583520 644058 584960 644148
rect 580901 644056 584960 644058
rect 580901 644000 580906 644056
rect 580962 644000 584960 644056
rect 580901 643998 584960 644000
rect 580901 643995 580967 643998
rect 583520 643908 584960 643998
rect 3374 632404 4048 632464
rect -960 632090 480 632180
rect 3374 632090 3434 632404
rect -960 632030 3434 632090
rect -960 631940 480 632030
rect 575920 631306 576410 631366
rect 576350 631274 576410 631306
rect 576350 631214 583586 631274
rect 583526 631002 583586 631214
rect 583342 630956 583586 631002
rect 583342 630942 584960 630956
rect 583342 630866 583402 630942
rect 583520 630866 584960 630942
rect 583342 630806 584960 630866
rect 583520 630716 584960 630806
rect 3374 619350 4048 619410
rect -960 619170 480 619260
rect 3374 619170 3434 619350
rect -960 619110 3434 619170
rect -960 619020 480 619110
rect 575920 617886 583586 617946
rect 583526 617674 583586 617886
rect 583342 617628 583586 617674
rect 583342 617614 584960 617628
rect 583342 617538 583402 617614
rect 583520 617538 584960 617614
rect 583342 617478 584960 617538
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3374 606174 4048 606234
rect 3374 606114 3434 606174
rect -960 606054 3434 606114
rect -960 605964 480 606054
rect 575920 604618 576410 604648
rect 575920 604588 576870 604618
rect 576350 604558 576870 604588
rect 576810 604482 576870 604558
rect 576810 604422 579722 604482
rect 579662 604210 579722 604422
rect 583520 604210 584960 604300
rect 579662 604150 584960 604210
rect 583520 604060 584960 604150
rect -960 593058 480 593148
rect 3374 593120 4048 593180
rect 3374 593058 3434 593120
rect -960 592998 3434 593058
rect -960 592908 480 592998
rect 575920 591290 576410 591350
rect 576350 591230 576870 591290
rect 576810 591018 576870 591230
rect 583520 591018 584960 591108
rect 576810 590958 584960 591018
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3374 580066 4048 580126
rect 3374 580002 3434 580066
rect -960 579942 3434 580002
rect -960 579852 480 579942
rect 575920 577870 576410 577930
rect 576350 577826 576410 577870
rect 576350 577766 576870 577826
rect 576810 577690 576870 577766
rect 583520 577690 584960 577780
rect 576810 577630 584960 577690
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3374 566946 4048 566950
rect -960 566890 4048 566946
rect -960 566886 3434 566890
rect -960 566796 480 566886
rect 575920 564572 576410 564632
rect 576350 564498 576410 564572
rect 576350 564438 579722 564498
rect 579662 564362 579722 564438
rect 583520 564362 584960 564452
rect 579662 564302 584960 564362
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3374 553890 4048 553896
rect -960 553836 4048 553890
rect -960 553830 3434 553836
rect -960 553740 480 553830
rect 575920 551170 576410 551212
rect 583520 551170 584960 551260
rect 575920 551152 584960 551170
rect 576350 551110 584960 551152
rect 583520 551020 584960 551110
rect -960 540834 480 540924
rect 3374 540834 4048 540842
rect -960 540782 4048 540834
rect -960 540774 3434 540782
rect -960 540684 480 540774
rect 575920 537854 576410 537914
rect 576350 537842 576410 537854
rect 583520 537842 584960 537932
rect 576350 537782 584960 537842
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect -960 527854 3434 527914
rect -960 527764 480 527854
rect 3374 527788 3434 527854
rect 3374 527728 4048 527788
rect 575920 524556 576410 524616
rect 576350 524514 576410 524556
rect 583520 524514 584960 524604
rect 576350 524454 584960 524514
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect -960 514798 3434 514858
rect -960 514708 480 514798
rect 3374 514612 3434 514798
rect 3374 514552 4048 514612
rect 583520 511322 584960 511412
rect 576350 511262 584960 511322
rect 576350 511196 576410 511262
rect 575920 511136 576410 511196
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect -960 501742 3434 501802
rect -960 501652 480 501742
rect 3374 501558 3434 501742
rect 3374 501498 4048 501558
rect 583520 497994 584960 498084
rect 576350 497934 584960 497994
rect 576350 497898 576410 497934
rect 575920 497838 576410 497898
rect 583520 497844 584960 497934
rect -960 488746 480 488836
rect -960 488686 3434 488746
rect -960 488596 480 488686
rect 3374 488504 3434 488686
rect 3374 488444 4048 488504
rect 583520 484666 584960 484756
rect 576350 484606 584960 484666
rect 576350 484600 576410 484606
rect 575920 484540 576410 484600
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect -960 475630 3434 475690
rect -960 475540 480 475630
rect 3374 475328 3434 475630
rect 3374 475268 4048 475328
rect 583520 471474 584960 471564
rect 576810 471414 584960 471474
rect 576810 471202 576870 471414
rect 583520 471324 584960 471414
rect 576350 471180 576870 471202
rect 575920 471142 576870 471180
rect 575920 471120 576410 471142
rect -960 462634 480 462724
rect -960 462574 3434 462634
rect -960 462484 480 462574
rect 3374 462274 3434 462574
rect 3374 462214 4048 462274
rect 583520 458146 584960 458236
rect 576810 458086 584960 458146
rect 576810 458010 576870 458086
rect 576350 457950 576870 458010
rect 583520 457996 584960 458086
rect 576350 457882 576410 457950
rect 575920 457822 576410 457882
rect -960 449578 480 449668
rect -960 449518 3434 449578
rect -960 449428 480 449518
rect 3374 449220 3434 449518
rect 3374 449160 4048 449220
rect 583520 444818 584960 444908
rect 576810 444758 584960 444818
rect 576810 444682 576870 444758
rect 576350 444622 576870 444682
rect 583520 444668 584960 444758
rect 576350 444584 576410 444622
rect 575920 444524 576410 444584
rect -960 436658 480 436748
rect 3417 436658 3483 436661
rect -960 436656 3483 436658
rect -960 436600 3422 436656
rect 3478 436600 3483 436656
rect -960 436598 3483 436600
rect -960 436508 480 436598
rect 3417 436595 3483 436598
rect 3417 436044 3483 436047
rect 3417 436042 4048 436044
rect 3417 435986 3422 436042
rect 3478 435986 4048 436042
rect 3417 435984 4048 435986
rect 3417 435981 3483 435984
rect 583520 431626 584960 431716
rect 583342 431566 584960 431626
rect 583342 431490 583402 431566
rect 583520 431490 584960 431566
rect 583342 431476 584960 431490
rect 583342 431430 583586 431476
rect 583526 431218 583586 431430
rect 576350 431164 583586 431218
rect 575920 431158 583586 431164
rect 575920 431104 576410 431158
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 3417 422990 3483 422993
rect 3417 422988 4048 422990
rect 3417 422932 3422 422988
rect 3478 422932 4048 422988
rect 3417 422930 4048 422932
rect 3417 422927 3483 422930
rect 583520 418298 584960 418388
rect 579662 418238 584960 418298
rect 579662 418162 579722 418238
rect 576810 418102 579722 418162
rect 583520 418148 584960 418238
rect 576810 417890 576870 418102
rect 576350 417866 576870 417890
rect 575920 417830 576870 417866
rect 575920 417806 576410 417830
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 3417 409936 3483 409939
rect 3417 409934 4048 409936
rect 3417 409878 3422 409934
rect 3478 409878 4048 409934
rect 3417 409876 4048 409878
rect 3417 409873 3483 409876
rect 583520 404970 584960 405060
rect 583342 404910 584960 404970
rect 583342 404834 583402 404910
rect 583520 404834 584960 404910
rect 583342 404820 584960 404834
rect 583342 404774 583586 404820
rect 583526 404562 583586 404774
rect 576350 404502 583586 404562
rect 576350 404446 576410 404502
rect 575920 404386 576410 404446
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 3417 396882 3483 396885
rect 3417 396880 4048 396882
rect 3417 396824 3422 396880
rect 3478 396824 4048 396880
rect 3417 396822 4048 396824
rect 3417 396819 3483 396822
rect 583520 391778 584960 391868
rect 583342 391718 584960 391778
rect 583342 391642 583402 391718
rect 583520 391642 584960 391718
rect 583342 391628 584960 391642
rect 583342 391582 583586 391628
rect 583526 391234 583586 391582
rect 576350 391174 583586 391234
rect 576350 391148 576410 391174
rect 575920 391088 576410 391148
rect -960 384434 480 384524
rect 3417 384434 3483 384437
rect -960 384432 3483 384434
rect -960 384376 3422 384432
rect 3478 384376 3483 384432
rect -960 384374 3483 384376
rect -960 384284 480 384374
rect 3417 384371 3483 384374
rect 3417 383706 3483 383709
rect 3417 383704 4048 383706
rect 3417 383648 3422 383704
rect 3478 383648 4048 383704
rect 3417 383646 4048 383648
rect 3417 383643 3483 383646
rect 583520 378450 584960 378540
rect 579662 378390 584960 378450
rect 579662 378178 579722 378390
rect 583520 378300 584960 378390
rect 579478 378118 579722 378178
rect 579478 377906 579538 378118
rect 576350 377850 579538 377906
rect 575920 377846 579538 377850
rect 575920 377790 576410 377846
rect -960 371378 480 371468
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 3417 370652 3483 370655
rect 3417 370650 4048 370652
rect 3417 370594 3422 370650
rect 3478 370594 4048 370650
rect 3417 370592 4048 370594
rect 3417 370589 3483 370592
rect 583520 365122 584960 365212
rect 583342 365062 584960 365122
rect 583342 364986 583402 365062
rect 583520 364986 584960 365062
rect 583342 364972 584960 364986
rect 583342 364926 583586 364972
rect 583526 364442 583586 364926
rect 576350 364430 583586 364442
rect 575920 364382 583586 364430
rect 575920 364370 576410 364382
rect -960 358458 480 358548
rect 3417 358458 3483 358461
rect -960 358456 3483 358458
rect -960 358400 3422 358456
rect 3478 358400 3483 358456
rect -960 358398 3483 358400
rect -960 358308 480 358398
rect 3417 358395 3483 358398
rect 3417 357598 3483 357601
rect 3417 357596 4048 357598
rect 3417 357540 3422 357596
rect 3478 357540 4048 357596
rect 3417 357538 4048 357540
rect 3417 357535 3483 357538
rect 579521 351930 579587 351933
rect 583520 351930 584960 352020
rect 579521 351928 584960 351930
rect 579521 351872 579526 351928
rect 579582 351872 584960 351928
rect 579521 351870 584960 351872
rect 579521 351867 579587 351870
rect 583520 351780 584960 351870
rect 575920 351114 576410 351132
rect 579521 351114 579587 351117
rect 575920 351112 579587 351114
rect 575920 351072 579526 351112
rect 576350 351056 579526 351072
rect 579582 351056 579587 351112
rect 576350 351054 579587 351056
rect 579521 351051 579587 351054
rect -960 345402 480 345492
rect 3417 345402 3483 345405
rect -960 345400 3483 345402
rect -960 345344 3422 345400
rect 3478 345344 3483 345400
rect -960 345342 3483 345344
rect -960 345252 480 345342
rect 3417 345339 3483 345342
rect 3417 344422 3483 344425
rect 3417 344420 4048 344422
rect 3417 344364 3422 344420
rect 3478 344364 4048 344420
rect 3417 344362 4048 344364
rect 3417 344359 3483 344362
rect 579613 338602 579679 338605
rect 583520 338602 584960 338692
rect 579613 338600 584960 338602
rect 579613 338544 579618 338600
rect 579674 338544 584960 338600
rect 579613 338542 584960 338544
rect 579613 338539 579679 338542
rect 583520 338452 584960 338542
rect 579521 337922 579587 337925
rect 576350 337920 579587 337922
rect 576350 337864 579526 337920
rect 579582 337864 579587 337920
rect 576350 337862 579587 337864
rect 576350 337834 576410 337862
rect 579521 337859 579587 337862
rect 575920 337774 576410 337834
rect -960 332346 480 332436
rect 3417 332346 3483 332349
rect -960 332344 3483 332346
rect -960 332288 3422 332344
rect 3478 332288 3483 332344
rect -960 332286 3483 332288
rect -960 332196 480 332286
rect 3417 332283 3483 332286
rect 3417 331368 3483 331371
rect 3417 331366 4048 331368
rect 3417 331310 3422 331366
rect 3478 331310 4048 331366
rect 3417 331308 4048 331310
rect 3417 331305 3483 331308
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 580165 324458 580231 324461
rect 576350 324456 580231 324458
rect 576350 324414 580170 324456
rect 575920 324400 580170 324414
rect 580226 324400 580231 324456
rect 575920 324398 580231 324400
rect 575920 324354 576410 324398
rect 580165 324395 580231 324398
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 3417 318314 3483 318317
rect 3417 318312 4048 318314
rect 3417 318256 3422 318312
rect 3478 318256 4048 318312
rect 3417 318254 4048 318256
rect 3417 318251 3483 318254
rect 579613 312082 579679 312085
rect 583520 312082 584960 312172
rect 579613 312080 584960 312082
rect 579613 312024 579618 312080
rect 579674 312024 584960 312080
rect 579613 312022 584960 312024
rect 579613 312019 579679 312022
rect 583520 311932 584960 312022
rect 579521 311130 579587 311133
rect 576350 311128 579587 311130
rect 576350 311116 579526 311128
rect 575920 311072 579526 311116
rect 579582 311072 579587 311128
rect 575920 311070 579587 311072
rect 575920 311056 576410 311070
rect 579521 311067 579587 311070
rect -960 306234 480 306324
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 3417 305138 3483 305141
rect 3417 305136 4048 305138
rect 3417 305080 3422 305136
rect 3478 305080 4048 305136
rect 3417 305078 4048 305080
rect 3417 305075 3483 305078
rect 579613 298754 579679 298757
rect 583520 298754 584960 298844
rect 579613 298752 584960 298754
rect 579613 298696 579618 298752
rect 579674 298696 584960 298752
rect 579613 298694 584960 298696
rect 579613 298691 579679 298694
rect 583520 298604 584960 298694
rect 575920 297802 576410 297818
rect 579521 297802 579587 297805
rect 575920 297800 579587 297802
rect 575920 297758 579526 297800
rect 576350 297744 579526 297758
rect 579582 297744 579587 297800
rect 576350 297742 579587 297744
rect 579521 297739 579587 297742
rect -960 293178 480 293268
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 3417 292084 3483 292087
rect 3417 292082 4048 292084
rect 3417 292026 3422 292082
rect 3478 292026 4048 292082
rect 3417 292024 4048 292026
rect 3417 292021 3483 292024
rect 580165 285426 580231 285429
rect 583520 285426 584960 285516
rect 580165 285424 584960 285426
rect 580165 285368 580170 285424
rect 580226 285368 584960 285424
rect 580165 285366 584960 285368
rect 580165 285363 580231 285366
rect 583520 285276 584960 285366
rect 580165 284474 580231 284477
rect 576350 284472 580231 284474
rect 576350 284416 580170 284472
rect 580226 284416 580231 284472
rect 576350 284414 580231 284416
rect 576350 284398 576410 284414
rect 580165 284411 580231 284414
rect 575920 284338 576410 284398
rect -960 280122 480 280212
rect 3417 280122 3483 280125
rect -960 280120 3483 280122
rect -960 280064 3422 280120
rect 3478 280064 3483 280120
rect -960 280062 3483 280064
rect -960 279972 480 280062
rect 3417 280059 3483 280062
rect 3417 279030 3483 279033
rect 3417 279028 4048 279030
rect 3417 278972 3422 279028
rect 3478 278972 4048 279028
rect 3417 278970 4048 278972
rect 3417 278967 3483 278970
rect 579613 272234 579679 272237
rect 583520 272234 584960 272324
rect 579613 272232 584960 272234
rect 579613 272176 579618 272232
rect 579674 272176 584960 272232
rect 579613 272174 584960 272176
rect 579613 272171 579679 272174
rect 583520 272084 584960 272174
rect 579521 271146 579587 271149
rect 576350 271144 579587 271146
rect 576350 271100 579526 271144
rect 575920 271088 579526 271100
rect 579582 271088 579587 271144
rect 575920 271086 579587 271088
rect 575920 271040 576410 271086
rect 579521 271083 579587 271086
rect -960 267202 480 267292
rect 3417 267202 3483 267205
rect -960 267200 3483 267202
rect -960 267144 3422 267200
rect 3478 267144 3483 267200
rect -960 267142 3483 267144
rect -960 267052 480 267142
rect 3417 267139 3483 267142
rect 3417 265976 3483 265979
rect 3417 265974 4048 265976
rect 3417 265918 3422 265974
rect 3478 265918 4048 265974
rect 3417 265916 4048 265918
rect 3417 265913 3483 265916
rect 580901 258906 580967 258909
rect 583520 258906 584960 258996
rect 580901 258904 584960 258906
rect 580901 258848 580906 258904
rect 580962 258848 584960 258904
rect 580901 258846 584960 258848
rect 580901 258843 580967 258846
rect 583520 258756 584960 258846
rect 578877 257682 578943 257685
rect 576350 257680 578943 257682
rect 575920 257624 578882 257680
rect 578938 257624 578943 257680
rect 575920 257622 578943 257624
rect 575920 257620 576410 257622
rect 578877 257619 578943 257622
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 3417 252800 3483 252803
rect 3417 252798 4048 252800
rect 3417 252742 3422 252798
rect 3478 252742 4048 252798
rect 3417 252740 4048 252742
rect 3417 252737 3483 252740
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 580165 244490 580231 244493
rect 576350 244488 580231 244490
rect 576350 244432 580170 244488
rect 580226 244432 580231 244488
rect 576350 244430 580231 244432
rect 576350 244382 576410 244430
rect 580165 244427 580231 244430
rect 575920 244322 576410 244382
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 3417 239746 3483 239749
rect 3417 239744 4048 239746
rect 3417 239688 3422 239744
rect 3478 239688 4048 239744
rect 3417 239686 4048 239688
rect 3417 239683 3483 239686
rect 579613 232386 579679 232389
rect 583520 232386 584960 232476
rect 579613 232384 584960 232386
rect 579613 232328 579618 232384
rect 579674 232328 584960 232384
rect 579613 232326 584960 232328
rect 579613 232323 579679 232326
rect 583520 232236 584960 232326
rect 579521 231162 579587 231165
rect 576350 231160 579587 231162
rect 576350 231104 579526 231160
rect 579582 231104 579587 231160
rect 576350 231102 579587 231104
rect 576350 231084 576410 231102
rect 579521 231099 579587 231102
rect 575920 231024 576410 231084
rect -960 228034 480 228124
rect 3417 228034 3483 228037
rect -960 228032 3483 228034
rect -960 227976 3422 228032
rect 3478 227976 3483 228032
rect -960 227974 3483 227976
rect -960 227884 480 227974
rect 3417 227971 3483 227974
rect 3417 226692 3483 226695
rect 3417 226690 4048 226692
rect 3417 226634 3422 226690
rect 3478 226634 4048 226690
rect 3417 226632 4048 226634
rect 3417 226629 3483 226632
rect 579613 219058 579679 219061
rect 583520 219058 584960 219148
rect 579613 219056 584960 219058
rect 579613 219000 579618 219056
rect 579674 219000 584960 219056
rect 579613 218998 584960 219000
rect 579613 218995 579679 218998
rect 583520 218908 584960 218998
rect 579521 217698 579587 217701
rect 576350 217696 579587 217698
rect 576350 217664 579526 217696
rect 575920 217640 579526 217664
rect 579582 217640 579587 217696
rect 575920 217638 579587 217640
rect 575920 217604 576410 217638
rect 579521 217635 579587 217638
rect -960 214978 480 215068
rect 3417 214978 3483 214981
rect -960 214976 3483 214978
rect -960 214920 3422 214976
rect 3478 214920 3483 214976
rect -960 214918 3483 214920
rect -960 214828 480 214918
rect 3417 214915 3483 214918
rect 3417 213516 3483 213519
rect 3417 213514 4048 213516
rect 3417 213458 3422 213514
rect 3478 213458 4048 213514
rect 3417 213456 4048 213458
rect 3417 213453 3483 213456
rect 579613 205730 579679 205733
rect 583520 205730 584960 205820
rect 579613 205728 584960 205730
rect 579613 205672 579618 205728
rect 579674 205672 584960 205728
rect 579613 205670 584960 205672
rect 579613 205667 579679 205670
rect 583520 205580 584960 205670
rect 579521 204370 579587 204373
rect 576350 204368 579587 204370
rect 576350 204366 579526 204368
rect 575920 204312 579526 204366
rect 579582 204312 579587 204368
rect 575920 204310 579587 204312
rect 575920 204306 576410 204310
rect 579521 204307 579587 204310
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 3417 200462 3483 200465
rect 3417 200460 4048 200462
rect 3417 200404 3422 200460
rect 3478 200404 4048 200460
rect 3417 200402 4048 200404
rect 3417 200399 3483 200402
rect 579613 192538 579679 192541
rect 583520 192538 584960 192628
rect 579613 192536 584960 192538
rect 579613 192480 579618 192536
rect 579674 192480 584960 192536
rect 579613 192478 584960 192480
rect 579613 192475 579679 192478
rect 583520 192388 584960 192478
rect 575920 191042 576410 191068
rect 579521 191042 579587 191045
rect 575920 191040 579587 191042
rect 575920 191008 579526 191040
rect 576350 190984 579526 191008
rect 579582 190984 579587 191040
rect 576350 190982 579587 190984
rect 579521 190979 579587 190982
rect -960 188866 480 188956
rect 3601 188866 3667 188869
rect -960 188864 3667 188866
rect -960 188808 3606 188864
rect 3662 188808 3667 188864
rect -960 188806 3667 188808
rect -960 188716 480 188806
rect 3601 188803 3667 188806
rect 3601 187408 3667 187411
rect 3601 187406 4048 187408
rect 3601 187350 3606 187406
rect 3662 187350 4048 187406
rect 3601 187348 4048 187350
rect 3601 187345 3667 187348
rect 579613 179210 579679 179213
rect 583520 179210 584960 179300
rect 579613 179208 584960 179210
rect 579613 179152 579618 179208
rect 579674 179152 584960 179208
rect 579613 179150 584960 179152
rect 579613 179147 579679 179150
rect 583520 179060 584960 179150
rect 579521 177714 579587 177717
rect 576350 177712 579587 177714
rect 576350 177656 579526 177712
rect 579582 177656 579587 177712
rect 576350 177654 579587 177656
rect 576350 177648 576410 177654
rect 579521 177651 579587 177654
rect 575920 177588 576410 177648
rect -960 175946 480 176036
rect 3417 175946 3483 175949
rect -960 175944 3483 175946
rect -960 175888 3422 175944
rect 3478 175888 3483 175944
rect -960 175886 3483 175888
rect -960 175796 480 175886
rect 3417 175883 3483 175886
rect 3417 174232 3483 174235
rect 3417 174230 4048 174232
rect 3417 174174 3422 174230
rect 3478 174174 4048 174230
rect 3417 174172 4048 174174
rect 3417 174169 3483 174172
rect 579613 165882 579679 165885
rect 583520 165882 584960 165972
rect 579613 165880 584960 165882
rect 579613 165824 579618 165880
rect 579674 165824 584960 165880
rect 579613 165822 584960 165824
rect 579613 165819 579679 165822
rect 583520 165732 584960 165822
rect 579521 164386 579587 164389
rect 576350 164384 579587 164386
rect 576350 164350 579526 164384
rect 575920 164328 579526 164350
rect 579582 164328 579587 164384
rect 575920 164326 579587 164328
rect 575920 164290 576410 164326
rect 579521 164323 579587 164326
rect -960 162890 480 162980
rect 2129 162890 2195 162893
rect -960 162888 2195 162890
rect -960 162832 2134 162888
rect 2190 162832 2195 162888
rect -960 162830 2195 162832
rect -960 162740 480 162830
rect 2129 162827 2195 162830
rect 2129 161122 2195 161125
rect 3374 161122 4048 161178
rect 2129 161120 4048 161122
rect 2129 161064 2134 161120
rect 2190 161118 4048 161120
rect 2190 161064 3434 161118
rect 2129 161062 3434 161064
rect 2129 161059 2195 161062
rect 580901 152690 580967 152693
rect 583520 152690 584960 152780
rect 580901 152688 584960 152690
rect 580901 152632 580906 152688
rect 580962 152632 584960 152688
rect 580901 152630 584960 152632
rect 580901 152627 580967 152630
rect 583520 152540 584960 152630
rect 578509 151058 578575 151061
rect 576350 151056 578575 151058
rect 576350 151052 578514 151056
rect 575920 151000 578514 151052
rect 578570 151000 578575 151056
rect 575920 150998 578575 151000
rect 575920 150992 576410 150998
rect 578509 150995 578575 150998
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 3417 148124 3483 148127
rect 3417 148122 4048 148124
rect 3417 148066 3422 148122
rect 3478 148066 4048 148122
rect 3417 148064 4048 148066
rect 3417 148061 3483 148064
rect 579613 139362 579679 139365
rect 583520 139362 584960 139452
rect 579613 139360 584960 139362
rect 579613 139304 579618 139360
rect 579674 139304 584960 139360
rect 579613 139302 584960 139304
rect 579613 139299 579679 139302
rect 583520 139212 584960 139302
rect 575920 137594 576410 137632
rect 579521 137594 579587 137597
rect 575920 137592 579587 137594
rect 575920 137572 579526 137592
rect 576350 137536 579526 137572
rect 579582 137536 579587 137592
rect 576350 137534 579587 137536
rect 579521 137531 579587 137534
rect -960 136778 480 136868
rect 2129 136778 2195 136781
rect -960 136776 2195 136778
rect -960 136720 2134 136776
rect 2190 136720 2195 136776
rect -960 136718 2195 136720
rect -960 136628 480 136718
rect 2129 136715 2195 136718
rect 2129 135010 2195 135013
rect 3374 135010 4048 135070
rect 2129 135008 3434 135010
rect 2129 134952 2134 135008
rect 2190 134952 3434 135008
rect 2129 134950 3434 134952
rect 2129 134947 2195 134950
rect 579613 126034 579679 126037
rect 583520 126034 584960 126124
rect 579613 126032 584960 126034
rect 579613 125976 579618 126032
rect 579674 125976 584960 126032
rect 579613 125974 584960 125976
rect 579613 125971 579679 125974
rect 583520 125884 584960 125974
rect 579521 124402 579587 124405
rect 576350 124400 579587 124402
rect 576350 124344 579526 124400
rect 579582 124344 579587 124400
rect 576350 124342 579587 124344
rect 576350 124334 576410 124342
rect 579521 124339 579587 124342
rect 575920 124274 576410 124334
rect -960 123722 480 123812
rect 3417 123722 3483 123725
rect -960 123720 3483 123722
rect -960 123664 3422 123720
rect 3478 123664 3483 123720
rect -960 123662 3483 123664
rect -960 123572 480 123662
rect 3417 123659 3483 123662
rect 3417 121894 3483 121897
rect 3417 121892 4048 121894
rect 3417 121836 3422 121892
rect 3478 121836 4048 121892
rect 3417 121834 4048 121836
rect 3417 121831 3483 121834
rect 579613 112842 579679 112845
rect 583520 112842 584960 112932
rect 579613 112840 584960 112842
rect 579613 112784 579618 112840
rect 579674 112784 584960 112840
rect 579613 112782 584960 112784
rect 579613 112779 579679 112782
rect 583520 112692 584960 112782
rect 579521 110938 579587 110941
rect 576350 110936 579587 110938
rect 576350 110914 579526 110936
rect 575920 110880 579526 110914
rect 579582 110880 579587 110936
rect 575920 110878 579587 110880
rect 575920 110854 576410 110878
rect 579521 110875 579587 110878
rect -960 110666 480 110756
rect 2129 110666 2195 110669
rect -960 110664 2195 110666
rect -960 110608 2134 110664
rect 2190 110608 2195 110664
rect -960 110606 2195 110608
rect -960 110516 480 110606
rect 2129 110603 2195 110606
rect 2129 108898 2195 108901
rect 2129 108896 3434 108898
rect 2129 108840 2134 108896
rect 2190 108840 3434 108896
rect 2129 108838 4048 108840
rect 2129 108835 2195 108838
rect 3374 108780 4048 108838
rect 579613 99514 579679 99517
rect 583520 99514 584960 99604
rect 579613 99512 584960 99514
rect 579613 99456 579618 99512
rect 579674 99456 584960 99512
rect 579613 99454 584960 99456
rect 579613 99451 579679 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect 575920 97610 576410 97616
rect 579521 97610 579587 97613
rect 575920 97608 579587 97610
rect 575920 97556 579526 97608
rect -960 97550 3483 97552
rect 576350 97552 579526 97556
rect 579582 97552 579587 97608
rect 576350 97550 579587 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 579521 97547 579587 97550
rect 3417 95786 3483 95789
rect 3417 95784 4048 95786
rect 3417 95728 3422 95784
rect 3478 95728 4048 95784
rect 3417 95726 4048 95728
rect 3417 95723 3483 95726
rect 579613 86186 579679 86189
rect 583520 86186 584960 86276
rect 579613 86184 584960 86186
rect 579613 86128 579618 86184
rect 579674 86128 584960 86184
rect 579613 86126 584960 86128
rect 579613 86123 579679 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 2129 84690 2195 84693
rect -960 84688 2195 84690
rect -960 84632 2134 84688
rect 2190 84632 2195 84688
rect -960 84630 2195 84632
rect -960 84540 480 84630
rect 2129 84627 2195 84630
rect 575920 84282 576410 84318
rect 579521 84282 579587 84285
rect 575920 84280 579587 84282
rect 575920 84258 579526 84280
rect 576350 84224 579526 84258
rect 579582 84224 579587 84280
rect 576350 84222 579587 84224
rect 579521 84219 579587 84222
rect 2129 82650 2195 82653
rect 2129 82648 3434 82650
rect 2129 82592 2134 82648
rect 2190 82610 3434 82648
rect 2190 82592 4048 82610
rect 2129 82590 4048 82592
rect 2129 82587 2195 82590
rect 3374 82550 4048 82590
rect 579613 72994 579679 72997
rect 583520 72994 584960 73084
rect 579613 72992 584960 72994
rect 579613 72936 579618 72992
rect 579674 72936 584960 72992
rect 579613 72934 584960 72936
rect 579613 72931 579679 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 579521 70954 579587 70957
rect 576350 70952 579587 70954
rect 576350 70898 579526 70952
rect 575920 70896 579526 70898
rect 579582 70896 579587 70952
rect 575920 70894 579587 70896
rect 575920 70838 576410 70894
rect 579521 70891 579587 70894
rect 3417 69556 3483 69559
rect 3417 69554 4048 69556
rect 3417 69498 3422 69554
rect 3478 69498 4048 69554
rect 3417 69496 4048 69498
rect 3417 69493 3483 69496
rect 579613 59666 579679 59669
rect 583520 59666 584960 59756
rect 579613 59664 584960 59666
rect 579613 59608 579618 59664
rect 579674 59608 584960 59664
rect 579613 59606 584960 59608
rect 579613 59603 579679 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 2129 58578 2195 58581
rect -960 58576 2195 58578
rect -960 58520 2134 58576
rect 2190 58520 2195 58576
rect -960 58518 2195 58520
rect -960 58428 480 58518
rect 2129 58515 2195 58518
rect 579521 57626 579587 57629
rect 576350 57624 579587 57626
rect 576350 57600 579526 57624
rect 575920 57568 579526 57600
rect 579582 57568 579587 57624
rect 575920 57566 579587 57568
rect 575920 57540 576410 57566
rect 579521 57563 579587 57566
rect 2129 56538 2195 56541
rect 2129 56536 3434 56538
rect 2129 56480 2134 56536
rect 2190 56502 3434 56536
rect 2190 56480 4048 56502
rect 2129 56478 4048 56480
rect 2129 56475 2195 56478
rect 3374 56442 4048 56478
rect 579981 46338 580047 46341
rect 583520 46338 584960 46428
rect 579981 46336 584960 46338
rect 579981 46280 579986 46336
rect 580042 46280 584960 46336
rect 579981 46278 584960 46280
rect 579981 46275 580047 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 575920 44298 576410 44302
rect 578325 44298 578391 44301
rect 575920 44296 578391 44298
rect 575920 44242 578330 44296
rect 576350 44240 578330 44242
rect 578386 44240 578391 44296
rect 576350 44238 578391 44240
rect 578325 44235 578391 44238
rect 3417 43326 3483 43329
rect 3417 43324 4048 43326
rect 3417 43268 3422 43324
rect 3478 43268 4048 43324
rect 3417 43266 4048 43268
rect 3417 43263 3483 43266
rect 579613 33146 579679 33149
rect 583520 33146 584960 33236
rect 579613 33144 584960 33146
rect 579613 33088 579618 33144
rect 579674 33088 584960 33144
rect 579613 33086 584960 33088
rect 579613 33083 579679 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2129 32466 2195 32469
rect -960 32464 2195 32466
rect -960 32408 2134 32464
rect 2190 32408 2195 32464
rect -960 32406 2195 32408
rect -960 32316 480 32406
rect 2129 32403 2195 32406
rect 579521 30970 579587 30973
rect 576350 30968 579587 30970
rect 576350 30912 579526 30968
rect 579582 30912 579587 30968
rect 576350 30910 579587 30912
rect 576350 30882 576410 30910
rect 579521 30907 579587 30910
rect 575920 30822 576410 30882
rect 2129 30290 2195 30293
rect 2129 30288 3434 30290
rect 2129 30232 2134 30288
rect 2190 30272 3434 30288
rect 2190 30232 4048 30272
rect 2129 30230 4048 30232
rect 2129 30227 2195 30230
rect 3374 30212 4048 30230
rect 579613 19818 579679 19821
rect 583520 19818 584960 19908
rect 579613 19816 584960 19818
rect 579613 19760 579618 19816
rect 579674 19760 584960 19816
rect 579613 19758 584960 19760
rect 579613 19755 579679 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 2037 19410 2103 19413
rect -960 19408 2103 19410
rect -960 19352 2042 19408
rect 2098 19352 2103 19408
rect -960 19350 2103 19352
rect -960 19260 480 19350
rect 2037 19347 2103 19350
rect 579521 17642 579587 17645
rect 576350 17640 579587 17642
rect 576350 17584 579526 17640
rect 579582 17584 579587 17640
rect 575920 17582 579587 17584
rect 575920 17524 576410 17582
rect 579521 17579 579587 17582
rect 2037 17234 2103 17237
rect 2037 17232 3434 17234
rect 2037 17176 2042 17232
rect 2098 17218 3434 17232
rect 2098 17176 4048 17218
rect 2037 17174 4048 17176
rect 2037 17171 2103 17174
rect 3374 17158 4048 17174
rect 579613 6626 579679 6629
rect 583520 6626 584960 6716
rect 579613 6624 584960 6626
rect -960 6490 480 6580
rect 579613 6568 579618 6624
rect 579674 6568 584960 6624
rect 579613 6566 584960 6568
rect 579613 6563 579679 6566
rect 2773 6490 2839 6493
rect -960 6488 2839 6490
rect -960 6432 2778 6488
rect 2834 6432 2839 6488
rect 583520 6476 584960 6566
rect -960 6430 2839 6432
rect -960 6340 480 6430
rect 2773 6427 2839 6430
rect 2773 4178 2839 4181
rect 579521 4178 579587 4181
rect 2773 4176 3802 4178
rect 2773 4120 2778 4176
rect 2834 4164 3802 4176
rect 576166 4176 579587 4178
rect 576166 4164 579526 4176
rect 2834 4120 4048 4164
rect 2773 4118 4048 4120
rect 2773 4115 2839 4118
rect 3742 4104 4048 4118
rect 575920 4120 579526 4164
rect 579582 4120 579587 4176
rect 575920 4118 579587 4120
rect 575920 4104 576226 4118
rect 579521 4115 579587 4118
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 674814 -8106 711002
rect -8726 674578 -8694 674814
rect -8458 674578 -8374 674814
rect -8138 674578 -8106 674814
rect -8726 674494 -8106 674578
rect -8726 674258 -8694 674494
rect -8458 674258 -8374 674494
rect -8138 674258 -8106 674494
rect -8726 634814 -8106 674258
rect -8726 634578 -8694 634814
rect -8458 634578 -8374 634814
rect -8138 634578 -8106 634814
rect -8726 634494 -8106 634578
rect -8726 634258 -8694 634494
rect -8458 634258 -8374 634494
rect -8138 634258 -8106 634494
rect -8726 594814 -8106 634258
rect -8726 594578 -8694 594814
rect -8458 594578 -8374 594814
rect -8138 594578 -8106 594814
rect -8726 594494 -8106 594578
rect -8726 594258 -8694 594494
rect -8458 594258 -8374 594494
rect -8138 594258 -8106 594494
rect -8726 554814 -8106 594258
rect -8726 554578 -8694 554814
rect -8458 554578 -8374 554814
rect -8138 554578 -8106 554814
rect -8726 554494 -8106 554578
rect -8726 554258 -8694 554494
rect -8458 554258 -8374 554494
rect -8138 554258 -8106 554494
rect -8726 514814 -8106 554258
rect -8726 514578 -8694 514814
rect -8458 514578 -8374 514814
rect -8138 514578 -8106 514814
rect -8726 514494 -8106 514578
rect -8726 514258 -8694 514494
rect -8458 514258 -8374 514494
rect -8138 514258 -8106 514494
rect -8726 474814 -8106 514258
rect -8726 474578 -8694 474814
rect -8458 474578 -8374 474814
rect -8138 474578 -8106 474814
rect -8726 474494 -8106 474578
rect -8726 474258 -8694 474494
rect -8458 474258 -8374 474494
rect -8138 474258 -8106 474494
rect -8726 434814 -8106 474258
rect -8726 434578 -8694 434814
rect -8458 434578 -8374 434814
rect -8138 434578 -8106 434814
rect -8726 434494 -8106 434578
rect -8726 434258 -8694 434494
rect -8458 434258 -8374 434494
rect -8138 434258 -8106 434494
rect -8726 394814 -8106 434258
rect -8726 394578 -8694 394814
rect -8458 394578 -8374 394814
rect -8138 394578 -8106 394814
rect -8726 394494 -8106 394578
rect -8726 394258 -8694 394494
rect -8458 394258 -8374 394494
rect -8138 394258 -8106 394494
rect -8726 354814 -8106 394258
rect -8726 354578 -8694 354814
rect -8458 354578 -8374 354814
rect -8138 354578 -8106 354814
rect -8726 354494 -8106 354578
rect -8726 354258 -8694 354494
rect -8458 354258 -8374 354494
rect -8138 354258 -8106 354494
rect -8726 314814 -8106 354258
rect -8726 314578 -8694 314814
rect -8458 314578 -8374 314814
rect -8138 314578 -8106 314814
rect -8726 314494 -8106 314578
rect -8726 314258 -8694 314494
rect -8458 314258 -8374 314494
rect -8138 314258 -8106 314494
rect -8726 274814 -8106 314258
rect -8726 274578 -8694 274814
rect -8458 274578 -8374 274814
rect -8138 274578 -8106 274814
rect -8726 274494 -8106 274578
rect -8726 274258 -8694 274494
rect -8458 274258 -8374 274494
rect -8138 274258 -8106 274494
rect -8726 234814 -8106 274258
rect -8726 234578 -8694 234814
rect -8458 234578 -8374 234814
rect -8138 234578 -8106 234814
rect -8726 234494 -8106 234578
rect -8726 234258 -8694 234494
rect -8458 234258 -8374 234494
rect -8138 234258 -8106 234494
rect -8726 194814 -8106 234258
rect -8726 194578 -8694 194814
rect -8458 194578 -8374 194814
rect -8138 194578 -8106 194814
rect -8726 194494 -8106 194578
rect -8726 194258 -8694 194494
rect -8458 194258 -8374 194494
rect -8138 194258 -8106 194494
rect -8726 154814 -8106 194258
rect -8726 154578 -8694 154814
rect -8458 154578 -8374 154814
rect -8138 154578 -8106 154814
rect -8726 154494 -8106 154578
rect -8726 154258 -8694 154494
rect -8458 154258 -8374 154494
rect -8138 154258 -8106 154494
rect -8726 114814 -8106 154258
rect -8726 114578 -8694 114814
rect -8458 114578 -8374 114814
rect -8138 114578 -8106 114814
rect -8726 114494 -8106 114578
rect -8726 114258 -8694 114494
rect -8458 114258 -8374 114494
rect -8138 114258 -8106 114494
rect -8726 74814 -8106 114258
rect -8726 74578 -8694 74814
rect -8458 74578 -8374 74814
rect -8138 74578 -8106 74814
rect -8726 74494 -8106 74578
rect -8726 74258 -8694 74494
rect -8458 74258 -8374 74494
rect -8138 74258 -8106 74494
rect -8726 34814 -8106 74258
rect -8726 34578 -8694 34814
rect -8458 34578 -8374 34814
rect -8138 34578 -8106 34814
rect -8726 34494 -8106 34578
rect -8726 34258 -8694 34494
rect -8458 34258 -8374 34494
rect -8138 34258 -8106 34494
rect -8726 -7066 -8106 34258
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 694814 -7146 710042
rect 13154 710598 13774 711590
rect 13154 710362 13186 710598
rect 13422 710362 13506 710598
rect 13742 710362 13774 710598
rect 13154 710278 13774 710362
rect 13154 710042 13186 710278
rect 13422 710042 13506 710278
rect 13742 710042 13774 710278
rect -7766 694578 -7734 694814
rect -7498 694578 -7414 694814
rect -7178 694578 -7146 694814
rect -7766 694494 -7146 694578
rect -7766 694258 -7734 694494
rect -7498 694258 -7414 694494
rect -7178 694258 -7146 694494
rect -7766 654814 -7146 694258
rect -7766 654578 -7734 654814
rect -7498 654578 -7414 654814
rect -7178 654578 -7146 654814
rect -7766 654494 -7146 654578
rect -7766 654258 -7734 654494
rect -7498 654258 -7414 654494
rect -7178 654258 -7146 654494
rect -7766 614814 -7146 654258
rect -7766 614578 -7734 614814
rect -7498 614578 -7414 614814
rect -7178 614578 -7146 614814
rect -7766 614494 -7146 614578
rect -7766 614258 -7734 614494
rect -7498 614258 -7414 614494
rect -7178 614258 -7146 614494
rect -7766 574814 -7146 614258
rect -7766 574578 -7734 574814
rect -7498 574578 -7414 574814
rect -7178 574578 -7146 574814
rect -7766 574494 -7146 574578
rect -7766 574258 -7734 574494
rect -7498 574258 -7414 574494
rect -7178 574258 -7146 574494
rect -7766 534814 -7146 574258
rect -7766 534578 -7734 534814
rect -7498 534578 -7414 534814
rect -7178 534578 -7146 534814
rect -7766 534494 -7146 534578
rect -7766 534258 -7734 534494
rect -7498 534258 -7414 534494
rect -7178 534258 -7146 534494
rect -7766 494814 -7146 534258
rect -7766 494578 -7734 494814
rect -7498 494578 -7414 494814
rect -7178 494578 -7146 494814
rect -7766 494494 -7146 494578
rect -7766 494258 -7734 494494
rect -7498 494258 -7414 494494
rect -7178 494258 -7146 494494
rect -7766 454814 -7146 494258
rect -7766 454578 -7734 454814
rect -7498 454578 -7414 454814
rect -7178 454578 -7146 454814
rect -7766 454494 -7146 454578
rect -7766 454258 -7734 454494
rect -7498 454258 -7414 454494
rect -7178 454258 -7146 454494
rect -7766 414814 -7146 454258
rect -7766 414578 -7734 414814
rect -7498 414578 -7414 414814
rect -7178 414578 -7146 414814
rect -7766 414494 -7146 414578
rect -7766 414258 -7734 414494
rect -7498 414258 -7414 414494
rect -7178 414258 -7146 414494
rect -7766 374814 -7146 414258
rect -7766 374578 -7734 374814
rect -7498 374578 -7414 374814
rect -7178 374578 -7146 374814
rect -7766 374494 -7146 374578
rect -7766 374258 -7734 374494
rect -7498 374258 -7414 374494
rect -7178 374258 -7146 374494
rect -7766 334814 -7146 374258
rect -7766 334578 -7734 334814
rect -7498 334578 -7414 334814
rect -7178 334578 -7146 334814
rect -7766 334494 -7146 334578
rect -7766 334258 -7734 334494
rect -7498 334258 -7414 334494
rect -7178 334258 -7146 334494
rect -7766 294814 -7146 334258
rect -7766 294578 -7734 294814
rect -7498 294578 -7414 294814
rect -7178 294578 -7146 294814
rect -7766 294494 -7146 294578
rect -7766 294258 -7734 294494
rect -7498 294258 -7414 294494
rect -7178 294258 -7146 294494
rect -7766 254814 -7146 294258
rect -7766 254578 -7734 254814
rect -7498 254578 -7414 254814
rect -7178 254578 -7146 254814
rect -7766 254494 -7146 254578
rect -7766 254258 -7734 254494
rect -7498 254258 -7414 254494
rect -7178 254258 -7146 254494
rect -7766 214814 -7146 254258
rect -7766 214578 -7734 214814
rect -7498 214578 -7414 214814
rect -7178 214578 -7146 214814
rect -7766 214494 -7146 214578
rect -7766 214258 -7734 214494
rect -7498 214258 -7414 214494
rect -7178 214258 -7146 214494
rect -7766 174814 -7146 214258
rect -7766 174578 -7734 174814
rect -7498 174578 -7414 174814
rect -7178 174578 -7146 174814
rect -7766 174494 -7146 174578
rect -7766 174258 -7734 174494
rect -7498 174258 -7414 174494
rect -7178 174258 -7146 174494
rect -7766 134814 -7146 174258
rect -7766 134578 -7734 134814
rect -7498 134578 -7414 134814
rect -7178 134578 -7146 134814
rect -7766 134494 -7146 134578
rect -7766 134258 -7734 134494
rect -7498 134258 -7414 134494
rect -7178 134258 -7146 134494
rect -7766 94814 -7146 134258
rect -7766 94578 -7734 94814
rect -7498 94578 -7414 94814
rect -7178 94578 -7146 94814
rect -7766 94494 -7146 94578
rect -7766 94258 -7734 94494
rect -7498 94258 -7414 94494
rect -7178 94258 -7146 94494
rect -7766 54814 -7146 94258
rect -7766 54578 -7734 54814
rect -7498 54578 -7414 54814
rect -7178 54578 -7146 54814
rect -7766 54494 -7146 54578
rect -7766 54258 -7734 54494
rect -7498 54258 -7414 54494
rect -7178 54258 -7146 54494
rect -7766 14814 -7146 54258
rect -7766 14578 -7734 14814
rect -7498 14578 -7414 14814
rect -7178 14578 -7146 14814
rect -7766 14494 -7146 14578
rect -7766 14258 -7734 14494
rect -7498 14258 -7414 14494
rect -7178 14258 -7146 14494
rect -7766 -6106 -7146 14258
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 671094 -6186 709082
rect -6806 670858 -6774 671094
rect -6538 670858 -6454 671094
rect -6218 670858 -6186 671094
rect -6806 670774 -6186 670858
rect -6806 670538 -6774 670774
rect -6538 670538 -6454 670774
rect -6218 670538 -6186 670774
rect -6806 631094 -6186 670538
rect -6806 630858 -6774 631094
rect -6538 630858 -6454 631094
rect -6218 630858 -6186 631094
rect -6806 630774 -6186 630858
rect -6806 630538 -6774 630774
rect -6538 630538 -6454 630774
rect -6218 630538 -6186 630774
rect -6806 591094 -6186 630538
rect -6806 590858 -6774 591094
rect -6538 590858 -6454 591094
rect -6218 590858 -6186 591094
rect -6806 590774 -6186 590858
rect -6806 590538 -6774 590774
rect -6538 590538 -6454 590774
rect -6218 590538 -6186 590774
rect -6806 551094 -6186 590538
rect -6806 550858 -6774 551094
rect -6538 550858 -6454 551094
rect -6218 550858 -6186 551094
rect -6806 550774 -6186 550858
rect -6806 550538 -6774 550774
rect -6538 550538 -6454 550774
rect -6218 550538 -6186 550774
rect -6806 511094 -6186 550538
rect -6806 510858 -6774 511094
rect -6538 510858 -6454 511094
rect -6218 510858 -6186 511094
rect -6806 510774 -6186 510858
rect -6806 510538 -6774 510774
rect -6538 510538 -6454 510774
rect -6218 510538 -6186 510774
rect -6806 471094 -6186 510538
rect -6806 470858 -6774 471094
rect -6538 470858 -6454 471094
rect -6218 470858 -6186 471094
rect -6806 470774 -6186 470858
rect -6806 470538 -6774 470774
rect -6538 470538 -6454 470774
rect -6218 470538 -6186 470774
rect -6806 431094 -6186 470538
rect -6806 430858 -6774 431094
rect -6538 430858 -6454 431094
rect -6218 430858 -6186 431094
rect -6806 430774 -6186 430858
rect -6806 430538 -6774 430774
rect -6538 430538 -6454 430774
rect -6218 430538 -6186 430774
rect -6806 391094 -6186 430538
rect -6806 390858 -6774 391094
rect -6538 390858 -6454 391094
rect -6218 390858 -6186 391094
rect -6806 390774 -6186 390858
rect -6806 390538 -6774 390774
rect -6538 390538 -6454 390774
rect -6218 390538 -6186 390774
rect -6806 351094 -6186 390538
rect -6806 350858 -6774 351094
rect -6538 350858 -6454 351094
rect -6218 350858 -6186 351094
rect -6806 350774 -6186 350858
rect -6806 350538 -6774 350774
rect -6538 350538 -6454 350774
rect -6218 350538 -6186 350774
rect -6806 311094 -6186 350538
rect -6806 310858 -6774 311094
rect -6538 310858 -6454 311094
rect -6218 310858 -6186 311094
rect -6806 310774 -6186 310858
rect -6806 310538 -6774 310774
rect -6538 310538 -6454 310774
rect -6218 310538 -6186 310774
rect -6806 271094 -6186 310538
rect -6806 270858 -6774 271094
rect -6538 270858 -6454 271094
rect -6218 270858 -6186 271094
rect -6806 270774 -6186 270858
rect -6806 270538 -6774 270774
rect -6538 270538 -6454 270774
rect -6218 270538 -6186 270774
rect -6806 231094 -6186 270538
rect -6806 230858 -6774 231094
rect -6538 230858 -6454 231094
rect -6218 230858 -6186 231094
rect -6806 230774 -6186 230858
rect -6806 230538 -6774 230774
rect -6538 230538 -6454 230774
rect -6218 230538 -6186 230774
rect -6806 191094 -6186 230538
rect -6806 190858 -6774 191094
rect -6538 190858 -6454 191094
rect -6218 190858 -6186 191094
rect -6806 190774 -6186 190858
rect -6806 190538 -6774 190774
rect -6538 190538 -6454 190774
rect -6218 190538 -6186 190774
rect -6806 151094 -6186 190538
rect -6806 150858 -6774 151094
rect -6538 150858 -6454 151094
rect -6218 150858 -6186 151094
rect -6806 150774 -6186 150858
rect -6806 150538 -6774 150774
rect -6538 150538 -6454 150774
rect -6218 150538 -6186 150774
rect -6806 111094 -6186 150538
rect -6806 110858 -6774 111094
rect -6538 110858 -6454 111094
rect -6218 110858 -6186 111094
rect -6806 110774 -6186 110858
rect -6806 110538 -6774 110774
rect -6538 110538 -6454 110774
rect -6218 110538 -6186 110774
rect -6806 71094 -6186 110538
rect -6806 70858 -6774 71094
rect -6538 70858 -6454 71094
rect -6218 70858 -6186 71094
rect -6806 70774 -6186 70858
rect -6806 70538 -6774 70774
rect -6538 70538 -6454 70774
rect -6218 70538 -6186 70774
rect -6806 31094 -6186 70538
rect -6806 30858 -6774 31094
rect -6538 30858 -6454 31094
rect -6218 30858 -6186 31094
rect -6806 30774 -6186 30858
rect -6806 30538 -6774 30774
rect -6538 30538 -6454 30774
rect -6218 30538 -6186 30774
rect -6806 -5146 -6186 30538
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 691094 -5226 708122
rect 9434 708678 10054 709670
rect 9434 708442 9466 708678
rect 9702 708442 9786 708678
rect 10022 708442 10054 708678
rect 9434 708358 10054 708442
rect 9434 708122 9466 708358
rect 9702 708122 9786 708358
rect 10022 708122 10054 708358
rect -5846 690858 -5814 691094
rect -5578 690858 -5494 691094
rect -5258 690858 -5226 691094
rect -5846 690774 -5226 690858
rect -5846 690538 -5814 690774
rect -5578 690538 -5494 690774
rect -5258 690538 -5226 690774
rect -5846 651094 -5226 690538
rect -5846 650858 -5814 651094
rect -5578 650858 -5494 651094
rect -5258 650858 -5226 651094
rect -5846 650774 -5226 650858
rect -5846 650538 -5814 650774
rect -5578 650538 -5494 650774
rect -5258 650538 -5226 650774
rect -5846 611094 -5226 650538
rect -5846 610858 -5814 611094
rect -5578 610858 -5494 611094
rect -5258 610858 -5226 611094
rect -5846 610774 -5226 610858
rect -5846 610538 -5814 610774
rect -5578 610538 -5494 610774
rect -5258 610538 -5226 610774
rect -5846 571094 -5226 610538
rect -5846 570858 -5814 571094
rect -5578 570858 -5494 571094
rect -5258 570858 -5226 571094
rect -5846 570774 -5226 570858
rect -5846 570538 -5814 570774
rect -5578 570538 -5494 570774
rect -5258 570538 -5226 570774
rect -5846 531094 -5226 570538
rect -5846 530858 -5814 531094
rect -5578 530858 -5494 531094
rect -5258 530858 -5226 531094
rect -5846 530774 -5226 530858
rect -5846 530538 -5814 530774
rect -5578 530538 -5494 530774
rect -5258 530538 -5226 530774
rect -5846 491094 -5226 530538
rect -5846 490858 -5814 491094
rect -5578 490858 -5494 491094
rect -5258 490858 -5226 491094
rect -5846 490774 -5226 490858
rect -5846 490538 -5814 490774
rect -5578 490538 -5494 490774
rect -5258 490538 -5226 490774
rect -5846 451094 -5226 490538
rect -5846 450858 -5814 451094
rect -5578 450858 -5494 451094
rect -5258 450858 -5226 451094
rect -5846 450774 -5226 450858
rect -5846 450538 -5814 450774
rect -5578 450538 -5494 450774
rect -5258 450538 -5226 450774
rect -5846 411094 -5226 450538
rect -5846 410858 -5814 411094
rect -5578 410858 -5494 411094
rect -5258 410858 -5226 411094
rect -5846 410774 -5226 410858
rect -5846 410538 -5814 410774
rect -5578 410538 -5494 410774
rect -5258 410538 -5226 410774
rect -5846 371094 -5226 410538
rect -5846 370858 -5814 371094
rect -5578 370858 -5494 371094
rect -5258 370858 -5226 371094
rect -5846 370774 -5226 370858
rect -5846 370538 -5814 370774
rect -5578 370538 -5494 370774
rect -5258 370538 -5226 370774
rect -5846 331094 -5226 370538
rect -5846 330858 -5814 331094
rect -5578 330858 -5494 331094
rect -5258 330858 -5226 331094
rect -5846 330774 -5226 330858
rect -5846 330538 -5814 330774
rect -5578 330538 -5494 330774
rect -5258 330538 -5226 330774
rect -5846 291094 -5226 330538
rect -5846 290858 -5814 291094
rect -5578 290858 -5494 291094
rect -5258 290858 -5226 291094
rect -5846 290774 -5226 290858
rect -5846 290538 -5814 290774
rect -5578 290538 -5494 290774
rect -5258 290538 -5226 290774
rect -5846 251094 -5226 290538
rect -5846 250858 -5814 251094
rect -5578 250858 -5494 251094
rect -5258 250858 -5226 251094
rect -5846 250774 -5226 250858
rect -5846 250538 -5814 250774
rect -5578 250538 -5494 250774
rect -5258 250538 -5226 250774
rect -5846 211094 -5226 250538
rect -5846 210858 -5814 211094
rect -5578 210858 -5494 211094
rect -5258 210858 -5226 211094
rect -5846 210774 -5226 210858
rect -5846 210538 -5814 210774
rect -5578 210538 -5494 210774
rect -5258 210538 -5226 210774
rect -5846 171094 -5226 210538
rect -5846 170858 -5814 171094
rect -5578 170858 -5494 171094
rect -5258 170858 -5226 171094
rect -5846 170774 -5226 170858
rect -5846 170538 -5814 170774
rect -5578 170538 -5494 170774
rect -5258 170538 -5226 170774
rect -5846 131094 -5226 170538
rect -5846 130858 -5814 131094
rect -5578 130858 -5494 131094
rect -5258 130858 -5226 131094
rect -5846 130774 -5226 130858
rect -5846 130538 -5814 130774
rect -5578 130538 -5494 130774
rect -5258 130538 -5226 130774
rect -5846 91094 -5226 130538
rect -5846 90858 -5814 91094
rect -5578 90858 -5494 91094
rect -5258 90858 -5226 91094
rect -5846 90774 -5226 90858
rect -5846 90538 -5814 90774
rect -5578 90538 -5494 90774
rect -5258 90538 -5226 90774
rect -5846 51094 -5226 90538
rect -5846 50858 -5814 51094
rect -5578 50858 -5494 51094
rect -5258 50858 -5226 51094
rect -5846 50774 -5226 50858
rect -5846 50538 -5814 50774
rect -5578 50538 -5494 50774
rect -5258 50538 -5226 50774
rect -5846 11094 -5226 50538
rect -5846 10858 -5814 11094
rect -5578 10858 -5494 11094
rect -5258 10858 -5226 11094
rect -5846 10774 -5226 10858
rect -5846 10538 -5814 10774
rect -5578 10538 -5494 10774
rect -5258 10538 -5226 10774
rect -5846 -4186 -5226 10538
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 667374 -4266 707162
rect -4886 667138 -4854 667374
rect -4618 667138 -4534 667374
rect -4298 667138 -4266 667374
rect -4886 667054 -4266 667138
rect -4886 666818 -4854 667054
rect -4618 666818 -4534 667054
rect -4298 666818 -4266 667054
rect -4886 627374 -4266 666818
rect -4886 627138 -4854 627374
rect -4618 627138 -4534 627374
rect -4298 627138 -4266 627374
rect -4886 627054 -4266 627138
rect -4886 626818 -4854 627054
rect -4618 626818 -4534 627054
rect -4298 626818 -4266 627054
rect -4886 587374 -4266 626818
rect -4886 587138 -4854 587374
rect -4618 587138 -4534 587374
rect -4298 587138 -4266 587374
rect -4886 587054 -4266 587138
rect -4886 586818 -4854 587054
rect -4618 586818 -4534 587054
rect -4298 586818 -4266 587054
rect -4886 547374 -4266 586818
rect -4886 547138 -4854 547374
rect -4618 547138 -4534 547374
rect -4298 547138 -4266 547374
rect -4886 547054 -4266 547138
rect -4886 546818 -4854 547054
rect -4618 546818 -4534 547054
rect -4298 546818 -4266 547054
rect -4886 507374 -4266 546818
rect -4886 507138 -4854 507374
rect -4618 507138 -4534 507374
rect -4298 507138 -4266 507374
rect -4886 507054 -4266 507138
rect -4886 506818 -4854 507054
rect -4618 506818 -4534 507054
rect -4298 506818 -4266 507054
rect -4886 467374 -4266 506818
rect -4886 467138 -4854 467374
rect -4618 467138 -4534 467374
rect -4298 467138 -4266 467374
rect -4886 467054 -4266 467138
rect -4886 466818 -4854 467054
rect -4618 466818 -4534 467054
rect -4298 466818 -4266 467054
rect -4886 427374 -4266 466818
rect -4886 427138 -4854 427374
rect -4618 427138 -4534 427374
rect -4298 427138 -4266 427374
rect -4886 427054 -4266 427138
rect -4886 426818 -4854 427054
rect -4618 426818 -4534 427054
rect -4298 426818 -4266 427054
rect -4886 387374 -4266 426818
rect -4886 387138 -4854 387374
rect -4618 387138 -4534 387374
rect -4298 387138 -4266 387374
rect -4886 387054 -4266 387138
rect -4886 386818 -4854 387054
rect -4618 386818 -4534 387054
rect -4298 386818 -4266 387054
rect -4886 347374 -4266 386818
rect -4886 347138 -4854 347374
rect -4618 347138 -4534 347374
rect -4298 347138 -4266 347374
rect -4886 347054 -4266 347138
rect -4886 346818 -4854 347054
rect -4618 346818 -4534 347054
rect -4298 346818 -4266 347054
rect -4886 307374 -4266 346818
rect -4886 307138 -4854 307374
rect -4618 307138 -4534 307374
rect -4298 307138 -4266 307374
rect -4886 307054 -4266 307138
rect -4886 306818 -4854 307054
rect -4618 306818 -4534 307054
rect -4298 306818 -4266 307054
rect -4886 267374 -4266 306818
rect -4886 267138 -4854 267374
rect -4618 267138 -4534 267374
rect -4298 267138 -4266 267374
rect -4886 267054 -4266 267138
rect -4886 266818 -4854 267054
rect -4618 266818 -4534 267054
rect -4298 266818 -4266 267054
rect -4886 227374 -4266 266818
rect -4886 227138 -4854 227374
rect -4618 227138 -4534 227374
rect -4298 227138 -4266 227374
rect -4886 227054 -4266 227138
rect -4886 226818 -4854 227054
rect -4618 226818 -4534 227054
rect -4298 226818 -4266 227054
rect -4886 187374 -4266 226818
rect -4886 187138 -4854 187374
rect -4618 187138 -4534 187374
rect -4298 187138 -4266 187374
rect -4886 187054 -4266 187138
rect -4886 186818 -4854 187054
rect -4618 186818 -4534 187054
rect -4298 186818 -4266 187054
rect -4886 147374 -4266 186818
rect -4886 147138 -4854 147374
rect -4618 147138 -4534 147374
rect -4298 147138 -4266 147374
rect -4886 147054 -4266 147138
rect -4886 146818 -4854 147054
rect -4618 146818 -4534 147054
rect -4298 146818 -4266 147054
rect -4886 107374 -4266 146818
rect -4886 107138 -4854 107374
rect -4618 107138 -4534 107374
rect -4298 107138 -4266 107374
rect -4886 107054 -4266 107138
rect -4886 106818 -4854 107054
rect -4618 106818 -4534 107054
rect -4298 106818 -4266 107054
rect -4886 67374 -4266 106818
rect -4886 67138 -4854 67374
rect -4618 67138 -4534 67374
rect -4298 67138 -4266 67374
rect -4886 67054 -4266 67138
rect -4886 66818 -4854 67054
rect -4618 66818 -4534 67054
rect -4298 66818 -4266 67054
rect -4886 27374 -4266 66818
rect -4886 27138 -4854 27374
rect -4618 27138 -4534 27374
rect -4298 27138 -4266 27374
rect -4886 27054 -4266 27138
rect -4886 26818 -4854 27054
rect -4618 26818 -4534 27054
rect -4298 26818 -4266 27054
rect -4886 -3226 -4266 26818
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 687374 -3306 706202
rect 5714 706758 6334 707750
rect 5714 706522 5746 706758
rect 5982 706522 6066 706758
rect 6302 706522 6334 706758
rect 5714 706438 6334 706522
rect 5714 706202 5746 706438
rect 5982 706202 6066 706438
rect 6302 706202 6334 706438
rect -3926 687138 -3894 687374
rect -3658 687138 -3574 687374
rect -3338 687138 -3306 687374
rect -3926 687054 -3306 687138
rect -3926 686818 -3894 687054
rect -3658 686818 -3574 687054
rect -3338 686818 -3306 687054
rect -3926 647374 -3306 686818
rect -3926 647138 -3894 647374
rect -3658 647138 -3574 647374
rect -3338 647138 -3306 647374
rect -3926 647054 -3306 647138
rect -3926 646818 -3894 647054
rect -3658 646818 -3574 647054
rect -3338 646818 -3306 647054
rect -3926 607374 -3306 646818
rect -3926 607138 -3894 607374
rect -3658 607138 -3574 607374
rect -3338 607138 -3306 607374
rect -3926 607054 -3306 607138
rect -3926 606818 -3894 607054
rect -3658 606818 -3574 607054
rect -3338 606818 -3306 607054
rect -3926 567374 -3306 606818
rect -3926 567138 -3894 567374
rect -3658 567138 -3574 567374
rect -3338 567138 -3306 567374
rect -3926 567054 -3306 567138
rect -3926 566818 -3894 567054
rect -3658 566818 -3574 567054
rect -3338 566818 -3306 567054
rect -3926 527374 -3306 566818
rect -3926 527138 -3894 527374
rect -3658 527138 -3574 527374
rect -3338 527138 -3306 527374
rect -3926 527054 -3306 527138
rect -3926 526818 -3894 527054
rect -3658 526818 -3574 527054
rect -3338 526818 -3306 527054
rect -3926 487374 -3306 526818
rect -3926 487138 -3894 487374
rect -3658 487138 -3574 487374
rect -3338 487138 -3306 487374
rect -3926 487054 -3306 487138
rect -3926 486818 -3894 487054
rect -3658 486818 -3574 487054
rect -3338 486818 -3306 487054
rect -3926 447374 -3306 486818
rect -3926 447138 -3894 447374
rect -3658 447138 -3574 447374
rect -3338 447138 -3306 447374
rect -3926 447054 -3306 447138
rect -3926 446818 -3894 447054
rect -3658 446818 -3574 447054
rect -3338 446818 -3306 447054
rect -3926 407374 -3306 446818
rect -3926 407138 -3894 407374
rect -3658 407138 -3574 407374
rect -3338 407138 -3306 407374
rect -3926 407054 -3306 407138
rect -3926 406818 -3894 407054
rect -3658 406818 -3574 407054
rect -3338 406818 -3306 407054
rect -3926 367374 -3306 406818
rect -3926 367138 -3894 367374
rect -3658 367138 -3574 367374
rect -3338 367138 -3306 367374
rect -3926 367054 -3306 367138
rect -3926 366818 -3894 367054
rect -3658 366818 -3574 367054
rect -3338 366818 -3306 367054
rect -3926 327374 -3306 366818
rect -3926 327138 -3894 327374
rect -3658 327138 -3574 327374
rect -3338 327138 -3306 327374
rect -3926 327054 -3306 327138
rect -3926 326818 -3894 327054
rect -3658 326818 -3574 327054
rect -3338 326818 -3306 327054
rect -3926 287374 -3306 326818
rect -3926 287138 -3894 287374
rect -3658 287138 -3574 287374
rect -3338 287138 -3306 287374
rect -3926 287054 -3306 287138
rect -3926 286818 -3894 287054
rect -3658 286818 -3574 287054
rect -3338 286818 -3306 287054
rect -3926 247374 -3306 286818
rect -3926 247138 -3894 247374
rect -3658 247138 -3574 247374
rect -3338 247138 -3306 247374
rect -3926 247054 -3306 247138
rect -3926 246818 -3894 247054
rect -3658 246818 -3574 247054
rect -3338 246818 -3306 247054
rect -3926 207374 -3306 246818
rect -3926 207138 -3894 207374
rect -3658 207138 -3574 207374
rect -3338 207138 -3306 207374
rect -3926 207054 -3306 207138
rect -3926 206818 -3894 207054
rect -3658 206818 -3574 207054
rect -3338 206818 -3306 207054
rect -3926 167374 -3306 206818
rect -3926 167138 -3894 167374
rect -3658 167138 -3574 167374
rect -3338 167138 -3306 167374
rect -3926 167054 -3306 167138
rect -3926 166818 -3894 167054
rect -3658 166818 -3574 167054
rect -3338 166818 -3306 167054
rect -3926 127374 -3306 166818
rect -3926 127138 -3894 127374
rect -3658 127138 -3574 127374
rect -3338 127138 -3306 127374
rect -3926 127054 -3306 127138
rect -3926 126818 -3894 127054
rect -3658 126818 -3574 127054
rect -3338 126818 -3306 127054
rect -3926 87374 -3306 126818
rect -3926 87138 -3894 87374
rect -3658 87138 -3574 87374
rect -3338 87138 -3306 87374
rect -3926 87054 -3306 87138
rect -3926 86818 -3894 87054
rect -3658 86818 -3574 87054
rect -3338 86818 -3306 87054
rect -3926 47374 -3306 86818
rect -3926 47138 -3894 47374
rect -3658 47138 -3574 47374
rect -3338 47138 -3306 47374
rect -3926 47054 -3306 47138
rect -3926 46818 -3894 47054
rect -3658 46818 -3574 47054
rect -3338 46818 -3306 47054
rect -3926 7374 -3306 46818
rect -3926 7138 -3894 7374
rect -3658 7138 -3574 7374
rect -3338 7138 -3306 7374
rect -3926 7054 -3306 7138
rect -3926 6818 -3894 7054
rect -3658 6818 -3574 7054
rect -3338 6818 -3306 7054
rect -3926 -2266 -3306 6818
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 663654 -2346 705242
rect -2966 663418 -2934 663654
rect -2698 663418 -2614 663654
rect -2378 663418 -2346 663654
rect -2966 663334 -2346 663418
rect -2966 663098 -2934 663334
rect -2698 663098 -2614 663334
rect -2378 663098 -2346 663334
rect -2966 623654 -2346 663098
rect -2966 623418 -2934 623654
rect -2698 623418 -2614 623654
rect -2378 623418 -2346 623654
rect -2966 623334 -2346 623418
rect -2966 623098 -2934 623334
rect -2698 623098 -2614 623334
rect -2378 623098 -2346 623334
rect -2966 583654 -2346 623098
rect -2966 583418 -2934 583654
rect -2698 583418 -2614 583654
rect -2378 583418 -2346 583654
rect -2966 583334 -2346 583418
rect -2966 583098 -2934 583334
rect -2698 583098 -2614 583334
rect -2378 583098 -2346 583334
rect -2966 543654 -2346 583098
rect -2966 543418 -2934 543654
rect -2698 543418 -2614 543654
rect -2378 543418 -2346 543654
rect -2966 543334 -2346 543418
rect -2966 543098 -2934 543334
rect -2698 543098 -2614 543334
rect -2378 543098 -2346 543334
rect -2966 503654 -2346 543098
rect -2966 503418 -2934 503654
rect -2698 503418 -2614 503654
rect -2378 503418 -2346 503654
rect -2966 503334 -2346 503418
rect -2966 503098 -2934 503334
rect -2698 503098 -2614 503334
rect -2378 503098 -2346 503334
rect -2966 463654 -2346 503098
rect -2966 463418 -2934 463654
rect -2698 463418 -2614 463654
rect -2378 463418 -2346 463654
rect -2966 463334 -2346 463418
rect -2966 463098 -2934 463334
rect -2698 463098 -2614 463334
rect -2378 463098 -2346 463334
rect -2966 423654 -2346 463098
rect -2966 423418 -2934 423654
rect -2698 423418 -2614 423654
rect -2378 423418 -2346 423654
rect -2966 423334 -2346 423418
rect -2966 423098 -2934 423334
rect -2698 423098 -2614 423334
rect -2378 423098 -2346 423334
rect -2966 383654 -2346 423098
rect -2966 383418 -2934 383654
rect -2698 383418 -2614 383654
rect -2378 383418 -2346 383654
rect -2966 383334 -2346 383418
rect -2966 383098 -2934 383334
rect -2698 383098 -2614 383334
rect -2378 383098 -2346 383334
rect -2966 343654 -2346 383098
rect -2966 343418 -2934 343654
rect -2698 343418 -2614 343654
rect -2378 343418 -2346 343654
rect -2966 343334 -2346 343418
rect -2966 343098 -2934 343334
rect -2698 343098 -2614 343334
rect -2378 343098 -2346 343334
rect -2966 303654 -2346 343098
rect -2966 303418 -2934 303654
rect -2698 303418 -2614 303654
rect -2378 303418 -2346 303654
rect -2966 303334 -2346 303418
rect -2966 303098 -2934 303334
rect -2698 303098 -2614 303334
rect -2378 303098 -2346 303334
rect -2966 263654 -2346 303098
rect -2966 263418 -2934 263654
rect -2698 263418 -2614 263654
rect -2378 263418 -2346 263654
rect -2966 263334 -2346 263418
rect -2966 263098 -2934 263334
rect -2698 263098 -2614 263334
rect -2378 263098 -2346 263334
rect -2966 223654 -2346 263098
rect -2966 223418 -2934 223654
rect -2698 223418 -2614 223654
rect -2378 223418 -2346 223654
rect -2966 223334 -2346 223418
rect -2966 223098 -2934 223334
rect -2698 223098 -2614 223334
rect -2378 223098 -2346 223334
rect -2966 183654 -2346 223098
rect -2966 183418 -2934 183654
rect -2698 183418 -2614 183654
rect -2378 183418 -2346 183654
rect -2966 183334 -2346 183418
rect -2966 183098 -2934 183334
rect -2698 183098 -2614 183334
rect -2378 183098 -2346 183334
rect -2966 143654 -2346 183098
rect -2966 143418 -2934 143654
rect -2698 143418 -2614 143654
rect -2378 143418 -2346 143654
rect -2966 143334 -2346 143418
rect -2966 143098 -2934 143334
rect -2698 143098 -2614 143334
rect -2378 143098 -2346 143334
rect -2966 103654 -2346 143098
rect -2966 103418 -2934 103654
rect -2698 103418 -2614 103654
rect -2378 103418 -2346 103654
rect -2966 103334 -2346 103418
rect -2966 103098 -2934 103334
rect -2698 103098 -2614 103334
rect -2378 103098 -2346 103334
rect -2966 63654 -2346 103098
rect -2966 63418 -2934 63654
rect -2698 63418 -2614 63654
rect -2378 63418 -2346 63654
rect -2966 63334 -2346 63418
rect -2966 63098 -2934 63334
rect -2698 63098 -2614 63334
rect -2378 63098 -2346 63334
rect -2966 23654 -2346 63098
rect -2966 23418 -2934 23654
rect -2698 23418 -2614 23654
rect -2378 23418 -2346 23654
rect -2966 23334 -2346 23418
rect -2966 23098 -2934 23334
rect -2698 23098 -2614 23334
rect -2378 23098 -2346 23334
rect -2966 -1306 -2346 23098
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 683654 -1386 704282
rect 1994 704838 2614 705830
rect 1994 704602 2026 704838
rect 2262 704602 2346 704838
rect 2582 704602 2614 704838
rect 1994 704518 2614 704602
rect 1994 704282 2026 704518
rect 2262 704282 2346 704518
rect 2582 704282 2614 704518
rect 1994 700008 2614 704282
rect 5714 700008 6334 706202
rect 9434 700008 10054 708122
rect 13154 700008 13774 710042
rect 33154 711558 33774 711590
rect 33154 711322 33186 711558
rect 33422 711322 33506 711558
rect 33742 711322 33774 711558
rect 33154 711238 33774 711322
rect 33154 711002 33186 711238
rect 33422 711002 33506 711238
rect 33742 711002 33774 711238
rect 29434 709638 30054 709670
rect 29434 709402 29466 709638
rect 29702 709402 29786 709638
rect 30022 709402 30054 709638
rect 29434 709318 30054 709402
rect 29434 709082 29466 709318
rect 29702 709082 29786 709318
rect 30022 709082 30054 709318
rect 25714 707718 26334 707750
rect 25714 707482 25746 707718
rect 25982 707482 26066 707718
rect 26302 707482 26334 707718
rect 25714 707398 26334 707482
rect 25714 707162 25746 707398
rect 25982 707162 26066 707398
rect 26302 707162 26334 707398
rect 21994 705798 22614 705830
rect 21994 705562 22026 705798
rect 22262 705562 22346 705798
rect 22582 705562 22614 705798
rect 21994 705478 22614 705562
rect 21994 705242 22026 705478
rect 22262 705242 22346 705478
rect 22582 705242 22614 705478
rect 21994 700008 22614 705242
rect 25714 700008 26334 707162
rect 29434 700008 30054 709082
rect 33154 700008 33774 711002
rect 53154 710598 53774 711590
rect 53154 710362 53186 710598
rect 53422 710362 53506 710598
rect 53742 710362 53774 710598
rect 53154 710278 53774 710362
rect 53154 710042 53186 710278
rect 53422 710042 53506 710278
rect 53742 710042 53774 710278
rect 49434 708678 50054 709670
rect 49434 708442 49466 708678
rect 49702 708442 49786 708678
rect 50022 708442 50054 708678
rect 49434 708358 50054 708442
rect 49434 708122 49466 708358
rect 49702 708122 49786 708358
rect 50022 708122 50054 708358
rect 45714 706758 46334 707750
rect 45714 706522 45746 706758
rect 45982 706522 46066 706758
rect 46302 706522 46334 706758
rect 45714 706438 46334 706522
rect 45714 706202 45746 706438
rect 45982 706202 46066 706438
rect 46302 706202 46334 706438
rect 41994 704838 42614 705830
rect 41994 704602 42026 704838
rect 42262 704602 42346 704838
rect 42582 704602 42614 704838
rect 41994 704518 42614 704602
rect 41994 704282 42026 704518
rect 42262 704282 42346 704518
rect 42582 704282 42614 704518
rect 41994 700008 42614 704282
rect 45714 700008 46334 706202
rect 49434 700008 50054 708122
rect 53154 700008 53774 710042
rect 73154 711558 73774 711590
rect 73154 711322 73186 711558
rect 73422 711322 73506 711558
rect 73742 711322 73774 711558
rect 73154 711238 73774 711322
rect 73154 711002 73186 711238
rect 73422 711002 73506 711238
rect 73742 711002 73774 711238
rect 69434 709638 70054 709670
rect 69434 709402 69466 709638
rect 69702 709402 69786 709638
rect 70022 709402 70054 709638
rect 69434 709318 70054 709402
rect 69434 709082 69466 709318
rect 69702 709082 69786 709318
rect 70022 709082 70054 709318
rect 65714 707718 66334 707750
rect 65714 707482 65746 707718
rect 65982 707482 66066 707718
rect 66302 707482 66334 707718
rect 65714 707398 66334 707482
rect 65714 707162 65746 707398
rect 65982 707162 66066 707398
rect 66302 707162 66334 707398
rect 61994 705798 62614 705830
rect 61994 705562 62026 705798
rect 62262 705562 62346 705798
rect 62582 705562 62614 705798
rect 61994 705478 62614 705562
rect 61994 705242 62026 705478
rect 62262 705242 62346 705478
rect 62582 705242 62614 705478
rect 61994 700008 62614 705242
rect 65714 700008 66334 707162
rect 69434 700008 70054 709082
rect 73154 700008 73774 711002
rect 93154 710598 93774 711590
rect 93154 710362 93186 710598
rect 93422 710362 93506 710598
rect 93742 710362 93774 710598
rect 93154 710278 93774 710362
rect 93154 710042 93186 710278
rect 93422 710042 93506 710278
rect 93742 710042 93774 710278
rect 89434 708678 90054 709670
rect 89434 708442 89466 708678
rect 89702 708442 89786 708678
rect 90022 708442 90054 708678
rect 89434 708358 90054 708442
rect 89434 708122 89466 708358
rect 89702 708122 89786 708358
rect 90022 708122 90054 708358
rect 85714 706758 86334 707750
rect 85714 706522 85746 706758
rect 85982 706522 86066 706758
rect 86302 706522 86334 706758
rect 85714 706438 86334 706522
rect 85714 706202 85746 706438
rect 85982 706202 86066 706438
rect 86302 706202 86334 706438
rect 81994 704838 82614 705830
rect 81994 704602 82026 704838
rect 82262 704602 82346 704838
rect 82582 704602 82614 704838
rect 81994 704518 82614 704602
rect 81994 704282 82026 704518
rect 82262 704282 82346 704518
rect 82582 704282 82614 704518
rect 81994 700008 82614 704282
rect 85714 700008 86334 706202
rect 89434 700008 90054 708122
rect 93154 700008 93774 710042
rect 113154 711558 113774 711590
rect 113154 711322 113186 711558
rect 113422 711322 113506 711558
rect 113742 711322 113774 711558
rect 113154 711238 113774 711322
rect 113154 711002 113186 711238
rect 113422 711002 113506 711238
rect 113742 711002 113774 711238
rect 109434 709638 110054 709670
rect 109434 709402 109466 709638
rect 109702 709402 109786 709638
rect 110022 709402 110054 709638
rect 109434 709318 110054 709402
rect 109434 709082 109466 709318
rect 109702 709082 109786 709318
rect 110022 709082 110054 709318
rect 105714 707718 106334 707750
rect 105714 707482 105746 707718
rect 105982 707482 106066 707718
rect 106302 707482 106334 707718
rect 105714 707398 106334 707482
rect 105714 707162 105746 707398
rect 105982 707162 106066 707398
rect 106302 707162 106334 707398
rect 101994 705798 102614 705830
rect 101994 705562 102026 705798
rect 102262 705562 102346 705798
rect 102582 705562 102614 705798
rect 101994 705478 102614 705562
rect 101994 705242 102026 705478
rect 102262 705242 102346 705478
rect 102582 705242 102614 705478
rect 101994 700008 102614 705242
rect 105714 700008 106334 707162
rect 109434 700008 110054 709082
rect 113154 700008 113774 711002
rect 133154 710598 133774 711590
rect 133154 710362 133186 710598
rect 133422 710362 133506 710598
rect 133742 710362 133774 710598
rect 133154 710278 133774 710362
rect 133154 710042 133186 710278
rect 133422 710042 133506 710278
rect 133742 710042 133774 710278
rect 129434 708678 130054 709670
rect 129434 708442 129466 708678
rect 129702 708442 129786 708678
rect 130022 708442 130054 708678
rect 129434 708358 130054 708442
rect 129434 708122 129466 708358
rect 129702 708122 129786 708358
rect 130022 708122 130054 708358
rect 125714 706758 126334 707750
rect 125714 706522 125746 706758
rect 125982 706522 126066 706758
rect 126302 706522 126334 706758
rect 125714 706438 126334 706522
rect 125714 706202 125746 706438
rect 125982 706202 126066 706438
rect 126302 706202 126334 706438
rect 121994 704838 122614 705830
rect 121994 704602 122026 704838
rect 122262 704602 122346 704838
rect 122582 704602 122614 704838
rect 121994 704518 122614 704602
rect 121994 704282 122026 704518
rect 122262 704282 122346 704518
rect 122582 704282 122614 704518
rect 121994 700008 122614 704282
rect 125714 700008 126334 706202
rect 129434 700008 130054 708122
rect 133154 700008 133774 710042
rect 153154 711558 153774 711590
rect 153154 711322 153186 711558
rect 153422 711322 153506 711558
rect 153742 711322 153774 711558
rect 153154 711238 153774 711322
rect 153154 711002 153186 711238
rect 153422 711002 153506 711238
rect 153742 711002 153774 711238
rect 149434 709638 150054 709670
rect 149434 709402 149466 709638
rect 149702 709402 149786 709638
rect 150022 709402 150054 709638
rect 149434 709318 150054 709402
rect 149434 709082 149466 709318
rect 149702 709082 149786 709318
rect 150022 709082 150054 709318
rect 145714 707718 146334 707750
rect 145714 707482 145746 707718
rect 145982 707482 146066 707718
rect 146302 707482 146334 707718
rect 145714 707398 146334 707482
rect 145714 707162 145746 707398
rect 145982 707162 146066 707398
rect 146302 707162 146334 707398
rect 141994 705798 142614 705830
rect 141994 705562 142026 705798
rect 142262 705562 142346 705798
rect 142582 705562 142614 705798
rect 141994 705478 142614 705562
rect 141994 705242 142026 705478
rect 142262 705242 142346 705478
rect 142582 705242 142614 705478
rect 141994 700008 142614 705242
rect 145714 700008 146334 707162
rect 149434 700008 150054 709082
rect 153154 700008 153774 711002
rect 173154 710598 173774 711590
rect 173154 710362 173186 710598
rect 173422 710362 173506 710598
rect 173742 710362 173774 710598
rect 173154 710278 173774 710362
rect 173154 710042 173186 710278
rect 173422 710042 173506 710278
rect 173742 710042 173774 710278
rect 169434 708678 170054 709670
rect 169434 708442 169466 708678
rect 169702 708442 169786 708678
rect 170022 708442 170054 708678
rect 169434 708358 170054 708442
rect 169434 708122 169466 708358
rect 169702 708122 169786 708358
rect 170022 708122 170054 708358
rect 165714 706758 166334 707750
rect 165714 706522 165746 706758
rect 165982 706522 166066 706758
rect 166302 706522 166334 706758
rect 165714 706438 166334 706522
rect 165714 706202 165746 706438
rect 165982 706202 166066 706438
rect 166302 706202 166334 706438
rect 161994 704838 162614 705830
rect 161994 704602 162026 704838
rect 162262 704602 162346 704838
rect 162582 704602 162614 704838
rect 161994 704518 162614 704602
rect 161994 704282 162026 704518
rect 162262 704282 162346 704518
rect 162582 704282 162614 704518
rect 161994 700008 162614 704282
rect 165714 700008 166334 706202
rect 169434 700008 170054 708122
rect 173154 700008 173774 710042
rect 193154 711558 193774 711590
rect 193154 711322 193186 711558
rect 193422 711322 193506 711558
rect 193742 711322 193774 711558
rect 193154 711238 193774 711322
rect 193154 711002 193186 711238
rect 193422 711002 193506 711238
rect 193742 711002 193774 711238
rect 189434 709638 190054 709670
rect 189434 709402 189466 709638
rect 189702 709402 189786 709638
rect 190022 709402 190054 709638
rect 189434 709318 190054 709402
rect 189434 709082 189466 709318
rect 189702 709082 189786 709318
rect 190022 709082 190054 709318
rect 185714 707718 186334 707750
rect 185714 707482 185746 707718
rect 185982 707482 186066 707718
rect 186302 707482 186334 707718
rect 185714 707398 186334 707482
rect 185714 707162 185746 707398
rect 185982 707162 186066 707398
rect 186302 707162 186334 707398
rect 181994 705798 182614 705830
rect 181994 705562 182026 705798
rect 182262 705562 182346 705798
rect 182582 705562 182614 705798
rect 181994 705478 182614 705562
rect 181994 705242 182026 705478
rect 182262 705242 182346 705478
rect 182582 705242 182614 705478
rect 181994 700008 182614 705242
rect 185714 700008 186334 707162
rect 189434 700008 190054 709082
rect 193154 700008 193774 711002
rect 213154 710598 213774 711590
rect 213154 710362 213186 710598
rect 213422 710362 213506 710598
rect 213742 710362 213774 710598
rect 213154 710278 213774 710362
rect 213154 710042 213186 710278
rect 213422 710042 213506 710278
rect 213742 710042 213774 710278
rect 209434 708678 210054 709670
rect 209434 708442 209466 708678
rect 209702 708442 209786 708678
rect 210022 708442 210054 708678
rect 209434 708358 210054 708442
rect 209434 708122 209466 708358
rect 209702 708122 209786 708358
rect 210022 708122 210054 708358
rect 205714 706758 206334 707750
rect 205714 706522 205746 706758
rect 205982 706522 206066 706758
rect 206302 706522 206334 706758
rect 205714 706438 206334 706522
rect 205714 706202 205746 706438
rect 205982 706202 206066 706438
rect 206302 706202 206334 706438
rect 201994 704838 202614 705830
rect 201994 704602 202026 704838
rect 202262 704602 202346 704838
rect 202582 704602 202614 704838
rect 201994 704518 202614 704602
rect 201994 704282 202026 704518
rect 202262 704282 202346 704518
rect 202582 704282 202614 704518
rect 201994 700008 202614 704282
rect 205714 700008 206334 706202
rect 209434 700008 210054 708122
rect 213154 700008 213774 710042
rect 233154 711558 233774 711590
rect 233154 711322 233186 711558
rect 233422 711322 233506 711558
rect 233742 711322 233774 711558
rect 233154 711238 233774 711322
rect 233154 711002 233186 711238
rect 233422 711002 233506 711238
rect 233742 711002 233774 711238
rect 229434 709638 230054 709670
rect 229434 709402 229466 709638
rect 229702 709402 229786 709638
rect 230022 709402 230054 709638
rect 229434 709318 230054 709402
rect 229434 709082 229466 709318
rect 229702 709082 229786 709318
rect 230022 709082 230054 709318
rect 225714 707718 226334 707750
rect 225714 707482 225746 707718
rect 225982 707482 226066 707718
rect 226302 707482 226334 707718
rect 225714 707398 226334 707482
rect 225714 707162 225746 707398
rect 225982 707162 226066 707398
rect 226302 707162 226334 707398
rect 221994 705798 222614 705830
rect 221994 705562 222026 705798
rect 222262 705562 222346 705798
rect 222582 705562 222614 705798
rect 221994 705478 222614 705562
rect 221994 705242 222026 705478
rect 222262 705242 222346 705478
rect 222582 705242 222614 705478
rect 221994 700008 222614 705242
rect 225714 700008 226334 707162
rect 229434 700008 230054 709082
rect 233154 700008 233774 711002
rect 253154 710598 253774 711590
rect 253154 710362 253186 710598
rect 253422 710362 253506 710598
rect 253742 710362 253774 710598
rect 253154 710278 253774 710362
rect 253154 710042 253186 710278
rect 253422 710042 253506 710278
rect 253742 710042 253774 710278
rect 249434 708678 250054 709670
rect 249434 708442 249466 708678
rect 249702 708442 249786 708678
rect 250022 708442 250054 708678
rect 249434 708358 250054 708442
rect 249434 708122 249466 708358
rect 249702 708122 249786 708358
rect 250022 708122 250054 708358
rect 245714 706758 246334 707750
rect 245714 706522 245746 706758
rect 245982 706522 246066 706758
rect 246302 706522 246334 706758
rect 245714 706438 246334 706522
rect 245714 706202 245746 706438
rect 245982 706202 246066 706438
rect 246302 706202 246334 706438
rect 241994 704838 242614 705830
rect 241994 704602 242026 704838
rect 242262 704602 242346 704838
rect 242582 704602 242614 704838
rect 241994 704518 242614 704602
rect 241994 704282 242026 704518
rect 242262 704282 242346 704518
rect 242582 704282 242614 704518
rect 241994 700008 242614 704282
rect 245714 700008 246334 706202
rect 249434 700008 250054 708122
rect 253154 700008 253774 710042
rect 273154 711558 273774 711590
rect 273154 711322 273186 711558
rect 273422 711322 273506 711558
rect 273742 711322 273774 711558
rect 273154 711238 273774 711322
rect 273154 711002 273186 711238
rect 273422 711002 273506 711238
rect 273742 711002 273774 711238
rect 269434 709638 270054 709670
rect 269434 709402 269466 709638
rect 269702 709402 269786 709638
rect 270022 709402 270054 709638
rect 269434 709318 270054 709402
rect 269434 709082 269466 709318
rect 269702 709082 269786 709318
rect 270022 709082 270054 709318
rect 265714 707718 266334 707750
rect 265714 707482 265746 707718
rect 265982 707482 266066 707718
rect 266302 707482 266334 707718
rect 265714 707398 266334 707482
rect 265714 707162 265746 707398
rect 265982 707162 266066 707398
rect 266302 707162 266334 707398
rect 261994 705798 262614 705830
rect 261994 705562 262026 705798
rect 262262 705562 262346 705798
rect 262582 705562 262614 705798
rect 261994 705478 262614 705562
rect 261994 705242 262026 705478
rect 262262 705242 262346 705478
rect 262582 705242 262614 705478
rect 261994 700008 262614 705242
rect 265714 700008 266334 707162
rect 269434 700008 270054 709082
rect 273154 700008 273774 711002
rect 293154 710598 293774 711590
rect 293154 710362 293186 710598
rect 293422 710362 293506 710598
rect 293742 710362 293774 710598
rect 293154 710278 293774 710362
rect 293154 710042 293186 710278
rect 293422 710042 293506 710278
rect 293742 710042 293774 710278
rect 289434 708678 290054 709670
rect 289434 708442 289466 708678
rect 289702 708442 289786 708678
rect 290022 708442 290054 708678
rect 289434 708358 290054 708442
rect 289434 708122 289466 708358
rect 289702 708122 289786 708358
rect 290022 708122 290054 708358
rect 285714 706758 286334 707750
rect 285714 706522 285746 706758
rect 285982 706522 286066 706758
rect 286302 706522 286334 706758
rect 285714 706438 286334 706522
rect 285714 706202 285746 706438
rect 285982 706202 286066 706438
rect 286302 706202 286334 706438
rect 281994 704838 282614 705830
rect 281994 704602 282026 704838
rect 282262 704602 282346 704838
rect 282582 704602 282614 704838
rect 281994 704518 282614 704602
rect 281994 704282 282026 704518
rect 282262 704282 282346 704518
rect 282582 704282 282614 704518
rect 281994 700008 282614 704282
rect 285714 700008 286334 706202
rect 289434 700008 290054 708122
rect 293154 700008 293774 710042
rect 313154 711558 313774 711590
rect 313154 711322 313186 711558
rect 313422 711322 313506 711558
rect 313742 711322 313774 711558
rect 313154 711238 313774 711322
rect 313154 711002 313186 711238
rect 313422 711002 313506 711238
rect 313742 711002 313774 711238
rect 309434 709638 310054 709670
rect 309434 709402 309466 709638
rect 309702 709402 309786 709638
rect 310022 709402 310054 709638
rect 309434 709318 310054 709402
rect 309434 709082 309466 709318
rect 309702 709082 309786 709318
rect 310022 709082 310054 709318
rect 305714 707718 306334 707750
rect 305714 707482 305746 707718
rect 305982 707482 306066 707718
rect 306302 707482 306334 707718
rect 305714 707398 306334 707482
rect 305714 707162 305746 707398
rect 305982 707162 306066 707398
rect 306302 707162 306334 707398
rect 301994 705798 302614 705830
rect 301994 705562 302026 705798
rect 302262 705562 302346 705798
rect 302582 705562 302614 705798
rect 301994 705478 302614 705562
rect 301994 705242 302026 705478
rect 302262 705242 302346 705478
rect 302582 705242 302614 705478
rect 301994 700008 302614 705242
rect 305714 700008 306334 707162
rect 309434 700008 310054 709082
rect 313154 700008 313774 711002
rect 333154 710598 333774 711590
rect 333154 710362 333186 710598
rect 333422 710362 333506 710598
rect 333742 710362 333774 710598
rect 333154 710278 333774 710362
rect 333154 710042 333186 710278
rect 333422 710042 333506 710278
rect 333742 710042 333774 710278
rect 329434 708678 330054 709670
rect 329434 708442 329466 708678
rect 329702 708442 329786 708678
rect 330022 708442 330054 708678
rect 329434 708358 330054 708442
rect 329434 708122 329466 708358
rect 329702 708122 329786 708358
rect 330022 708122 330054 708358
rect 325714 706758 326334 707750
rect 325714 706522 325746 706758
rect 325982 706522 326066 706758
rect 326302 706522 326334 706758
rect 325714 706438 326334 706522
rect 325714 706202 325746 706438
rect 325982 706202 326066 706438
rect 326302 706202 326334 706438
rect 321994 704838 322614 705830
rect 321994 704602 322026 704838
rect 322262 704602 322346 704838
rect 322582 704602 322614 704838
rect 321994 704518 322614 704602
rect 321994 704282 322026 704518
rect 322262 704282 322346 704518
rect 322582 704282 322614 704518
rect 321994 700008 322614 704282
rect 325714 700008 326334 706202
rect 329434 700008 330054 708122
rect 333154 700008 333774 710042
rect 353154 711558 353774 711590
rect 353154 711322 353186 711558
rect 353422 711322 353506 711558
rect 353742 711322 353774 711558
rect 353154 711238 353774 711322
rect 353154 711002 353186 711238
rect 353422 711002 353506 711238
rect 353742 711002 353774 711238
rect 349434 709638 350054 709670
rect 349434 709402 349466 709638
rect 349702 709402 349786 709638
rect 350022 709402 350054 709638
rect 349434 709318 350054 709402
rect 349434 709082 349466 709318
rect 349702 709082 349786 709318
rect 350022 709082 350054 709318
rect 345714 707718 346334 707750
rect 345714 707482 345746 707718
rect 345982 707482 346066 707718
rect 346302 707482 346334 707718
rect 345714 707398 346334 707482
rect 345714 707162 345746 707398
rect 345982 707162 346066 707398
rect 346302 707162 346334 707398
rect 341994 705798 342614 705830
rect 341994 705562 342026 705798
rect 342262 705562 342346 705798
rect 342582 705562 342614 705798
rect 341994 705478 342614 705562
rect 341994 705242 342026 705478
rect 342262 705242 342346 705478
rect 342582 705242 342614 705478
rect 341994 700008 342614 705242
rect 345714 700008 346334 707162
rect 349434 700008 350054 709082
rect 353154 700008 353774 711002
rect 373154 710598 373774 711590
rect 373154 710362 373186 710598
rect 373422 710362 373506 710598
rect 373742 710362 373774 710598
rect 373154 710278 373774 710362
rect 373154 710042 373186 710278
rect 373422 710042 373506 710278
rect 373742 710042 373774 710278
rect 369434 708678 370054 709670
rect 369434 708442 369466 708678
rect 369702 708442 369786 708678
rect 370022 708442 370054 708678
rect 369434 708358 370054 708442
rect 369434 708122 369466 708358
rect 369702 708122 369786 708358
rect 370022 708122 370054 708358
rect 365714 706758 366334 707750
rect 365714 706522 365746 706758
rect 365982 706522 366066 706758
rect 366302 706522 366334 706758
rect 365714 706438 366334 706522
rect 365714 706202 365746 706438
rect 365982 706202 366066 706438
rect 366302 706202 366334 706438
rect 361994 704838 362614 705830
rect 361994 704602 362026 704838
rect 362262 704602 362346 704838
rect 362582 704602 362614 704838
rect 361994 704518 362614 704602
rect 361994 704282 362026 704518
rect 362262 704282 362346 704518
rect 362582 704282 362614 704518
rect 361994 700008 362614 704282
rect 365714 700008 366334 706202
rect 369434 700008 370054 708122
rect 373154 700008 373774 710042
rect 393154 711558 393774 711590
rect 393154 711322 393186 711558
rect 393422 711322 393506 711558
rect 393742 711322 393774 711558
rect 393154 711238 393774 711322
rect 393154 711002 393186 711238
rect 393422 711002 393506 711238
rect 393742 711002 393774 711238
rect 389434 709638 390054 709670
rect 389434 709402 389466 709638
rect 389702 709402 389786 709638
rect 390022 709402 390054 709638
rect 389434 709318 390054 709402
rect 389434 709082 389466 709318
rect 389702 709082 389786 709318
rect 390022 709082 390054 709318
rect 385714 707718 386334 707750
rect 385714 707482 385746 707718
rect 385982 707482 386066 707718
rect 386302 707482 386334 707718
rect 385714 707398 386334 707482
rect 385714 707162 385746 707398
rect 385982 707162 386066 707398
rect 386302 707162 386334 707398
rect 381994 705798 382614 705830
rect 381994 705562 382026 705798
rect 382262 705562 382346 705798
rect 382582 705562 382614 705798
rect 381994 705478 382614 705562
rect 381994 705242 382026 705478
rect 382262 705242 382346 705478
rect 382582 705242 382614 705478
rect 381994 700008 382614 705242
rect 385714 700008 386334 707162
rect 389434 700008 390054 709082
rect 393154 700008 393774 711002
rect 413154 710598 413774 711590
rect 413154 710362 413186 710598
rect 413422 710362 413506 710598
rect 413742 710362 413774 710598
rect 413154 710278 413774 710362
rect 413154 710042 413186 710278
rect 413422 710042 413506 710278
rect 413742 710042 413774 710278
rect 409434 708678 410054 709670
rect 409434 708442 409466 708678
rect 409702 708442 409786 708678
rect 410022 708442 410054 708678
rect 409434 708358 410054 708442
rect 409434 708122 409466 708358
rect 409702 708122 409786 708358
rect 410022 708122 410054 708358
rect 405714 706758 406334 707750
rect 405714 706522 405746 706758
rect 405982 706522 406066 706758
rect 406302 706522 406334 706758
rect 405714 706438 406334 706522
rect 405714 706202 405746 706438
rect 405982 706202 406066 706438
rect 406302 706202 406334 706438
rect 401994 704838 402614 705830
rect 401994 704602 402026 704838
rect 402262 704602 402346 704838
rect 402582 704602 402614 704838
rect 401994 704518 402614 704602
rect 401994 704282 402026 704518
rect 402262 704282 402346 704518
rect 402582 704282 402614 704518
rect 401994 700008 402614 704282
rect 405714 700008 406334 706202
rect 409434 700008 410054 708122
rect 413154 700008 413774 710042
rect 433154 711558 433774 711590
rect 433154 711322 433186 711558
rect 433422 711322 433506 711558
rect 433742 711322 433774 711558
rect 433154 711238 433774 711322
rect 433154 711002 433186 711238
rect 433422 711002 433506 711238
rect 433742 711002 433774 711238
rect 429434 709638 430054 709670
rect 429434 709402 429466 709638
rect 429702 709402 429786 709638
rect 430022 709402 430054 709638
rect 429434 709318 430054 709402
rect 429434 709082 429466 709318
rect 429702 709082 429786 709318
rect 430022 709082 430054 709318
rect 425714 707718 426334 707750
rect 425714 707482 425746 707718
rect 425982 707482 426066 707718
rect 426302 707482 426334 707718
rect 425714 707398 426334 707482
rect 425714 707162 425746 707398
rect 425982 707162 426066 707398
rect 426302 707162 426334 707398
rect 421994 705798 422614 705830
rect 421994 705562 422026 705798
rect 422262 705562 422346 705798
rect 422582 705562 422614 705798
rect 421994 705478 422614 705562
rect 421994 705242 422026 705478
rect 422262 705242 422346 705478
rect 422582 705242 422614 705478
rect 421994 700008 422614 705242
rect 425714 700008 426334 707162
rect 429434 700008 430054 709082
rect 433154 700008 433774 711002
rect 453154 710598 453774 711590
rect 453154 710362 453186 710598
rect 453422 710362 453506 710598
rect 453742 710362 453774 710598
rect 453154 710278 453774 710362
rect 453154 710042 453186 710278
rect 453422 710042 453506 710278
rect 453742 710042 453774 710278
rect 449434 708678 450054 709670
rect 449434 708442 449466 708678
rect 449702 708442 449786 708678
rect 450022 708442 450054 708678
rect 449434 708358 450054 708442
rect 449434 708122 449466 708358
rect 449702 708122 449786 708358
rect 450022 708122 450054 708358
rect 445714 706758 446334 707750
rect 445714 706522 445746 706758
rect 445982 706522 446066 706758
rect 446302 706522 446334 706758
rect 445714 706438 446334 706522
rect 445714 706202 445746 706438
rect 445982 706202 446066 706438
rect 446302 706202 446334 706438
rect 441994 704838 442614 705830
rect 441994 704602 442026 704838
rect 442262 704602 442346 704838
rect 442582 704602 442614 704838
rect 441994 704518 442614 704602
rect 441994 704282 442026 704518
rect 442262 704282 442346 704518
rect 442582 704282 442614 704518
rect 441994 700008 442614 704282
rect 445714 700008 446334 706202
rect 449434 700008 450054 708122
rect 453154 700008 453774 710042
rect 473154 711558 473774 711590
rect 473154 711322 473186 711558
rect 473422 711322 473506 711558
rect 473742 711322 473774 711558
rect 473154 711238 473774 711322
rect 473154 711002 473186 711238
rect 473422 711002 473506 711238
rect 473742 711002 473774 711238
rect 469434 709638 470054 709670
rect 469434 709402 469466 709638
rect 469702 709402 469786 709638
rect 470022 709402 470054 709638
rect 469434 709318 470054 709402
rect 469434 709082 469466 709318
rect 469702 709082 469786 709318
rect 470022 709082 470054 709318
rect 465714 707718 466334 707750
rect 465714 707482 465746 707718
rect 465982 707482 466066 707718
rect 466302 707482 466334 707718
rect 465714 707398 466334 707482
rect 465714 707162 465746 707398
rect 465982 707162 466066 707398
rect 466302 707162 466334 707398
rect 461994 705798 462614 705830
rect 461994 705562 462026 705798
rect 462262 705562 462346 705798
rect 462582 705562 462614 705798
rect 461994 705478 462614 705562
rect 461994 705242 462026 705478
rect 462262 705242 462346 705478
rect 462582 705242 462614 705478
rect 461994 700008 462614 705242
rect 465714 700008 466334 707162
rect 469434 700008 470054 709082
rect 473154 700008 473774 711002
rect 493154 710598 493774 711590
rect 493154 710362 493186 710598
rect 493422 710362 493506 710598
rect 493742 710362 493774 710598
rect 493154 710278 493774 710362
rect 493154 710042 493186 710278
rect 493422 710042 493506 710278
rect 493742 710042 493774 710278
rect 489434 708678 490054 709670
rect 489434 708442 489466 708678
rect 489702 708442 489786 708678
rect 490022 708442 490054 708678
rect 489434 708358 490054 708442
rect 489434 708122 489466 708358
rect 489702 708122 489786 708358
rect 490022 708122 490054 708358
rect 485714 706758 486334 707750
rect 485714 706522 485746 706758
rect 485982 706522 486066 706758
rect 486302 706522 486334 706758
rect 485714 706438 486334 706522
rect 485714 706202 485746 706438
rect 485982 706202 486066 706438
rect 486302 706202 486334 706438
rect 481994 704838 482614 705830
rect 481994 704602 482026 704838
rect 482262 704602 482346 704838
rect 482582 704602 482614 704838
rect 481994 704518 482614 704602
rect 481994 704282 482026 704518
rect 482262 704282 482346 704518
rect 482582 704282 482614 704518
rect 481994 700008 482614 704282
rect 485714 700008 486334 706202
rect 489434 700008 490054 708122
rect 493154 700008 493774 710042
rect 513154 711558 513774 711590
rect 513154 711322 513186 711558
rect 513422 711322 513506 711558
rect 513742 711322 513774 711558
rect 513154 711238 513774 711322
rect 513154 711002 513186 711238
rect 513422 711002 513506 711238
rect 513742 711002 513774 711238
rect 509434 709638 510054 709670
rect 509434 709402 509466 709638
rect 509702 709402 509786 709638
rect 510022 709402 510054 709638
rect 509434 709318 510054 709402
rect 509434 709082 509466 709318
rect 509702 709082 509786 709318
rect 510022 709082 510054 709318
rect 505714 707718 506334 707750
rect 505714 707482 505746 707718
rect 505982 707482 506066 707718
rect 506302 707482 506334 707718
rect 505714 707398 506334 707482
rect 505714 707162 505746 707398
rect 505982 707162 506066 707398
rect 506302 707162 506334 707398
rect 501994 705798 502614 705830
rect 501994 705562 502026 705798
rect 502262 705562 502346 705798
rect 502582 705562 502614 705798
rect 501994 705478 502614 705562
rect 501994 705242 502026 705478
rect 502262 705242 502346 705478
rect 502582 705242 502614 705478
rect 501994 700008 502614 705242
rect 505714 700008 506334 707162
rect 509434 700008 510054 709082
rect 513154 700008 513774 711002
rect 533154 710598 533774 711590
rect 533154 710362 533186 710598
rect 533422 710362 533506 710598
rect 533742 710362 533774 710598
rect 533154 710278 533774 710362
rect 533154 710042 533186 710278
rect 533422 710042 533506 710278
rect 533742 710042 533774 710278
rect 529434 708678 530054 709670
rect 529434 708442 529466 708678
rect 529702 708442 529786 708678
rect 530022 708442 530054 708678
rect 529434 708358 530054 708442
rect 529434 708122 529466 708358
rect 529702 708122 529786 708358
rect 530022 708122 530054 708358
rect 525714 706758 526334 707750
rect 525714 706522 525746 706758
rect 525982 706522 526066 706758
rect 526302 706522 526334 706758
rect 525714 706438 526334 706522
rect 525714 706202 525746 706438
rect 525982 706202 526066 706438
rect 526302 706202 526334 706438
rect 521994 704838 522614 705830
rect 521994 704602 522026 704838
rect 522262 704602 522346 704838
rect 522582 704602 522614 704838
rect 521994 704518 522614 704602
rect 521994 704282 522026 704518
rect 522262 704282 522346 704518
rect 522582 704282 522614 704518
rect 521994 700008 522614 704282
rect 525714 700008 526334 706202
rect 529434 700008 530054 708122
rect 533154 700008 533774 710042
rect 553154 711558 553774 711590
rect 553154 711322 553186 711558
rect 553422 711322 553506 711558
rect 553742 711322 553774 711558
rect 553154 711238 553774 711322
rect 553154 711002 553186 711238
rect 553422 711002 553506 711238
rect 553742 711002 553774 711238
rect 549434 709638 550054 709670
rect 549434 709402 549466 709638
rect 549702 709402 549786 709638
rect 550022 709402 550054 709638
rect 549434 709318 550054 709402
rect 549434 709082 549466 709318
rect 549702 709082 549786 709318
rect 550022 709082 550054 709318
rect 545714 707718 546334 707750
rect 545714 707482 545746 707718
rect 545982 707482 546066 707718
rect 546302 707482 546334 707718
rect 545714 707398 546334 707482
rect 545714 707162 545746 707398
rect 545982 707162 546066 707398
rect 546302 707162 546334 707398
rect 541994 705798 542614 705830
rect 541994 705562 542026 705798
rect 542262 705562 542346 705798
rect 542582 705562 542614 705798
rect 541994 705478 542614 705562
rect 541994 705242 542026 705478
rect 542262 705242 542346 705478
rect 542582 705242 542614 705478
rect 541994 700008 542614 705242
rect 545714 700008 546334 707162
rect 549434 700008 550054 709082
rect 553154 700008 553774 711002
rect 573154 710598 573774 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 573154 710362 573186 710598
rect 573422 710362 573506 710598
rect 573742 710362 573774 710598
rect 573154 710278 573774 710362
rect 573154 710042 573186 710278
rect 573422 710042 573506 710278
rect 573742 710042 573774 710278
rect 569434 708678 570054 709670
rect 569434 708442 569466 708678
rect 569702 708442 569786 708678
rect 570022 708442 570054 708678
rect 569434 708358 570054 708442
rect 569434 708122 569466 708358
rect 569702 708122 569786 708358
rect 570022 708122 570054 708358
rect 565714 706758 566334 707750
rect 565714 706522 565746 706758
rect 565982 706522 566066 706758
rect 566302 706522 566334 706758
rect 565714 706438 566334 706522
rect 565714 706202 565746 706438
rect 565982 706202 566066 706438
rect 566302 706202 566334 706438
rect 561994 704838 562614 705830
rect 561994 704602 562026 704838
rect 562262 704602 562346 704838
rect 562582 704602 562614 704838
rect 561994 704518 562614 704602
rect 561994 704282 562026 704518
rect 562262 704282 562346 704518
rect 562582 704282 562614 704518
rect 561994 700008 562614 704282
rect 565714 700008 566334 706202
rect 569434 700008 570054 708122
rect 573154 700008 573774 710042
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 683418 -1974 683654
rect -1738 683418 -1654 683654
rect -1418 683418 -1386 683654
rect -2006 683334 -1386 683418
rect -2006 683098 -1974 683334
rect -1738 683098 -1654 683334
rect -1418 683098 -1386 683334
rect -2006 643654 -1386 683098
rect 9084 683654 9704 683686
rect 9084 683418 9116 683654
rect 9352 683418 9436 683654
rect 9672 683418 9704 683654
rect 9084 683334 9704 683418
rect 9084 683098 9116 683334
rect 9352 683098 9436 683334
rect 9672 683098 9704 683334
rect 9084 683066 9704 683098
rect 56620 683654 57240 683686
rect 56620 683418 56652 683654
rect 56888 683418 56972 683654
rect 57208 683418 57240 683654
rect 56620 683334 57240 683418
rect 56620 683098 56652 683334
rect 56888 683098 56972 683334
rect 57208 683098 57240 683334
rect 56620 683066 57240 683098
rect 92620 683654 93240 683686
rect 92620 683418 92652 683654
rect 92888 683418 92972 683654
rect 93208 683418 93240 683654
rect 92620 683334 93240 683418
rect 92620 683098 92652 683334
rect 92888 683098 92972 683334
rect 93208 683098 93240 683334
rect 92620 683066 93240 683098
rect 128620 683654 129240 683686
rect 128620 683418 128652 683654
rect 128888 683418 128972 683654
rect 129208 683418 129240 683654
rect 128620 683334 129240 683418
rect 128620 683098 128652 683334
rect 128888 683098 128972 683334
rect 129208 683098 129240 683334
rect 128620 683066 129240 683098
rect 164620 683654 165240 683686
rect 164620 683418 164652 683654
rect 164888 683418 164972 683654
rect 165208 683418 165240 683654
rect 164620 683334 165240 683418
rect 164620 683098 164652 683334
rect 164888 683098 164972 683334
rect 165208 683098 165240 683334
rect 164620 683066 165240 683098
rect 200620 683654 201240 683686
rect 200620 683418 200652 683654
rect 200888 683418 200972 683654
rect 201208 683418 201240 683654
rect 200620 683334 201240 683418
rect 200620 683098 200652 683334
rect 200888 683098 200972 683334
rect 201208 683098 201240 683334
rect 200620 683066 201240 683098
rect 236620 683654 237240 683686
rect 236620 683418 236652 683654
rect 236888 683418 236972 683654
rect 237208 683418 237240 683654
rect 236620 683334 237240 683418
rect 236620 683098 236652 683334
rect 236888 683098 236972 683334
rect 237208 683098 237240 683334
rect 236620 683066 237240 683098
rect 272620 683654 273240 683686
rect 272620 683418 272652 683654
rect 272888 683418 272972 683654
rect 273208 683418 273240 683654
rect 272620 683334 273240 683418
rect 272620 683098 272652 683334
rect 272888 683098 272972 683334
rect 273208 683098 273240 683334
rect 272620 683066 273240 683098
rect 308620 683654 309240 683686
rect 308620 683418 308652 683654
rect 308888 683418 308972 683654
rect 309208 683418 309240 683654
rect 308620 683334 309240 683418
rect 308620 683098 308652 683334
rect 308888 683098 308972 683334
rect 309208 683098 309240 683334
rect 308620 683066 309240 683098
rect 344620 683654 345240 683686
rect 344620 683418 344652 683654
rect 344888 683418 344972 683654
rect 345208 683418 345240 683654
rect 344620 683334 345240 683418
rect 344620 683098 344652 683334
rect 344888 683098 344972 683334
rect 345208 683098 345240 683334
rect 344620 683066 345240 683098
rect 380620 683654 381240 683686
rect 380620 683418 380652 683654
rect 380888 683418 380972 683654
rect 381208 683418 381240 683654
rect 380620 683334 381240 683418
rect 380620 683098 380652 683334
rect 380888 683098 380972 683334
rect 381208 683098 381240 683334
rect 380620 683066 381240 683098
rect 416620 683654 417240 683686
rect 416620 683418 416652 683654
rect 416888 683418 416972 683654
rect 417208 683418 417240 683654
rect 416620 683334 417240 683418
rect 416620 683098 416652 683334
rect 416888 683098 416972 683334
rect 417208 683098 417240 683334
rect 416620 683066 417240 683098
rect 452620 683654 453240 683686
rect 452620 683418 452652 683654
rect 452888 683418 452972 683654
rect 453208 683418 453240 683654
rect 452620 683334 453240 683418
rect 452620 683098 452652 683334
rect 452888 683098 452972 683334
rect 453208 683098 453240 683334
rect 452620 683066 453240 683098
rect 488620 683654 489240 683686
rect 488620 683418 488652 683654
rect 488888 683418 488972 683654
rect 489208 683418 489240 683654
rect 488620 683334 489240 683418
rect 488620 683098 488652 683334
rect 488888 683098 488972 683334
rect 489208 683098 489240 683334
rect 488620 683066 489240 683098
rect 524620 683654 525240 683686
rect 524620 683418 524652 683654
rect 524888 683418 524972 683654
rect 525208 683418 525240 683654
rect 524620 683334 525240 683418
rect 524620 683098 524652 683334
rect 524888 683098 524972 683334
rect 525208 683098 525240 683334
rect 524620 683066 525240 683098
rect 560620 683654 561240 683686
rect 560620 683418 560652 683654
rect 560888 683418 560972 683654
rect 561208 683418 561240 683654
rect 560620 683334 561240 683418
rect 560620 683098 560652 683334
rect 560888 683098 560972 683334
rect 561208 683098 561240 683334
rect 560620 683066 561240 683098
rect 570260 683654 570880 683686
rect 570260 683418 570292 683654
rect 570528 683418 570612 683654
rect 570848 683418 570880 683654
rect 570260 683334 570880 683418
rect 570260 683098 570292 683334
rect 570528 683098 570612 683334
rect 570848 683098 570880 683334
rect 570260 683066 570880 683098
rect 585310 683654 585930 704282
rect 585310 683418 585342 683654
rect 585578 683418 585662 683654
rect 585898 683418 585930 683654
rect 585310 683334 585930 683418
rect 585310 683098 585342 683334
rect 585578 683098 585662 683334
rect 585898 683098 585930 683334
rect 7844 663654 8464 663686
rect 7844 663418 7876 663654
rect 8112 663418 8196 663654
rect 8432 663418 8464 663654
rect 7844 663334 8464 663418
rect 7844 663098 7876 663334
rect 8112 663098 8196 663334
rect 8432 663098 8464 663334
rect 7844 663066 8464 663098
rect 38000 663654 38620 663686
rect 38000 663418 38032 663654
rect 38268 663418 38352 663654
rect 38588 663418 38620 663654
rect 38000 663334 38620 663418
rect 38000 663098 38032 663334
rect 38268 663098 38352 663334
rect 38588 663098 38620 663334
rect 38000 663066 38620 663098
rect 74000 663654 74620 663686
rect 74000 663418 74032 663654
rect 74268 663418 74352 663654
rect 74588 663418 74620 663654
rect 74000 663334 74620 663418
rect 74000 663098 74032 663334
rect 74268 663098 74352 663334
rect 74588 663098 74620 663334
rect 74000 663066 74620 663098
rect 110000 663654 110620 663686
rect 110000 663418 110032 663654
rect 110268 663418 110352 663654
rect 110588 663418 110620 663654
rect 110000 663334 110620 663418
rect 110000 663098 110032 663334
rect 110268 663098 110352 663334
rect 110588 663098 110620 663334
rect 110000 663066 110620 663098
rect 146000 663654 146620 663686
rect 146000 663418 146032 663654
rect 146268 663418 146352 663654
rect 146588 663418 146620 663654
rect 146000 663334 146620 663418
rect 146000 663098 146032 663334
rect 146268 663098 146352 663334
rect 146588 663098 146620 663334
rect 146000 663066 146620 663098
rect 182000 663654 182620 663686
rect 182000 663418 182032 663654
rect 182268 663418 182352 663654
rect 182588 663418 182620 663654
rect 182000 663334 182620 663418
rect 182000 663098 182032 663334
rect 182268 663098 182352 663334
rect 182588 663098 182620 663334
rect 182000 663066 182620 663098
rect 218000 663654 218620 663686
rect 218000 663418 218032 663654
rect 218268 663418 218352 663654
rect 218588 663418 218620 663654
rect 218000 663334 218620 663418
rect 218000 663098 218032 663334
rect 218268 663098 218352 663334
rect 218588 663098 218620 663334
rect 218000 663066 218620 663098
rect 254000 663654 254620 663686
rect 254000 663418 254032 663654
rect 254268 663418 254352 663654
rect 254588 663418 254620 663654
rect 254000 663334 254620 663418
rect 254000 663098 254032 663334
rect 254268 663098 254352 663334
rect 254588 663098 254620 663334
rect 254000 663066 254620 663098
rect 290000 663654 290620 663686
rect 290000 663418 290032 663654
rect 290268 663418 290352 663654
rect 290588 663418 290620 663654
rect 290000 663334 290620 663418
rect 290000 663098 290032 663334
rect 290268 663098 290352 663334
rect 290588 663098 290620 663334
rect 290000 663066 290620 663098
rect 326000 663654 326620 663686
rect 326000 663418 326032 663654
rect 326268 663418 326352 663654
rect 326588 663418 326620 663654
rect 326000 663334 326620 663418
rect 326000 663098 326032 663334
rect 326268 663098 326352 663334
rect 326588 663098 326620 663334
rect 326000 663066 326620 663098
rect 362000 663654 362620 663686
rect 362000 663418 362032 663654
rect 362268 663418 362352 663654
rect 362588 663418 362620 663654
rect 362000 663334 362620 663418
rect 362000 663098 362032 663334
rect 362268 663098 362352 663334
rect 362588 663098 362620 663334
rect 362000 663066 362620 663098
rect 398000 663654 398620 663686
rect 398000 663418 398032 663654
rect 398268 663418 398352 663654
rect 398588 663418 398620 663654
rect 398000 663334 398620 663418
rect 398000 663098 398032 663334
rect 398268 663098 398352 663334
rect 398588 663098 398620 663334
rect 398000 663066 398620 663098
rect 434000 663654 434620 663686
rect 434000 663418 434032 663654
rect 434268 663418 434352 663654
rect 434588 663418 434620 663654
rect 434000 663334 434620 663418
rect 434000 663098 434032 663334
rect 434268 663098 434352 663334
rect 434588 663098 434620 663334
rect 434000 663066 434620 663098
rect 470000 663654 470620 663686
rect 470000 663418 470032 663654
rect 470268 663418 470352 663654
rect 470588 663418 470620 663654
rect 470000 663334 470620 663418
rect 470000 663098 470032 663334
rect 470268 663098 470352 663334
rect 470588 663098 470620 663334
rect 470000 663066 470620 663098
rect 506000 663654 506620 663686
rect 506000 663418 506032 663654
rect 506268 663418 506352 663654
rect 506588 663418 506620 663654
rect 506000 663334 506620 663418
rect 506000 663098 506032 663334
rect 506268 663098 506352 663334
rect 506588 663098 506620 663334
rect 506000 663066 506620 663098
rect 542000 663654 542620 663686
rect 542000 663418 542032 663654
rect 542268 663418 542352 663654
rect 542588 663418 542620 663654
rect 542000 663334 542620 663418
rect 542000 663098 542032 663334
rect 542268 663098 542352 663334
rect 542588 663098 542620 663334
rect 542000 663066 542620 663098
rect 571500 663654 572120 663686
rect 571500 663418 571532 663654
rect 571768 663418 571852 663654
rect 572088 663418 572120 663654
rect 571500 663334 572120 663418
rect 571500 663098 571532 663334
rect 571768 663098 571852 663334
rect 572088 663098 572120 663334
rect 571500 663066 572120 663098
rect -2006 643418 -1974 643654
rect -1738 643418 -1654 643654
rect -1418 643418 -1386 643654
rect -2006 643334 -1386 643418
rect -2006 643098 -1974 643334
rect -1738 643098 -1654 643334
rect -1418 643098 -1386 643334
rect -2006 603654 -1386 643098
rect 9084 643654 9704 643686
rect 9084 643418 9116 643654
rect 9352 643418 9436 643654
rect 9672 643418 9704 643654
rect 9084 643334 9704 643418
rect 9084 643098 9116 643334
rect 9352 643098 9436 643334
rect 9672 643098 9704 643334
rect 9084 643066 9704 643098
rect 56620 643654 57240 643686
rect 56620 643418 56652 643654
rect 56888 643418 56972 643654
rect 57208 643418 57240 643654
rect 56620 643334 57240 643418
rect 56620 643098 56652 643334
rect 56888 643098 56972 643334
rect 57208 643098 57240 643334
rect 56620 643066 57240 643098
rect 92620 643654 93240 643686
rect 92620 643418 92652 643654
rect 92888 643418 92972 643654
rect 93208 643418 93240 643654
rect 92620 643334 93240 643418
rect 92620 643098 92652 643334
rect 92888 643098 92972 643334
rect 93208 643098 93240 643334
rect 92620 643066 93240 643098
rect 128620 643654 129240 643686
rect 128620 643418 128652 643654
rect 128888 643418 128972 643654
rect 129208 643418 129240 643654
rect 128620 643334 129240 643418
rect 128620 643098 128652 643334
rect 128888 643098 128972 643334
rect 129208 643098 129240 643334
rect 128620 643066 129240 643098
rect 164620 643654 165240 643686
rect 164620 643418 164652 643654
rect 164888 643418 164972 643654
rect 165208 643418 165240 643654
rect 164620 643334 165240 643418
rect 164620 643098 164652 643334
rect 164888 643098 164972 643334
rect 165208 643098 165240 643334
rect 164620 643066 165240 643098
rect 200620 643654 201240 643686
rect 200620 643418 200652 643654
rect 200888 643418 200972 643654
rect 201208 643418 201240 643654
rect 200620 643334 201240 643418
rect 200620 643098 200652 643334
rect 200888 643098 200972 643334
rect 201208 643098 201240 643334
rect 200620 643066 201240 643098
rect 236620 643654 237240 643686
rect 236620 643418 236652 643654
rect 236888 643418 236972 643654
rect 237208 643418 237240 643654
rect 236620 643334 237240 643418
rect 236620 643098 236652 643334
rect 236888 643098 236972 643334
rect 237208 643098 237240 643334
rect 236620 643066 237240 643098
rect 272620 643654 273240 643686
rect 272620 643418 272652 643654
rect 272888 643418 272972 643654
rect 273208 643418 273240 643654
rect 272620 643334 273240 643418
rect 272620 643098 272652 643334
rect 272888 643098 272972 643334
rect 273208 643098 273240 643334
rect 272620 643066 273240 643098
rect 308620 643654 309240 643686
rect 308620 643418 308652 643654
rect 308888 643418 308972 643654
rect 309208 643418 309240 643654
rect 308620 643334 309240 643418
rect 308620 643098 308652 643334
rect 308888 643098 308972 643334
rect 309208 643098 309240 643334
rect 308620 643066 309240 643098
rect 344620 643654 345240 643686
rect 344620 643418 344652 643654
rect 344888 643418 344972 643654
rect 345208 643418 345240 643654
rect 344620 643334 345240 643418
rect 344620 643098 344652 643334
rect 344888 643098 344972 643334
rect 345208 643098 345240 643334
rect 344620 643066 345240 643098
rect 380620 643654 381240 643686
rect 380620 643418 380652 643654
rect 380888 643418 380972 643654
rect 381208 643418 381240 643654
rect 380620 643334 381240 643418
rect 380620 643098 380652 643334
rect 380888 643098 380972 643334
rect 381208 643098 381240 643334
rect 380620 643066 381240 643098
rect 416620 643654 417240 643686
rect 416620 643418 416652 643654
rect 416888 643418 416972 643654
rect 417208 643418 417240 643654
rect 416620 643334 417240 643418
rect 416620 643098 416652 643334
rect 416888 643098 416972 643334
rect 417208 643098 417240 643334
rect 416620 643066 417240 643098
rect 452620 643654 453240 643686
rect 452620 643418 452652 643654
rect 452888 643418 452972 643654
rect 453208 643418 453240 643654
rect 452620 643334 453240 643418
rect 452620 643098 452652 643334
rect 452888 643098 452972 643334
rect 453208 643098 453240 643334
rect 452620 643066 453240 643098
rect 488620 643654 489240 643686
rect 488620 643418 488652 643654
rect 488888 643418 488972 643654
rect 489208 643418 489240 643654
rect 488620 643334 489240 643418
rect 488620 643098 488652 643334
rect 488888 643098 488972 643334
rect 489208 643098 489240 643334
rect 488620 643066 489240 643098
rect 524620 643654 525240 643686
rect 524620 643418 524652 643654
rect 524888 643418 524972 643654
rect 525208 643418 525240 643654
rect 524620 643334 525240 643418
rect 524620 643098 524652 643334
rect 524888 643098 524972 643334
rect 525208 643098 525240 643334
rect 524620 643066 525240 643098
rect 560620 643654 561240 643686
rect 560620 643418 560652 643654
rect 560888 643418 560972 643654
rect 561208 643418 561240 643654
rect 560620 643334 561240 643418
rect 560620 643098 560652 643334
rect 560888 643098 560972 643334
rect 561208 643098 561240 643334
rect 560620 643066 561240 643098
rect 570260 643654 570880 643686
rect 570260 643418 570292 643654
rect 570528 643418 570612 643654
rect 570848 643418 570880 643654
rect 570260 643334 570880 643418
rect 570260 643098 570292 643334
rect 570528 643098 570612 643334
rect 570848 643098 570880 643334
rect 570260 643066 570880 643098
rect 585310 643654 585930 683098
rect 585310 643418 585342 643654
rect 585578 643418 585662 643654
rect 585898 643418 585930 643654
rect 585310 643334 585930 643418
rect 585310 643098 585342 643334
rect 585578 643098 585662 643334
rect 585898 643098 585930 643334
rect 7844 623654 8464 623686
rect 7844 623418 7876 623654
rect 8112 623418 8196 623654
rect 8432 623418 8464 623654
rect 7844 623334 8464 623418
rect 7844 623098 7876 623334
rect 8112 623098 8196 623334
rect 8432 623098 8464 623334
rect 7844 623066 8464 623098
rect 38000 623654 38620 623686
rect 38000 623418 38032 623654
rect 38268 623418 38352 623654
rect 38588 623418 38620 623654
rect 38000 623334 38620 623418
rect 38000 623098 38032 623334
rect 38268 623098 38352 623334
rect 38588 623098 38620 623334
rect 38000 623066 38620 623098
rect 74000 623654 74620 623686
rect 74000 623418 74032 623654
rect 74268 623418 74352 623654
rect 74588 623418 74620 623654
rect 74000 623334 74620 623418
rect 74000 623098 74032 623334
rect 74268 623098 74352 623334
rect 74588 623098 74620 623334
rect 74000 623066 74620 623098
rect 110000 623654 110620 623686
rect 110000 623418 110032 623654
rect 110268 623418 110352 623654
rect 110588 623418 110620 623654
rect 110000 623334 110620 623418
rect 110000 623098 110032 623334
rect 110268 623098 110352 623334
rect 110588 623098 110620 623334
rect 110000 623066 110620 623098
rect 146000 623654 146620 623686
rect 146000 623418 146032 623654
rect 146268 623418 146352 623654
rect 146588 623418 146620 623654
rect 146000 623334 146620 623418
rect 146000 623098 146032 623334
rect 146268 623098 146352 623334
rect 146588 623098 146620 623334
rect 146000 623066 146620 623098
rect 182000 623654 182620 623686
rect 182000 623418 182032 623654
rect 182268 623418 182352 623654
rect 182588 623418 182620 623654
rect 182000 623334 182620 623418
rect 182000 623098 182032 623334
rect 182268 623098 182352 623334
rect 182588 623098 182620 623334
rect 182000 623066 182620 623098
rect 218000 623654 218620 623686
rect 218000 623418 218032 623654
rect 218268 623418 218352 623654
rect 218588 623418 218620 623654
rect 218000 623334 218620 623418
rect 218000 623098 218032 623334
rect 218268 623098 218352 623334
rect 218588 623098 218620 623334
rect 218000 623066 218620 623098
rect 254000 623654 254620 623686
rect 254000 623418 254032 623654
rect 254268 623418 254352 623654
rect 254588 623418 254620 623654
rect 254000 623334 254620 623418
rect 254000 623098 254032 623334
rect 254268 623098 254352 623334
rect 254588 623098 254620 623334
rect 254000 623066 254620 623098
rect 290000 623654 290620 623686
rect 290000 623418 290032 623654
rect 290268 623418 290352 623654
rect 290588 623418 290620 623654
rect 290000 623334 290620 623418
rect 290000 623098 290032 623334
rect 290268 623098 290352 623334
rect 290588 623098 290620 623334
rect 290000 623066 290620 623098
rect 326000 623654 326620 623686
rect 326000 623418 326032 623654
rect 326268 623418 326352 623654
rect 326588 623418 326620 623654
rect 326000 623334 326620 623418
rect 326000 623098 326032 623334
rect 326268 623098 326352 623334
rect 326588 623098 326620 623334
rect 326000 623066 326620 623098
rect 362000 623654 362620 623686
rect 362000 623418 362032 623654
rect 362268 623418 362352 623654
rect 362588 623418 362620 623654
rect 362000 623334 362620 623418
rect 362000 623098 362032 623334
rect 362268 623098 362352 623334
rect 362588 623098 362620 623334
rect 362000 623066 362620 623098
rect 398000 623654 398620 623686
rect 398000 623418 398032 623654
rect 398268 623418 398352 623654
rect 398588 623418 398620 623654
rect 398000 623334 398620 623418
rect 398000 623098 398032 623334
rect 398268 623098 398352 623334
rect 398588 623098 398620 623334
rect 398000 623066 398620 623098
rect 434000 623654 434620 623686
rect 434000 623418 434032 623654
rect 434268 623418 434352 623654
rect 434588 623418 434620 623654
rect 434000 623334 434620 623418
rect 434000 623098 434032 623334
rect 434268 623098 434352 623334
rect 434588 623098 434620 623334
rect 434000 623066 434620 623098
rect 470000 623654 470620 623686
rect 470000 623418 470032 623654
rect 470268 623418 470352 623654
rect 470588 623418 470620 623654
rect 470000 623334 470620 623418
rect 470000 623098 470032 623334
rect 470268 623098 470352 623334
rect 470588 623098 470620 623334
rect 470000 623066 470620 623098
rect 506000 623654 506620 623686
rect 506000 623418 506032 623654
rect 506268 623418 506352 623654
rect 506588 623418 506620 623654
rect 506000 623334 506620 623418
rect 506000 623098 506032 623334
rect 506268 623098 506352 623334
rect 506588 623098 506620 623334
rect 506000 623066 506620 623098
rect 542000 623654 542620 623686
rect 542000 623418 542032 623654
rect 542268 623418 542352 623654
rect 542588 623418 542620 623654
rect 542000 623334 542620 623418
rect 542000 623098 542032 623334
rect 542268 623098 542352 623334
rect 542588 623098 542620 623334
rect 542000 623066 542620 623098
rect 571500 623654 572120 623686
rect 571500 623418 571532 623654
rect 571768 623418 571852 623654
rect 572088 623418 572120 623654
rect 571500 623334 572120 623418
rect 571500 623098 571532 623334
rect 571768 623098 571852 623334
rect 572088 623098 572120 623334
rect 571500 623066 572120 623098
rect -2006 603418 -1974 603654
rect -1738 603418 -1654 603654
rect -1418 603418 -1386 603654
rect -2006 603334 -1386 603418
rect -2006 603098 -1974 603334
rect -1738 603098 -1654 603334
rect -1418 603098 -1386 603334
rect -2006 563654 -1386 603098
rect 9084 603654 9704 603686
rect 9084 603418 9116 603654
rect 9352 603418 9436 603654
rect 9672 603418 9704 603654
rect 9084 603334 9704 603418
rect 9084 603098 9116 603334
rect 9352 603098 9436 603334
rect 9672 603098 9704 603334
rect 9084 603066 9704 603098
rect 56620 603654 57240 603686
rect 56620 603418 56652 603654
rect 56888 603418 56972 603654
rect 57208 603418 57240 603654
rect 56620 603334 57240 603418
rect 56620 603098 56652 603334
rect 56888 603098 56972 603334
rect 57208 603098 57240 603334
rect 56620 603066 57240 603098
rect 92620 603654 93240 603686
rect 92620 603418 92652 603654
rect 92888 603418 92972 603654
rect 93208 603418 93240 603654
rect 92620 603334 93240 603418
rect 92620 603098 92652 603334
rect 92888 603098 92972 603334
rect 93208 603098 93240 603334
rect 92620 603066 93240 603098
rect 128620 603654 129240 603686
rect 128620 603418 128652 603654
rect 128888 603418 128972 603654
rect 129208 603418 129240 603654
rect 128620 603334 129240 603418
rect 128620 603098 128652 603334
rect 128888 603098 128972 603334
rect 129208 603098 129240 603334
rect 128620 603066 129240 603098
rect 164620 603654 165240 603686
rect 164620 603418 164652 603654
rect 164888 603418 164972 603654
rect 165208 603418 165240 603654
rect 164620 603334 165240 603418
rect 164620 603098 164652 603334
rect 164888 603098 164972 603334
rect 165208 603098 165240 603334
rect 164620 603066 165240 603098
rect 200620 603654 201240 603686
rect 200620 603418 200652 603654
rect 200888 603418 200972 603654
rect 201208 603418 201240 603654
rect 200620 603334 201240 603418
rect 200620 603098 200652 603334
rect 200888 603098 200972 603334
rect 201208 603098 201240 603334
rect 200620 603066 201240 603098
rect 236620 603654 237240 603686
rect 236620 603418 236652 603654
rect 236888 603418 236972 603654
rect 237208 603418 237240 603654
rect 236620 603334 237240 603418
rect 236620 603098 236652 603334
rect 236888 603098 236972 603334
rect 237208 603098 237240 603334
rect 236620 603066 237240 603098
rect 272620 603654 273240 603686
rect 272620 603418 272652 603654
rect 272888 603418 272972 603654
rect 273208 603418 273240 603654
rect 272620 603334 273240 603418
rect 272620 603098 272652 603334
rect 272888 603098 272972 603334
rect 273208 603098 273240 603334
rect 272620 603066 273240 603098
rect 308620 603654 309240 603686
rect 308620 603418 308652 603654
rect 308888 603418 308972 603654
rect 309208 603418 309240 603654
rect 308620 603334 309240 603418
rect 308620 603098 308652 603334
rect 308888 603098 308972 603334
rect 309208 603098 309240 603334
rect 308620 603066 309240 603098
rect 344620 603654 345240 603686
rect 344620 603418 344652 603654
rect 344888 603418 344972 603654
rect 345208 603418 345240 603654
rect 344620 603334 345240 603418
rect 344620 603098 344652 603334
rect 344888 603098 344972 603334
rect 345208 603098 345240 603334
rect 344620 603066 345240 603098
rect 380620 603654 381240 603686
rect 380620 603418 380652 603654
rect 380888 603418 380972 603654
rect 381208 603418 381240 603654
rect 380620 603334 381240 603418
rect 380620 603098 380652 603334
rect 380888 603098 380972 603334
rect 381208 603098 381240 603334
rect 380620 603066 381240 603098
rect 416620 603654 417240 603686
rect 416620 603418 416652 603654
rect 416888 603418 416972 603654
rect 417208 603418 417240 603654
rect 416620 603334 417240 603418
rect 416620 603098 416652 603334
rect 416888 603098 416972 603334
rect 417208 603098 417240 603334
rect 416620 603066 417240 603098
rect 452620 603654 453240 603686
rect 452620 603418 452652 603654
rect 452888 603418 452972 603654
rect 453208 603418 453240 603654
rect 452620 603334 453240 603418
rect 452620 603098 452652 603334
rect 452888 603098 452972 603334
rect 453208 603098 453240 603334
rect 452620 603066 453240 603098
rect 488620 603654 489240 603686
rect 488620 603418 488652 603654
rect 488888 603418 488972 603654
rect 489208 603418 489240 603654
rect 488620 603334 489240 603418
rect 488620 603098 488652 603334
rect 488888 603098 488972 603334
rect 489208 603098 489240 603334
rect 488620 603066 489240 603098
rect 524620 603654 525240 603686
rect 524620 603418 524652 603654
rect 524888 603418 524972 603654
rect 525208 603418 525240 603654
rect 524620 603334 525240 603418
rect 524620 603098 524652 603334
rect 524888 603098 524972 603334
rect 525208 603098 525240 603334
rect 524620 603066 525240 603098
rect 560620 603654 561240 603686
rect 560620 603418 560652 603654
rect 560888 603418 560972 603654
rect 561208 603418 561240 603654
rect 560620 603334 561240 603418
rect 560620 603098 560652 603334
rect 560888 603098 560972 603334
rect 561208 603098 561240 603334
rect 560620 603066 561240 603098
rect 570260 603654 570880 603686
rect 570260 603418 570292 603654
rect 570528 603418 570612 603654
rect 570848 603418 570880 603654
rect 570260 603334 570880 603418
rect 570260 603098 570292 603334
rect 570528 603098 570612 603334
rect 570848 603098 570880 603334
rect 570260 603066 570880 603098
rect 585310 603654 585930 643098
rect 585310 603418 585342 603654
rect 585578 603418 585662 603654
rect 585898 603418 585930 603654
rect 585310 603334 585930 603418
rect 585310 603098 585342 603334
rect 585578 603098 585662 603334
rect 585898 603098 585930 603334
rect 7844 583654 8464 583686
rect 7844 583418 7876 583654
rect 8112 583418 8196 583654
rect 8432 583418 8464 583654
rect 7844 583334 8464 583418
rect 7844 583098 7876 583334
rect 8112 583098 8196 583334
rect 8432 583098 8464 583334
rect 7844 583066 8464 583098
rect 38000 583654 38620 583686
rect 38000 583418 38032 583654
rect 38268 583418 38352 583654
rect 38588 583418 38620 583654
rect 38000 583334 38620 583418
rect 38000 583098 38032 583334
rect 38268 583098 38352 583334
rect 38588 583098 38620 583334
rect 38000 583066 38620 583098
rect 74000 583654 74620 583686
rect 74000 583418 74032 583654
rect 74268 583418 74352 583654
rect 74588 583418 74620 583654
rect 74000 583334 74620 583418
rect 74000 583098 74032 583334
rect 74268 583098 74352 583334
rect 74588 583098 74620 583334
rect 74000 583066 74620 583098
rect 110000 583654 110620 583686
rect 110000 583418 110032 583654
rect 110268 583418 110352 583654
rect 110588 583418 110620 583654
rect 110000 583334 110620 583418
rect 110000 583098 110032 583334
rect 110268 583098 110352 583334
rect 110588 583098 110620 583334
rect 110000 583066 110620 583098
rect 146000 583654 146620 583686
rect 146000 583418 146032 583654
rect 146268 583418 146352 583654
rect 146588 583418 146620 583654
rect 146000 583334 146620 583418
rect 146000 583098 146032 583334
rect 146268 583098 146352 583334
rect 146588 583098 146620 583334
rect 146000 583066 146620 583098
rect 182000 583654 182620 583686
rect 182000 583418 182032 583654
rect 182268 583418 182352 583654
rect 182588 583418 182620 583654
rect 182000 583334 182620 583418
rect 182000 583098 182032 583334
rect 182268 583098 182352 583334
rect 182588 583098 182620 583334
rect 182000 583066 182620 583098
rect 218000 583654 218620 583686
rect 218000 583418 218032 583654
rect 218268 583418 218352 583654
rect 218588 583418 218620 583654
rect 218000 583334 218620 583418
rect 218000 583098 218032 583334
rect 218268 583098 218352 583334
rect 218588 583098 218620 583334
rect 218000 583066 218620 583098
rect 254000 583654 254620 583686
rect 254000 583418 254032 583654
rect 254268 583418 254352 583654
rect 254588 583418 254620 583654
rect 254000 583334 254620 583418
rect 254000 583098 254032 583334
rect 254268 583098 254352 583334
rect 254588 583098 254620 583334
rect 254000 583066 254620 583098
rect 290000 583654 290620 583686
rect 290000 583418 290032 583654
rect 290268 583418 290352 583654
rect 290588 583418 290620 583654
rect 290000 583334 290620 583418
rect 290000 583098 290032 583334
rect 290268 583098 290352 583334
rect 290588 583098 290620 583334
rect 290000 583066 290620 583098
rect 326000 583654 326620 583686
rect 326000 583418 326032 583654
rect 326268 583418 326352 583654
rect 326588 583418 326620 583654
rect 326000 583334 326620 583418
rect 326000 583098 326032 583334
rect 326268 583098 326352 583334
rect 326588 583098 326620 583334
rect 326000 583066 326620 583098
rect 362000 583654 362620 583686
rect 362000 583418 362032 583654
rect 362268 583418 362352 583654
rect 362588 583418 362620 583654
rect 362000 583334 362620 583418
rect 362000 583098 362032 583334
rect 362268 583098 362352 583334
rect 362588 583098 362620 583334
rect 362000 583066 362620 583098
rect 398000 583654 398620 583686
rect 398000 583418 398032 583654
rect 398268 583418 398352 583654
rect 398588 583418 398620 583654
rect 398000 583334 398620 583418
rect 398000 583098 398032 583334
rect 398268 583098 398352 583334
rect 398588 583098 398620 583334
rect 398000 583066 398620 583098
rect 434000 583654 434620 583686
rect 434000 583418 434032 583654
rect 434268 583418 434352 583654
rect 434588 583418 434620 583654
rect 434000 583334 434620 583418
rect 434000 583098 434032 583334
rect 434268 583098 434352 583334
rect 434588 583098 434620 583334
rect 434000 583066 434620 583098
rect 470000 583654 470620 583686
rect 470000 583418 470032 583654
rect 470268 583418 470352 583654
rect 470588 583418 470620 583654
rect 470000 583334 470620 583418
rect 470000 583098 470032 583334
rect 470268 583098 470352 583334
rect 470588 583098 470620 583334
rect 470000 583066 470620 583098
rect 506000 583654 506620 583686
rect 506000 583418 506032 583654
rect 506268 583418 506352 583654
rect 506588 583418 506620 583654
rect 506000 583334 506620 583418
rect 506000 583098 506032 583334
rect 506268 583098 506352 583334
rect 506588 583098 506620 583334
rect 506000 583066 506620 583098
rect 542000 583654 542620 583686
rect 542000 583418 542032 583654
rect 542268 583418 542352 583654
rect 542588 583418 542620 583654
rect 542000 583334 542620 583418
rect 542000 583098 542032 583334
rect 542268 583098 542352 583334
rect 542588 583098 542620 583334
rect 542000 583066 542620 583098
rect 571500 583654 572120 583686
rect 571500 583418 571532 583654
rect 571768 583418 571852 583654
rect 572088 583418 572120 583654
rect 571500 583334 572120 583418
rect 571500 583098 571532 583334
rect 571768 583098 571852 583334
rect 572088 583098 572120 583334
rect 571500 583066 572120 583098
rect -2006 563418 -1974 563654
rect -1738 563418 -1654 563654
rect -1418 563418 -1386 563654
rect -2006 563334 -1386 563418
rect -2006 563098 -1974 563334
rect -1738 563098 -1654 563334
rect -1418 563098 -1386 563334
rect -2006 523654 -1386 563098
rect 9084 563654 9704 563686
rect 9084 563418 9116 563654
rect 9352 563418 9436 563654
rect 9672 563418 9704 563654
rect 9084 563334 9704 563418
rect 9084 563098 9116 563334
rect 9352 563098 9436 563334
rect 9672 563098 9704 563334
rect 9084 563066 9704 563098
rect 56620 563654 57240 563686
rect 56620 563418 56652 563654
rect 56888 563418 56972 563654
rect 57208 563418 57240 563654
rect 56620 563334 57240 563418
rect 56620 563098 56652 563334
rect 56888 563098 56972 563334
rect 57208 563098 57240 563334
rect 56620 563066 57240 563098
rect 92620 563654 93240 563686
rect 92620 563418 92652 563654
rect 92888 563418 92972 563654
rect 93208 563418 93240 563654
rect 92620 563334 93240 563418
rect 92620 563098 92652 563334
rect 92888 563098 92972 563334
rect 93208 563098 93240 563334
rect 92620 563066 93240 563098
rect 128620 563654 129240 563686
rect 128620 563418 128652 563654
rect 128888 563418 128972 563654
rect 129208 563418 129240 563654
rect 128620 563334 129240 563418
rect 128620 563098 128652 563334
rect 128888 563098 128972 563334
rect 129208 563098 129240 563334
rect 128620 563066 129240 563098
rect 164620 563654 165240 563686
rect 164620 563418 164652 563654
rect 164888 563418 164972 563654
rect 165208 563418 165240 563654
rect 164620 563334 165240 563418
rect 164620 563098 164652 563334
rect 164888 563098 164972 563334
rect 165208 563098 165240 563334
rect 164620 563066 165240 563098
rect 200620 563654 201240 563686
rect 200620 563418 200652 563654
rect 200888 563418 200972 563654
rect 201208 563418 201240 563654
rect 200620 563334 201240 563418
rect 200620 563098 200652 563334
rect 200888 563098 200972 563334
rect 201208 563098 201240 563334
rect 200620 563066 201240 563098
rect 236620 563654 237240 563686
rect 236620 563418 236652 563654
rect 236888 563418 236972 563654
rect 237208 563418 237240 563654
rect 236620 563334 237240 563418
rect 236620 563098 236652 563334
rect 236888 563098 236972 563334
rect 237208 563098 237240 563334
rect 236620 563066 237240 563098
rect 272620 563654 273240 563686
rect 272620 563418 272652 563654
rect 272888 563418 272972 563654
rect 273208 563418 273240 563654
rect 272620 563334 273240 563418
rect 272620 563098 272652 563334
rect 272888 563098 272972 563334
rect 273208 563098 273240 563334
rect 272620 563066 273240 563098
rect 308620 563654 309240 563686
rect 308620 563418 308652 563654
rect 308888 563418 308972 563654
rect 309208 563418 309240 563654
rect 308620 563334 309240 563418
rect 308620 563098 308652 563334
rect 308888 563098 308972 563334
rect 309208 563098 309240 563334
rect 308620 563066 309240 563098
rect 344620 563654 345240 563686
rect 344620 563418 344652 563654
rect 344888 563418 344972 563654
rect 345208 563418 345240 563654
rect 344620 563334 345240 563418
rect 344620 563098 344652 563334
rect 344888 563098 344972 563334
rect 345208 563098 345240 563334
rect 344620 563066 345240 563098
rect 380620 563654 381240 563686
rect 380620 563418 380652 563654
rect 380888 563418 380972 563654
rect 381208 563418 381240 563654
rect 380620 563334 381240 563418
rect 380620 563098 380652 563334
rect 380888 563098 380972 563334
rect 381208 563098 381240 563334
rect 380620 563066 381240 563098
rect 416620 563654 417240 563686
rect 416620 563418 416652 563654
rect 416888 563418 416972 563654
rect 417208 563418 417240 563654
rect 416620 563334 417240 563418
rect 416620 563098 416652 563334
rect 416888 563098 416972 563334
rect 417208 563098 417240 563334
rect 416620 563066 417240 563098
rect 452620 563654 453240 563686
rect 452620 563418 452652 563654
rect 452888 563418 452972 563654
rect 453208 563418 453240 563654
rect 452620 563334 453240 563418
rect 452620 563098 452652 563334
rect 452888 563098 452972 563334
rect 453208 563098 453240 563334
rect 452620 563066 453240 563098
rect 488620 563654 489240 563686
rect 488620 563418 488652 563654
rect 488888 563418 488972 563654
rect 489208 563418 489240 563654
rect 488620 563334 489240 563418
rect 488620 563098 488652 563334
rect 488888 563098 488972 563334
rect 489208 563098 489240 563334
rect 488620 563066 489240 563098
rect 524620 563654 525240 563686
rect 524620 563418 524652 563654
rect 524888 563418 524972 563654
rect 525208 563418 525240 563654
rect 524620 563334 525240 563418
rect 524620 563098 524652 563334
rect 524888 563098 524972 563334
rect 525208 563098 525240 563334
rect 524620 563066 525240 563098
rect 560620 563654 561240 563686
rect 560620 563418 560652 563654
rect 560888 563418 560972 563654
rect 561208 563418 561240 563654
rect 560620 563334 561240 563418
rect 560620 563098 560652 563334
rect 560888 563098 560972 563334
rect 561208 563098 561240 563334
rect 560620 563066 561240 563098
rect 570260 563654 570880 563686
rect 570260 563418 570292 563654
rect 570528 563418 570612 563654
rect 570848 563418 570880 563654
rect 570260 563334 570880 563418
rect 570260 563098 570292 563334
rect 570528 563098 570612 563334
rect 570848 563098 570880 563334
rect 570260 563066 570880 563098
rect 585310 563654 585930 603098
rect 585310 563418 585342 563654
rect 585578 563418 585662 563654
rect 585898 563418 585930 563654
rect 585310 563334 585930 563418
rect 585310 563098 585342 563334
rect 585578 563098 585662 563334
rect 585898 563098 585930 563334
rect 7844 543654 8464 543686
rect 7844 543418 7876 543654
rect 8112 543418 8196 543654
rect 8432 543418 8464 543654
rect 7844 543334 8464 543418
rect 7844 543098 7876 543334
rect 8112 543098 8196 543334
rect 8432 543098 8464 543334
rect 7844 543066 8464 543098
rect 38000 543654 38620 543686
rect 38000 543418 38032 543654
rect 38268 543418 38352 543654
rect 38588 543418 38620 543654
rect 38000 543334 38620 543418
rect 38000 543098 38032 543334
rect 38268 543098 38352 543334
rect 38588 543098 38620 543334
rect 38000 543066 38620 543098
rect 74000 543654 74620 543686
rect 74000 543418 74032 543654
rect 74268 543418 74352 543654
rect 74588 543418 74620 543654
rect 74000 543334 74620 543418
rect 74000 543098 74032 543334
rect 74268 543098 74352 543334
rect 74588 543098 74620 543334
rect 74000 543066 74620 543098
rect 110000 543654 110620 543686
rect 110000 543418 110032 543654
rect 110268 543418 110352 543654
rect 110588 543418 110620 543654
rect 110000 543334 110620 543418
rect 110000 543098 110032 543334
rect 110268 543098 110352 543334
rect 110588 543098 110620 543334
rect 110000 543066 110620 543098
rect 146000 543654 146620 543686
rect 146000 543418 146032 543654
rect 146268 543418 146352 543654
rect 146588 543418 146620 543654
rect 146000 543334 146620 543418
rect 146000 543098 146032 543334
rect 146268 543098 146352 543334
rect 146588 543098 146620 543334
rect 146000 543066 146620 543098
rect 182000 543654 182620 543686
rect 182000 543418 182032 543654
rect 182268 543418 182352 543654
rect 182588 543418 182620 543654
rect 182000 543334 182620 543418
rect 182000 543098 182032 543334
rect 182268 543098 182352 543334
rect 182588 543098 182620 543334
rect 182000 543066 182620 543098
rect 218000 543654 218620 543686
rect 218000 543418 218032 543654
rect 218268 543418 218352 543654
rect 218588 543418 218620 543654
rect 218000 543334 218620 543418
rect 218000 543098 218032 543334
rect 218268 543098 218352 543334
rect 218588 543098 218620 543334
rect 218000 543066 218620 543098
rect 254000 543654 254620 543686
rect 254000 543418 254032 543654
rect 254268 543418 254352 543654
rect 254588 543418 254620 543654
rect 254000 543334 254620 543418
rect 254000 543098 254032 543334
rect 254268 543098 254352 543334
rect 254588 543098 254620 543334
rect 254000 543066 254620 543098
rect 290000 543654 290620 543686
rect 290000 543418 290032 543654
rect 290268 543418 290352 543654
rect 290588 543418 290620 543654
rect 290000 543334 290620 543418
rect 290000 543098 290032 543334
rect 290268 543098 290352 543334
rect 290588 543098 290620 543334
rect 290000 543066 290620 543098
rect 326000 543654 326620 543686
rect 326000 543418 326032 543654
rect 326268 543418 326352 543654
rect 326588 543418 326620 543654
rect 326000 543334 326620 543418
rect 326000 543098 326032 543334
rect 326268 543098 326352 543334
rect 326588 543098 326620 543334
rect 326000 543066 326620 543098
rect 362000 543654 362620 543686
rect 362000 543418 362032 543654
rect 362268 543418 362352 543654
rect 362588 543418 362620 543654
rect 362000 543334 362620 543418
rect 362000 543098 362032 543334
rect 362268 543098 362352 543334
rect 362588 543098 362620 543334
rect 362000 543066 362620 543098
rect 398000 543654 398620 543686
rect 398000 543418 398032 543654
rect 398268 543418 398352 543654
rect 398588 543418 398620 543654
rect 398000 543334 398620 543418
rect 398000 543098 398032 543334
rect 398268 543098 398352 543334
rect 398588 543098 398620 543334
rect 398000 543066 398620 543098
rect 434000 543654 434620 543686
rect 434000 543418 434032 543654
rect 434268 543418 434352 543654
rect 434588 543418 434620 543654
rect 434000 543334 434620 543418
rect 434000 543098 434032 543334
rect 434268 543098 434352 543334
rect 434588 543098 434620 543334
rect 434000 543066 434620 543098
rect 470000 543654 470620 543686
rect 470000 543418 470032 543654
rect 470268 543418 470352 543654
rect 470588 543418 470620 543654
rect 470000 543334 470620 543418
rect 470000 543098 470032 543334
rect 470268 543098 470352 543334
rect 470588 543098 470620 543334
rect 470000 543066 470620 543098
rect 506000 543654 506620 543686
rect 506000 543418 506032 543654
rect 506268 543418 506352 543654
rect 506588 543418 506620 543654
rect 506000 543334 506620 543418
rect 506000 543098 506032 543334
rect 506268 543098 506352 543334
rect 506588 543098 506620 543334
rect 506000 543066 506620 543098
rect 542000 543654 542620 543686
rect 542000 543418 542032 543654
rect 542268 543418 542352 543654
rect 542588 543418 542620 543654
rect 542000 543334 542620 543418
rect 542000 543098 542032 543334
rect 542268 543098 542352 543334
rect 542588 543098 542620 543334
rect 542000 543066 542620 543098
rect 571500 543654 572120 543686
rect 571500 543418 571532 543654
rect 571768 543418 571852 543654
rect 572088 543418 572120 543654
rect 571500 543334 572120 543418
rect 571500 543098 571532 543334
rect 571768 543098 571852 543334
rect 572088 543098 572120 543334
rect 571500 543066 572120 543098
rect -2006 523418 -1974 523654
rect -1738 523418 -1654 523654
rect -1418 523418 -1386 523654
rect -2006 523334 -1386 523418
rect -2006 523098 -1974 523334
rect -1738 523098 -1654 523334
rect -1418 523098 -1386 523334
rect -2006 483654 -1386 523098
rect 9084 523654 9704 523686
rect 9084 523418 9116 523654
rect 9352 523418 9436 523654
rect 9672 523418 9704 523654
rect 9084 523334 9704 523418
rect 9084 523098 9116 523334
rect 9352 523098 9436 523334
rect 9672 523098 9704 523334
rect 9084 523066 9704 523098
rect 56620 523654 57240 523686
rect 56620 523418 56652 523654
rect 56888 523418 56972 523654
rect 57208 523418 57240 523654
rect 56620 523334 57240 523418
rect 56620 523098 56652 523334
rect 56888 523098 56972 523334
rect 57208 523098 57240 523334
rect 56620 523066 57240 523098
rect 92620 523654 93240 523686
rect 92620 523418 92652 523654
rect 92888 523418 92972 523654
rect 93208 523418 93240 523654
rect 92620 523334 93240 523418
rect 92620 523098 92652 523334
rect 92888 523098 92972 523334
rect 93208 523098 93240 523334
rect 92620 523066 93240 523098
rect 128620 523654 129240 523686
rect 128620 523418 128652 523654
rect 128888 523418 128972 523654
rect 129208 523418 129240 523654
rect 128620 523334 129240 523418
rect 128620 523098 128652 523334
rect 128888 523098 128972 523334
rect 129208 523098 129240 523334
rect 128620 523066 129240 523098
rect 164620 523654 165240 523686
rect 164620 523418 164652 523654
rect 164888 523418 164972 523654
rect 165208 523418 165240 523654
rect 164620 523334 165240 523418
rect 164620 523098 164652 523334
rect 164888 523098 164972 523334
rect 165208 523098 165240 523334
rect 164620 523066 165240 523098
rect 200620 523654 201240 523686
rect 200620 523418 200652 523654
rect 200888 523418 200972 523654
rect 201208 523418 201240 523654
rect 200620 523334 201240 523418
rect 200620 523098 200652 523334
rect 200888 523098 200972 523334
rect 201208 523098 201240 523334
rect 200620 523066 201240 523098
rect 236620 523654 237240 523686
rect 236620 523418 236652 523654
rect 236888 523418 236972 523654
rect 237208 523418 237240 523654
rect 236620 523334 237240 523418
rect 236620 523098 236652 523334
rect 236888 523098 236972 523334
rect 237208 523098 237240 523334
rect 236620 523066 237240 523098
rect 272620 523654 273240 523686
rect 272620 523418 272652 523654
rect 272888 523418 272972 523654
rect 273208 523418 273240 523654
rect 272620 523334 273240 523418
rect 272620 523098 272652 523334
rect 272888 523098 272972 523334
rect 273208 523098 273240 523334
rect 272620 523066 273240 523098
rect 308620 523654 309240 523686
rect 308620 523418 308652 523654
rect 308888 523418 308972 523654
rect 309208 523418 309240 523654
rect 308620 523334 309240 523418
rect 308620 523098 308652 523334
rect 308888 523098 308972 523334
rect 309208 523098 309240 523334
rect 308620 523066 309240 523098
rect 344620 523654 345240 523686
rect 344620 523418 344652 523654
rect 344888 523418 344972 523654
rect 345208 523418 345240 523654
rect 344620 523334 345240 523418
rect 344620 523098 344652 523334
rect 344888 523098 344972 523334
rect 345208 523098 345240 523334
rect 344620 523066 345240 523098
rect 380620 523654 381240 523686
rect 380620 523418 380652 523654
rect 380888 523418 380972 523654
rect 381208 523418 381240 523654
rect 380620 523334 381240 523418
rect 380620 523098 380652 523334
rect 380888 523098 380972 523334
rect 381208 523098 381240 523334
rect 380620 523066 381240 523098
rect 416620 523654 417240 523686
rect 416620 523418 416652 523654
rect 416888 523418 416972 523654
rect 417208 523418 417240 523654
rect 416620 523334 417240 523418
rect 416620 523098 416652 523334
rect 416888 523098 416972 523334
rect 417208 523098 417240 523334
rect 416620 523066 417240 523098
rect 452620 523654 453240 523686
rect 452620 523418 452652 523654
rect 452888 523418 452972 523654
rect 453208 523418 453240 523654
rect 452620 523334 453240 523418
rect 452620 523098 452652 523334
rect 452888 523098 452972 523334
rect 453208 523098 453240 523334
rect 452620 523066 453240 523098
rect 488620 523654 489240 523686
rect 488620 523418 488652 523654
rect 488888 523418 488972 523654
rect 489208 523418 489240 523654
rect 488620 523334 489240 523418
rect 488620 523098 488652 523334
rect 488888 523098 488972 523334
rect 489208 523098 489240 523334
rect 488620 523066 489240 523098
rect 524620 523654 525240 523686
rect 524620 523418 524652 523654
rect 524888 523418 524972 523654
rect 525208 523418 525240 523654
rect 524620 523334 525240 523418
rect 524620 523098 524652 523334
rect 524888 523098 524972 523334
rect 525208 523098 525240 523334
rect 524620 523066 525240 523098
rect 560620 523654 561240 523686
rect 560620 523418 560652 523654
rect 560888 523418 560972 523654
rect 561208 523418 561240 523654
rect 560620 523334 561240 523418
rect 560620 523098 560652 523334
rect 560888 523098 560972 523334
rect 561208 523098 561240 523334
rect 560620 523066 561240 523098
rect 570260 523654 570880 523686
rect 570260 523418 570292 523654
rect 570528 523418 570612 523654
rect 570848 523418 570880 523654
rect 570260 523334 570880 523418
rect 570260 523098 570292 523334
rect 570528 523098 570612 523334
rect 570848 523098 570880 523334
rect 570260 523066 570880 523098
rect 585310 523654 585930 563098
rect 585310 523418 585342 523654
rect 585578 523418 585662 523654
rect 585898 523418 585930 523654
rect 585310 523334 585930 523418
rect 585310 523098 585342 523334
rect 585578 523098 585662 523334
rect 585898 523098 585930 523334
rect 7844 503654 8464 503686
rect 7844 503418 7876 503654
rect 8112 503418 8196 503654
rect 8432 503418 8464 503654
rect 7844 503334 8464 503418
rect 7844 503098 7876 503334
rect 8112 503098 8196 503334
rect 8432 503098 8464 503334
rect 7844 503066 8464 503098
rect 38000 503654 38620 503686
rect 38000 503418 38032 503654
rect 38268 503418 38352 503654
rect 38588 503418 38620 503654
rect 38000 503334 38620 503418
rect 38000 503098 38032 503334
rect 38268 503098 38352 503334
rect 38588 503098 38620 503334
rect 38000 503066 38620 503098
rect 60560 503654 60920 503686
rect 60560 503418 60622 503654
rect 60858 503418 60920 503654
rect 60560 503334 60920 503418
rect 60560 503098 60622 503334
rect 60858 503098 60920 503334
rect 60560 503066 60920 503098
rect 159036 503654 159396 503686
rect 159036 503418 159098 503654
rect 159334 503418 159396 503654
rect 159036 503334 159396 503418
rect 159036 503098 159098 503334
rect 159334 503098 159396 503334
rect 159036 503066 159396 503098
rect 182000 503654 182620 503686
rect 182000 503418 182032 503654
rect 182268 503418 182352 503654
rect 182588 503418 182620 503654
rect 182000 503334 182620 503418
rect 182000 503098 182032 503334
rect 182268 503098 182352 503334
rect 182588 503098 182620 503334
rect 182000 503066 182620 503098
rect 185560 503654 185920 503686
rect 185560 503418 185622 503654
rect 185858 503418 185920 503654
rect 185560 503334 185920 503418
rect 185560 503098 185622 503334
rect 185858 503098 185920 503334
rect 185560 503066 185920 503098
rect 284036 503654 284396 503686
rect 284036 503418 284098 503654
rect 284334 503418 284396 503654
rect 284036 503334 284396 503418
rect 284036 503098 284098 503334
rect 284334 503098 284396 503334
rect 284036 503066 284396 503098
rect 290000 503654 290620 503686
rect 290000 503418 290032 503654
rect 290268 503418 290352 503654
rect 290588 503418 290620 503654
rect 290000 503334 290620 503418
rect 290000 503098 290032 503334
rect 290268 503098 290352 503334
rect 290588 503098 290620 503334
rect 290000 503066 290620 503098
rect 310560 503654 310920 503686
rect 310560 503418 310622 503654
rect 310858 503418 310920 503654
rect 310560 503334 310920 503418
rect 310560 503098 310622 503334
rect 310858 503098 310920 503334
rect 310560 503066 310920 503098
rect 409036 503654 409396 503686
rect 409036 503418 409098 503654
rect 409334 503418 409396 503654
rect 409036 503334 409396 503418
rect 409036 503098 409098 503334
rect 409334 503098 409396 503334
rect 409036 503066 409396 503098
rect 434000 503654 434620 503686
rect 434000 503418 434032 503654
rect 434268 503418 434352 503654
rect 434588 503418 434620 503654
rect 434000 503334 434620 503418
rect 434000 503098 434032 503334
rect 434268 503098 434352 503334
rect 434588 503098 434620 503334
rect 434000 503066 434620 503098
rect 436560 503654 436920 503686
rect 436560 503418 436622 503654
rect 436858 503418 436920 503654
rect 436560 503334 436920 503418
rect 436560 503098 436622 503334
rect 436858 503098 436920 503334
rect 436560 503066 436920 503098
rect 535036 503654 535396 503686
rect 535036 503418 535098 503654
rect 535334 503418 535396 503654
rect 535036 503334 535396 503418
rect 535036 503098 535098 503334
rect 535334 503098 535396 503334
rect 535036 503066 535396 503098
rect 542000 503654 542620 503686
rect 542000 503418 542032 503654
rect 542268 503418 542352 503654
rect 542588 503418 542620 503654
rect 542000 503334 542620 503418
rect 542000 503098 542032 503334
rect 542268 503098 542352 503334
rect 542588 503098 542620 503334
rect 542000 503066 542620 503098
rect 571500 503654 572120 503686
rect 571500 503418 571532 503654
rect 571768 503418 571852 503654
rect 572088 503418 572120 503654
rect 571500 503334 572120 503418
rect 571500 503098 571532 503334
rect 571768 503098 571852 503334
rect 572088 503098 572120 503334
rect 571500 503066 572120 503098
rect -2006 483418 -1974 483654
rect -1738 483418 -1654 483654
rect -1418 483418 -1386 483654
rect -2006 483334 -1386 483418
rect -2006 483098 -1974 483334
rect -1738 483098 -1654 483334
rect -1418 483098 -1386 483334
rect -2006 443654 -1386 483098
rect 9084 483654 9704 483686
rect 9084 483418 9116 483654
rect 9352 483418 9436 483654
rect 9672 483418 9704 483654
rect 9084 483334 9704 483418
rect 9084 483098 9116 483334
rect 9352 483098 9436 483334
rect 9672 483098 9704 483334
rect 9084 483066 9704 483098
rect 56620 483654 57240 483686
rect 56620 483418 56652 483654
rect 56888 483418 56972 483654
rect 57208 483418 57240 483654
rect 56620 483334 57240 483418
rect 56620 483098 56652 483334
rect 56888 483098 56972 483334
rect 57208 483098 57240 483334
rect 56620 483066 57240 483098
rect 61280 483654 61640 483686
rect 61280 483418 61342 483654
rect 61578 483418 61640 483654
rect 61280 483334 61640 483418
rect 61280 483098 61342 483334
rect 61578 483098 61640 483334
rect 61280 483066 61640 483098
rect 158316 483654 158676 483686
rect 158316 483418 158378 483654
rect 158614 483418 158676 483654
rect 158316 483334 158676 483418
rect 158316 483098 158378 483334
rect 158614 483098 158676 483334
rect 158316 483066 158676 483098
rect 164620 483654 165240 483686
rect 164620 483418 164652 483654
rect 164888 483418 164972 483654
rect 165208 483418 165240 483654
rect 164620 483334 165240 483418
rect 164620 483098 164652 483334
rect 164888 483098 164972 483334
rect 165208 483098 165240 483334
rect 164620 483066 165240 483098
rect 186280 483654 186640 483686
rect 186280 483418 186342 483654
rect 186578 483418 186640 483654
rect 186280 483334 186640 483418
rect 186280 483098 186342 483334
rect 186578 483098 186640 483334
rect 186280 483066 186640 483098
rect 283316 483654 283676 483686
rect 283316 483418 283378 483654
rect 283614 483418 283676 483654
rect 283316 483334 283676 483418
rect 283316 483098 283378 483334
rect 283614 483098 283676 483334
rect 283316 483066 283676 483098
rect 308620 483654 309240 483686
rect 308620 483418 308652 483654
rect 308888 483418 308972 483654
rect 309208 483418 309240 483654
rect 308620 483334 309240 483418
rect 308620 483098 308652 483334
rect 308888 483098 308972 483334
rect 309208 483098 309240 483334
rect 308620 483066 309240 483098
rect 311280 483654 311640 483686
rect 311280 483418 311342 483654
rect 311578 483418 311640 483654
rect 311280 483334 311640 483418
rect 311280 483098 311342 483334
rect 311578 483098 311640 483334
rect 311280 483066 311640 483098
rect 408316 483654 408676 483686
rect 408316 483418 408378 483654
rect 408614 483418 408676 483654
rect 408316 483334 408676 483418
rect 408316 483098 408378 483334
rect 408614 483098 408676 483334
rect 408316 483066 408676 483098
rect 416620 483654 417240 483686
rect 416620 483418 416652 483654
rect 416888 483418 416972 483654
rect 417208 483418 417240 483654
rect 416620 483334 417240 483418
rect 416620 483098 416652 483334
rect 416888 483098 416972 483334
rect 417208 483098 417240 483334
rect 416620 483066 417240 483098
rect 437280 483654 437640 483686
rect 437280 483418 437342 483654
rect 437578 483418 437640 483654
rect 437280 483334 437640 483418
rect 437280 483098 437342 483334
rect 437578 483098 437640 483334
rect 437280 483066 437640 483098
rect 534316 483654 534676 483686
rect 534316 483418 534378 483654
rect 534614 483418 534676 483654
rect 534316 483334 534676 483418
rect 534316 483098 534378 483334
rect 534614 483098 534676 483334
rect 534316 483066 534676 483098
rect 560620 483654 561240 483686
rect 560620 483418 560652 483654
rect 560888 483418 560972 483654
rect 561208 483418 561240 483654
rect 560620 483334 561240 483418
rect 560620 483098 560652 483334
rect 560888 483098 560972 483334
rect 561208 483098 561240 483334
rect 560620 483066 561240 483098
rect 570260 483654 570880 483686
rect 570260 483418 570292 483654
rect 570528 483418 570612 483654
rect 570848 483418 570880 483654
rect 570260 483334 570880 483418
rect 570260 483098 570292 483334
rect 570528 483098 570612 483334
rect 570848 483098 570880 483334
rect 570260 483066 570880 483098
rect 585310 483654 585930 523098
rect 585310 483418 585342 483654
rect 585578 483418 585662 483654
rect 585898 483418 585930 483654
rect 585310 483334 585930 483418
rect 585310 483098 585342 483334
rect 585578 483098 585662 483334
rect 585898 483098 585930 483334
rect 7844 463654 8464 463686
rect 7844 463418 7876 463654
rect 8112 463418 8196 463654
rect 8432 463418 8464 463654
rect 7844 463334 8464 463418
rect 7844 463098 7876 463334
rect 8112 463098 8196 463334
rect 8432 463098 8464 463334
rect 7844 463066 8464 463098
rect 38000 463654 38620 463686
rect 38000 463418 38032 463654
rect 38268 463418 38352 463654
rect 38588 463418 38620 463654
rect 38000 463334 38620 463418
rect 38000 463098 38032 463334
rect 38268 463098 38352 463334
rect 38588 463098 38620 463334
rect 38000 463066 38620 463098
rect 60560 463654 60920 463686
rect 60560 463418 60622 463654
rect 60858 463418 60920 463654
rect 60560 463334 60920 463418
rect 60560 463098 60622 463334
rect 60858 463098 60920 463334
rect 60560 463066 60920 463098
rect 159036 463654 159396 463686
rect 159036 463418 159098 463654
rect 159334 463418 159396 463654
rect 159036 463334 159396 463418
rect 159036 463098 159098 463334
rect 159334 463098 159396 463334
rect 159036 463066 159396 463098
rect 182000 463654 182620 463686
rect 182000 463418 182032 463654
rect 182268 463418 182352 463654
rect 182588 463418 182620 463654
rect 182000 463334 182620 463418
rect 182000 463098 182032 463334
rect 182268 463098 182352 463334
rect 182588 463098 182620 463334
rect 182000 463066 182620 463098
rect 185560 463654 185920 463686
rect 185560 463418 185622 463654
rect 185858 463418 185920 463654
rect 185560 463334 185920 463418
rect 185560 463098 185622 463334
rect 185858 463098 185920 463334
rect 185560 463066 185920 463098
rect 284036 463654 284396 463686
rect 284036 463418 284098 463654
rect 284334 463418 284396 463654
rect 284036 463334 284396 463418
rect 284036 463098 284098 463334
rect 284334 463098 284396 463334
rect 284036 463066 284396 463098
rect 290000 463654 290620 463686
rect 290000 463418 290032 463654
rect 290268 463418 290352 463654
rect 290588 463418 290620 463654
rect 290000 463334 290620 463418
rect 290000 463098 290032 463334
rect 290268 463098 290352 463334
rect 290588 463098 290620 463334
rect 290000 463066 290620 463098
rect 310560 463654 310920 463686
rect 310560 463418 310622 463654
rect 310858 463418 310920 463654
rect 310560 463334 310920 463418
rect 310560 463098 310622 463334
rect 310858 463098 310920 463334
rect 310560 463066 310920 463098
rect 409036 463654 409396 463686
rect 409036 463418 409098 463654
rect 409334 463418 409396 463654
rect 409036 463334 409396 463418
rect 409036 463098 409098 463334
rect 409334 463098 409396 463334
rect 409036 463066 409396 463098
rect 434000 463654 434620 463686
rect 434000 463418 434032 463654
rect 434268 463418 434352 463654
rect 434588 463418 434620 463654
rect 434000 463334 434620 463418
rect 434000 463098 434032 463334
rect 434268 463098 434352 463334
rect 434588 463098 434620 463334
rect 434000 463066 434620 463098
rect 436560 463654 436920 463686
rect 436560 463418 436622 463654
rect 436858 463418 436920 463654
rect 436560 463334 436920 463418
rect 436560 463098 436622 463334
rect 436858 463098 436920 463334
rect 436560 463066 436920 463098
rect 535036 463654 535396 463686
rect 535036 463418 535098 463654
rect 535334 463418 535396 463654
rect 535036 463334 535396 463418
rect 535036 463098 535098 463334
rect 535334 463098 535396 463334
rect 535036 463066 535396 463098
rect 542000 463654 542620 463686
rect 542000 463418 542032 463654
rect 542268 463418 542352 463654
rect 542588 463418 542620 463654
rect 542000 463334 542620 463418
rect 542000 463098 542032 463334
rect 542268 463098 542352 463334
rect 542588 463098 542620 463334
rect 542000 463066 542620 463098
rect 571500 463654 572120 463686
rect 571500 463418 571532 463654
rect 571768 463418 571852 463654
rect 572088 463418 572120 463654
rect 571500 463334 572120 463418
rect 571500 463098 571532 463334
rect 571768 463098 571852 463334
rect 572088 463098 572120 463334
rect 571500 463066 572120 463098
rect -2006 443418 -1974 443654
rect -1738 443418 -1654 443654
rect -1418 443418 -1386 443654
rect -2006 443334 -1386 443418
rect -2006 443098 -1974 443334
rect -1738 443098 -1654 443334
rect -1418 443098 -1386 443334
rect -2006 403654 -1386 443098
rect 9084 443654 9704 443686
rect 9084 443418 9116 443654
rect 9352 443418 9436 443654
rect 9672 443418 9704 443654
rect 9084 443334 9704 443418
rect 9084 443098 9116 443334
rect 9352 443098 9436 443334
rect 9672 443098 9704 443334
rect 9084 443066 9704 443098
rect 56620 443654 57240 443686
rect 56620 443418 56652 443654
rect 56888 443418 56972 443654
rect 57208 443418 57240 443654
rect 56620 443334 57240 443418
rect 56620 443098 56652 443334
rect 56888 443098 56972 443334
rect 57208 443098 57240 443334
rect 56620 443066 57240 443098
rect 61280 443654 61640 443686
rect 61280 443418 61342 443654
rect 61578 443418 61640 443654
rect 61280 443334 61640 443418
rect 61280 443098 61342 443334
rect 61578 443098 61640 443334
rect 61280 443066 61640 443098
rect 158316 443654 158676 443686
rect 158316 443418 158378 443654
rect 158614 443418 158676 443654
rect 158316 443334 158676 443418
rect 158316 443098 158378 443334
rect 158614 443098 158676 443334
rect 158316 443066 158676 443098
rect 164620 443654 165240 443686
rect 164620 443418 164652 443654
rect 164888 443418 164972 443654
rect 165208 443418 165240 443654
rect 164620 443334 165240 443418
rect 164620 443098 164652 443334
rect 164888 443098 164972 443334
rect 165208 443098 165240 443334
rect 164620 443066 165240 443098
rect 186280 443654 186640 443686
rect 186280 443418 186342 443654
rect 186578 443418 186640 443654
rect 186280 443334 186640 443418
rect 186280 443098 186342 443334
rect 186578 443098 186640 443334
rect 186280 443066 186640 443098
rect 283316 443654 283676 443686
rect 283316 443418 283378 443654
rect 283614 443418 283676 443654
rect 283316 443334 283676 443418
rect 283316 443098 283378 443334
rect 283614 443098 283676 443334
rect 283316 443066 283676 443098
rect 308620 443654 309240 443686
rect 308620 443418 308652 443654
rect 308888 443418 308972 443654
rect 309208 443418 309240 443654
rect 308620 443334 309240 443418
rect 308620 443098 308652 443334
rect 308888 443098 308972 443334
rect 309208 443098 309240 443334
rect 308620 443066 309240 443098
rect 311280 443654 311640 443686
rect 311280 443418 311342 443654
rect 311578 443418 311640 443654
rect 311280 443334 311640 443418
rect 311280 443098 311342 443334
rect 311578 443098 311640 443334
rect 311280 443066 311640 443098
rect 408316 443654 408676 443686
rect 408316 443418 408378 443654
rect 408614 443418 408676 443654
rect 408316 443334 408676 443418
rect 408316 443098 408378 443334
rect 408614 443098 408676 443334
rect 408316 443066 408676 443098
rect 416620 443654 417240 443686
rect 416620 443418 416652 443654
rect 416888 443418 416972 443654
rect 417208 443418 417240 443654
rect 416620 443334 417240 443418
rect 416620 443098 416652 443334
rect 416888 443098 416972 443334
rect 417208 443098 417240 443334
rect 416620 443066 417240 443098
rect 437280 443654 437640 443686
rect 437280 443418 437342 443654
rect 437578 443418 437640 443654
rect 437280 443334 437640 443418
rect 437280 443098 437342 443334
rect 437578 443098 437640 443334
rect 437280 443066 437640 443098
rect 534316 443654 534676 443686
rect 534316 443418 534378 443654
rect 534614 443418 534676 443654
rect 534316 443334 534676 443418
rect 534316 443098 534378 443334
rect 534614 443098 534676 443334
rect 534316 443066 534676 443098
rect 560620 443654 561240 443686
rect 560620 443418 560652 443654
rect 560888 443418 560972 443654
rect 561208 443418 561240 443654
rect 560620 443334 561240 443418
rect 560620 443098 560652 443334
rect 560888 443098 560972 443334
rect 561208 443098 561240 443334
rect 560620 443066 561240 443098
rect 570260 443654 570880 443686
rect 570260 443418 570292 443654
rect 570528 443418 570612 443654
rect 570848 443418 570880 443654
rect 570260 443334 570880 443418
rect 570260 443098 570292 443334
rect 570528 443098 570612 443334
rect 570848 443098 570880 443334
rect 570260 443066 570880 443098
rect 585310 443654 585930 483098
rect 585310 443418 585342 443654
rect 585578 443418 585662 443654
rect 585898 443418 585930 443654
rect 585310 443334 585930 443418
rect 585310 443098 585342 443334
rect 585578 443098 585662 443334
rect 585898 443098 585930 443334
rect 7844 423654 8464 423686
rect 7844 423418 7876 423654
rect 8112 423418 8196 423654
rect 8432 423418 8464 423654
rect 7844 423334 8464 423418
rect 7844 423098 7876 423334
rect 8112 423098 8196 423334
rect 8432 423098 8464 423334
rect 7844 423066 8464 423098
rect 38000 423654 38620 423686
rect 38000 423418 38032 423654
rect 38268 423418 38352 423654
rect 38588 423418 38620 423654
rect 38000 423334 38620 423418
rect 38000 423098 38032 423334
rect 38268 423098 38352 423334
rect 38588 423098 38620 423334
rect 38000 423066 38620 423098
rect 74000 423654 74620 423686
rect 74000 423418 74032 423654
rect 74268 423418 74352 423654
rect 74588 423418 74620 423654
rect 74000 423334 74620 423418
rect 74000 423098 74032 423334
rect 74268 423098 74352 423334
rect 74588 423098 74620 423334
rect 74000 423066 74620 423098
rect 110000 423654 110620 423686
rect 110000 423418 110032 423654
rect 110268 423418 110352 423654
rect 110588 423418 110620 423654
rect 110000 423334 110620 423418
rect 110000 423098 110032 423334
rect 110268 423098 110352 423334
rect 110588 423098 110620 423334
rect 110000 423066 110620 423098
rect 146000 423654 146620 423686
rect 146000 423418 146032 423654
rect 146268 423418 146352 423654
rect 146588 423418 146620 423654
rect 146000 423334 146620 423418
rect 146000 423098 146032 423334
rect 146268 423098 146352 423334
rect 146588 423098 146620 423334
rect 146000 423066 146620 423098
rect 182000 423654 182620 423686
rect 182000 423418 182032 423654
rect 182268 423418 182352 423654
rect 182588 423418 182620 423654
rect 182000 423334 182620 423418
rect 182000 423098 182032 423334
rect 182268 423098 182352 423334
rect 182588 423098 182620 423334
rect 182000 423066 182620 423098
rect 218000 423654 218620 423686
rect 218000 423418 218032 423654
rect 218268 423418 218352 423654
rect 218588 423418 218620 423654
rect 218000 423334 218620 423418
rect 218000 423098 218032 423334
rect 218268 423098 218352 423334
rect 218588 423098 218620 423334
rect 218000 423066 218620 423098
rect 254000 423654 254620 423686
rect 254000 423418 254032 423654
rect 254268 423418 254352 423654
rect 254588 423418 254620 423654
rect 254000 423334 254620 423418
rect 254000 423098 254032 423334
rect 254268 423098 254352 423334
rect 254588 423098 254620 423334
rect 254000 423066 254620 423098
rect 290000 423654 290620 423686
rect 290000 423418 290032 423654
rect 290268 423418 290352 423654
rect 290588 423418 290620 423654
rect 290000 423334 290620 423418
rect 290000 423098 290032 423334
rect 290268 423098 290352 423334
rect 290588 423098 290620 423334
rect 290000 423066 290620 423098
rect 326000 423654 326620 423686
rect 326000 423418 326032 423654
rect 326268 423418 326352 423654
rect 326588 423418 326620 423654
rect 326000 423334 326620 423418
rect 326000 423098 326032 423334
rect 326268 423098 326352 423334
rect 326588 423098 326620 423334
rect 326000 423066 326620 423098
rect 362000 423654 362620 423686
rect 362000 423418 362032 423654
rect 362268 423418 362352 423654
rect 362588 423418 362620 423654
rect 362000 423334 362620 423418
rect 362000 423098 362032 423334
rect 362268 423098 362352 423334
rect 362588 423098 362620 423334
rect 362000 423066 362620 423098
rect 398000 423654 398620 423686
rect 398000 423418 398032 423654
rect 398268 423418 398352 423654
rect 398588 423418 398620 423654
rect 398000 423334 398620 423418
rect 398000 423098 398032 423334
rect 398268 423098 398352 423334
rect 398588 423098 398620 423334
rect 398000 423066 398620 423098
rect 434000 423654 434620 423686
rect 434000 423418 434032 423654
rect 434268 423418 434352 423654
rect 434588 423418 434620 423654
rect 434000 423334 434620 423418
rect 434000 423098 434032 423334
rect 434268 423098 434352 423334
rect 434588 423098 434620 423334
rect 434000 423066 434620 423098
rect 470000 423654 470620 423686
rect 470000 423418 470032 423654
rect 470268 423418 470352 423654
rect 470588 423418 470620 423654
rect 470000 423334 470620 423418
rect 470000 423098 470032 423334
rect 470268 423098 470352 423334
rect 470588 423098 470620 423334
rect 470000 423066 470620 423098
rect 506000 423654 506620 423686
rect 506000 423418 506032 423654
rect 506268 423418 506352 423654
rect 506588 423418 506620 423654
rect 506000 423334 506620 423418
rect 506000 423098 506032 423334
rect 506268 423098 506352 423334
rect 506588 423098 506620 423334
rect 506000 423066 506620 423098
rect 542000 423654 542620 423686
rect 542000 423418 542032 423654
rect 542268 423418 542352 423654
rect 542588 423418 542620 423654
rect 542000 423334 542620 423418
rect 542000 423098 542032 423334
rect 542268 423098 542352 423334
rect 542588 423098 542620 423334
rect 542000 423066 542620 423098
rect 571500 423654 572120 423686
rect 571500 423418 571532 423654
rect 571768 423418 571852 423654
rect 572088 423418 572120 423654
rect 571500 423334 572120 423418
rect 571500 423098 571532 423334
rect 571768 423098 571852 423334
rect 572088 423098 572120 423334
rect 571500 423066 572120 423098
rect -2006 403418 -1974 403654
rect -1738 403418 -1654 403654
rect -1418 403418 -1386 403654
rect -2006 403334 -1386 403418
rect -2006 403098 -1974 403334
rect -1738 403098 -1654 403334
rect -1418 403098 -1386 403334
rect -2006 363654 -1386 403098
rect 9084 403654 9704 403686
rect 9084 403418 9116 403654
rect 9352 403418 9436 403654
rect 9672 403418 9704 403654
rect 9084 403334 9704 403418
rect 9084 403098 9116 403334
rect 9352 403098 9436 403334
rect 9672 403098 9704 403334
rect 9084 403066 9704 403098
rect 56620 403654 57240 403686
rect 56620 403418 56652 403654
rect 56888 403418 56972 403654
rect 57208 403418 57240 403654
rect 56620 403334 57240 403418
rect 56620 403098 56652 403334
rect 56888 403098 56972 403334
rect 57208 403098 57240 403334
rect 56620 403066 57240 403098
rect 92620 403654 93240 403686
rect 92620 403418 92652 403654
rect 92888 403418 92972 403654
rect 93208 403418 93240 403654
rect 92620 403334 93240 403418
rect 92620 403098 92652 403334
rect 92888 403098 92972 403334
rect 93208 403098 93240 403334
rect 92620 403066 93240 403098
rect 128620 403654 129240 403686
rect 128620 403418 128652 403654
rect 128888 403418 128972 403654
rect 129208 403418 129240 403654
rect 128620 403334 129240 403418
rect 128620 403098 128652 403334
rect 128888 403098 128972 403334
rect 129208 403098 129240 403334
rect 128620 403066 129240 403098
rect 164620 403654 165240 403686
rect 164620 403418 164652 403654
rect 164888 403418 164972 403654
rect 165208 403418 165240 403654
rect 164620 403334 165240 403418
rect 164620 403098 164652 403334
rect 164888 403098 164972 403334
rect 165208 403098 165240 403334
rect 164620 403066 165240 403098
rect 200620 403654 201240 403686
rect 200620 403418 200652 403654
rect 200888 403418 200972 403654
rect 201208 403418 201240 403654
rect 200620 403334 201240 403418
rect 200620 403098 200652 403334
rect 200888 403098 200972 403334
rect 201208 403098 201240 403334
rect 200620 403066 201240 403098
rect 236620 403654 237240 403686
rect 236620 403418 236652 403654
rect 236888 403418 236972 403654
rect 237208 403418 237240 403654
rect 236620 403334 237240 403418
rect 236620 403098 236652 403334
rect 236888 403098 236972 403334
rect 237208 403098 237240 403334
rect 236620 403066 237240 403098
rect 272620 403654 273240 403686
rect 272620 403418 272652 403654
rect 272888 403418 272972 403654
rect 273208 403418 273240 403654
rect 272620 403334 273240 403418
rect 272620 403098 272652 403334
rect 272888 403098 272972 403334
rect 273208 403098 273240 403334
rect 272620 403066 273240 403098
rect 308620 403654 309240 403686
rect 308620 403418 308652 403654
rect 308888 403418 308972 403654
rect 309208 403418 309240 403654
rect 308620 403334 309240 403418
rect 308620 403098 308652 403334
rect 308888 403098 308972 403334
rect 309208 403098 309240 403334
rect 308620 403066 309240 403098
rect 344620 403654 345240 403686
rect 344620 403418 344652 403654
rect 344888 403418 344972 403654
rect 345208 403418 345240 403654
rect 344620 403334 345240 403418
rect 344620 403098 344652 403334
rect 344888 403098 344972 403334
rect 345208 403098 345240 403334
rect 344620 403066 345240 403098
rect 380620 403654 381240 403686
rect 380620 403418 380652 403654
rect 380888 403418 380972 403654
rect 381208 403418 381240 403654
rect 380620 403334 381240 403418
rect 380620 403098 380652 403334
rect 380888 403098 380972 403334
rect 381208 403098 381240 403334
rect 380620 403066 381240 403098
rect 416620 403654 417240 403686
rect 416620 403418 416652 403654
rect 416888 403418 416972 403654
rect 417208 403418 417240 403654
rect 416620 403334 417240 403418
rect 416620 403098 416652 403334
rect 416888 403098 416972 403334
rect 417208 403098 417240 403334
rect 416620 403066 417240 403098
rect 452620 403654 453240 403686
rect 452620 403418 452652 403654
rect 452888 403418 452972 403654
rect 453208 403418 453240 403654
rect 452620 403334 453240 403418
rect 452620 403098 452652 403334
rect 452888 403098 452972 403334
rect 453208 403098 453240 403334
rect 452620 403066 453240 403098
rect 488620 403654 489240 403686
rect 488620 403418 488652 403654
rect 488888 403418 488972 403654
rect 489208 403418 489240 403654
rect 488620 403334 489240 403418
rect 488620 403098 488652 403334
rect 488888 403098 488972 403334
rect 489208 403098 489240 403334
rect 488620 403066 489240 403098
rect 524620 403654 525240 403686
rect 524620 403418 524652 403654
rect 524888 403418 524972 403654
rect 525208 403418 525240 403654
rect 524620 403334 525240 403418
rect 524620 403098 524652 403334
rect 524888 403098 524972 403334
rect 525208 403098 525240 403334
rect 524620 403066 525240 403098
rect 560620 403654 561240 403686
rect 560620 403418 560652 403654
rect 560888 403418 560972 403654
rect 561208 403418 561240 403654
rect 560620 403334 561240 403418
rect 560620 403098 560652 403334
rect 560888 403098 560972 403334
rect 561208 403098 561240 403334
rect 560620 403066 561240 403098
rect 570260 403654 570880 403686
rect 570260 403418 570292 403654
rect 570528 403418 570612 403654
rect 570848 403418 570880 403654
rect 570260 403334 570880 403418
rect 570260 403098 570292 403334
rect 570528 403098 570612 403334
rect 570848 403098 570880 403334
rect 570260 403066 570880 403098
rect 585310 403654 585930 443098
rect 585310 403418 585342 403654
rect 585578 403418 585662 403654
rect 585898 403418 585930 403654
rect 585310 403334 585930 403418
rect 585310 403098 585342 403334
rect 585578 403098 585662 403334
rect 585898 403098 585930 403334
rect 7844 383654 8464 383686
rect 7844 383418 7876 383654
rect 8112 383418 8196 383654
rect 8432 383418 8464 383654
rect 7844 383334 8464 383418
rect 7844 383098 7876 383334
rect 8112 383098 8196 383334
rect 8432 383098 8464 383334
rect 7844 383066 8464 383098
rect 38000 383654 38620 383686
rect 38000 383418 38032 383654
rect 38268 383418 38352 383654
rect 38588 383418 38620 383654
rect 38000 383334 38620 383418
rect 38000 383098 38032 383334
rect 38268 383098 38352 383334
rect 38588 383098 38620 383334
rect 38000 383066 38620 383098
rect 74000 383654 74620 383686
rect 74000 383418 74032 383654
rect 74268 383418 74352 383654
rect 74588 383418 74620 383654
rect 74000 383334 74620 383418
rect 74000 383098 74032 383334
rect 74268 383098 74352 383334
rect 74588 383098 74620 383334
rect 74000 383066 74620 383098
rect 110000 383654 110620 383686
rect 110000 383418 110032 383654
rect 110268 383418 110352 383654
rect 110588 383418 110620 383654
rect 110000 383334 110620 383418
rect 110000 383098 110032 383334
rect 110268 383098 110352 383334
rect 110588 383098 110620 383334
rect 110000 383066 110620 383098
rect 146000 383654 146620 383686
rect 146000 383418 146032 383654
rect 146268 383418 146352 383654
rect 146588 383418 146620 383654
rect 146000 383334 146620 383418
rect 146000 383098 146032 383334
rect 146268 383098 146352 383334
rect 146588 383098 146620 383334
rect 146000 383066 146620 383098
rect 182000 383654 182620 383686
rect 182000 383418 182032 383654
rect 182268 383418 182352 383654
rect 182588 383418 182620 383654
rect 182000 383334 182620 383418
rect 182000 383098 182032 383334
rect 182268 383098 182352 383334
rect 182588 383098 182620 383334
rect 182000 383066 182620 383098
rect 218000 383654 218620 383686
rect 218000 383418 218032 383654
rect 218268 383418 218352 383654
rect 218588 383418 218620 383654
rect 218000 383334 218620 383418
rect 218000 383098 218032 383334
rect 218268 383098 218352 383334
rect 218588 383098 218620 383334
rect 218000 383066 218620 383098
rect 254000 383654 254620 383686
rect 254000 383418 254032 383654
rect 254268 383418 254352 383654
rect 254588 383418 254620 383654
rect 254000 383334 254620 383418
rect 254000 383098 254032 383334
rect 254268 383098 254352 383334
rect 254588 383098 254620 383334
rect 254000 383066 254620 383098
rect 290000 383654 290620 383686
rect 290000 383418 290032 383654
rect 290268 383418 290352 383654
rect 290588 383418 290620 383654
rect 290000 383334 290620 383418
rect 290000 383098 290032 383334
rect 290268 383098 290352 383334
rect 290588 383098 290620 383334
rect 290000 383066 290620 383098
rect 326000 383654 326620 383686
rect 326000 383418 326032 383654
rect 326268 383418 326352 383654
rect 326588 383418 326620 383654
rect 326000 383334 326620 383418
rect 326000 383098 326032 383334
rect 326268 383098 326352 383334
rect 326588 383098 326620 383334
rect 326000 383066 326620 383098
rect 362000 383654 362620 383686
rect 362000 383418 362032 383654
rect 362268 383418 362352 383654
rect 362588 383418 362620 383654
rect 362000 383334 362620 383418
rect 362000 383098 362032 383334
rect 362268 383098 362352 383334
rect 362588 383098 362620 383334
rect 362000 383066 362620 383098
rect 398000 383654 398620 383686
rect 398000 383418 398032 383654
rect 398268 383418 398352 383654
rect 398588 383418 398620 383654
rect 398000 383334 398620 383418
rect 398000 383098 398032 383334
rect 398268 383098 398352 383334
rect 398588 383098 398620 383334
rect 398000 383066 398620 383098
rect 434000 383654 434620 383686
rect 434000 383418 434032 383654
rect 434268 383418 434352 383654
rect 434588 383418 434620 383654
rect 434000 383334 434620 383418
rect 434000 383098 434032 383334
rect 434268 383098 434352 383334
rect 434588 383098 434620 383334
rect 434000 383066 434620 383098
rect 470000 383654 470620 383686
rect 470000 383418 470032 383654
rect 470268 383418 470352 383654
rect 470588 383418 470620 383654
rect 470000 383334 470620 383418
rect 470000 383098 470032 383334
rect 470268 383098 470352 383334
rect 470588 383098 470620 383334
rect 470000 383066 470620 383098
rect 506000 383654 506620 383686
rect 506000 383418 506032 383654
rect 506268 383418 506352 383654
rect 506588 383418 506620 383654
rect 506000 383334 506620 383418
rect 506000 383098 506032 383334
rect 506268 383098 506352 383334
rect 506588 383098 506620 383334
rect 506000 383066 506620 383098
rect 542000 383654 542620 383686
rect 542000 383418 542032 383654
rect 542268 383418 542352 383654
rect 542588 383418 542620 383654
rect 542000 383334 542620 383418
rect 542000 383098 542032 383334
rect 542268 383098 542352 383334
rect 542588 383098 542620 383334
rect 542000 383066 542620 383098
rect 571500 383654 572120 383686
rect 571500 383418 571532 383654
rect 571768 383418 571852 383654
rect 572088 383418 572120 383654
rect 571500 383334 572120 383418
rect 571500 383098 571532 383334
rect 571768 383098 571852 383334
rect 572088 383098 572120 383334
rect 571500 383066 572120 383098
rect -2006 363418 -1974 363654
rect -1738 363418 -1654 363654
rect -1418 363418 -1386 363654
rect -2006 363334 -1386 363418
rect -2006 363098 -1974 363334
rect -1738 363098 -1654 363334
rect -1418 363098 -1386 363334
rect -2006 323654 -1386 363098
rect 9084 363654 9704 363686
rect 9084 363418 9116 363654
rect 9352 363418 9436 363654
rect 9672 363418 9704 363654
rect 9084 363334 9704 363418
rect 9084 363098 9116 363334
rect 9352 363098 9436 363334
rect 9672 363098 9704 363334
rect 9084 363066 9704 363098
rect 56620 363654 57240 363686
rect 56620 363418 56652 363654
rect 56888 363418 56972 363654
rect 57208 363418 57240 363654
rect 56620 363334 57240 363418
rect 56620 363098 56652 363334
rect 56888 363098 56972 363334
rect 57208 363098 57240 363334
rect 56620 363066 57240 363098
rect 92620 363654 93240 363686
rect 92620 363418 92652 363654
rect 92888 363418 92972 363654
rect 93208 363418 93240 363654
rect 92620 363334 93240 363418
rect 92620 363098 92652 363334
rect 92888 363098 92972 363334
rect 93208 363098 93240 363334
rect 92620 363066 93240 363098
rect 128620 363654 129240 363686
rect 128620 363418 128652 363654
rect 128888 363418 128972 363654
rect 129208 363418 129240 363654
rect 128620 363334 129240 363418
rect 128620 363098 128652 363334
rect 128888 363098 128972 363334
rect 129208 363098 129240 363334
rect 128620 363066 129240 363098
rect 164620 363654 165240 363686
rect 164620 363418 164652 363654
rect 164888 363418 164972 363654
rect 165208 363418 165240 363654
rect 164620 363334 165240 363418
rect 164620 363098 164652 363334
rect 164888 363098 164972 363334
rect 165208 363098 165240 363334
rect 164620 363066 165240 363098
rect 200620 363654 201240 363686
rect 200620 363418 200652 363654
rect 200888 363418 200972 363654
rect 201208 363418 201240 363654
rect 200620 363334 201240 363418
rect 200620 363098 200652 363334
rect 200888 363098 200972 363334
rect 201208 363098 201240 363334
rect 200620 363066 201240 363098
rect 236620 363654 237240 363686
rect 236620 363418 236652 363654
rect 236888 363418 236972 363654
rect 237208 363418 237240 363654
rect 236620 363334 237240 363418
rect 236620 363098 236652 363334
rect 236888 363098 236972 363334
rect 237208 363098 237240 363334
rect 236620 363066 237240 363098
rect 272620 363654 273240 363686
rect 272620 363418 272652 363654
rect 272888 363418 272972 363654
rect 273208 363418 273240 363654
rect 272620 363334 273240 363418
rect 272620 363098 272652 363334
rect 272888 363098 272972 363334
rect 273208 363098 273240 363334
rect 272620 363066 273240 363098
rect 308620 363654 309240 363686
rect 308620 363418 308652 363654
rect 308888 363418 308972 363654
rect 309208 363418 309240 363654
rect 308620 363334 309240 363418
rect 308620 363098 308652 363334
rect 308888 363098 308972 363334
rect 309208 363098 309240 363334
rect 308620 363066 309240 363098
rect 344620 363654 345240 363686
rect 344620 363418 344652 363654
rect 344888 363418 344972 363654
rect 345208 363418 345240 363654
rect 344620 363334 345240 363418
rect 344620 363098 344652 363334
rect 344888 363098 344972 363334
rect 345208 363098 345240 363334
rect 344620 363066 345240 363098
rect 380620 363654 381240 363686
rect 380620 363418 380652 363654
rect 380888 363418 380972 363654
rect 381208 363418 381240 363654
rect 380620 363334 381240 363418
rect 380620 363098 380652 363334
rect 380888 363098 380972 363334
rect 381208 363098 381240 363334
rect 380620 363066 381240 363098
rect 416620 363654 417240 363686
rect 416620 363418 416652 363654
rect 416888 363418 416972 363654
rect 417208 363418 417240 363654
rect 416620 363334 417240 363418
rect 416620 363098 416652 363334
rect 416888 363098 416972 363334
rect 417208 363098 417240 363334
rect 416620 363066 417240 363098
rect 452620 363654 453240 363686
rect 452620 363418 452652 363654
rect 452888 363418 452972 363654
rect 453208 363418 453240 363654
rect 452620 363334 453240 363418
rect 452620 363098 452652 363334
rect 452888 363098 452972 363334
rect 453208 363098 453240 363334
rect 452620 363066 453240 363098
rect 488620 363654 489240 363686
rect 488620 363418 488652 363654
rect 488888 363418 488972 363654
rect 489208 363418 489240 363654
rect 488620 363334 489240 363418
rect 488620 363098 488652 363334
rect 488888 363098 488972 363334
rect 489208 363098 489240 363334
rect 488620 363066 489240 363098
rect 524620 363654 525240 363686
rect 524620 363418 524652 363654
rect 524888 363418 524972 363654
rect 525208 363418 525240 363654
rect 524620 363334 525240 363418
rect 524620 363098 524652 363334
rect 524888 363098 524972 363334
rect 525208 363098 525240 363334
rect 524620 363066 525240 363098
rect 560620 363654 561240 363686
rect 560620 363418 560652 363654
rect 560888 363418 560972 363654
rect 561208 363418 561240 363654
rect 560620 363334 561240 363418
rect 560620 363098 560652 363334
rect 560888 363098 560972 363334
rect 561208 363098 561240 363334
rect 560620 363066 561240 363098
rect 570260 363654 570880 363686
rect 570260 363418 570292 363654
rect 570528 363418 570612 363654
rect 570848 363418 570880 363654
rect 570260 363334 570880 363418
rect 570260 363098 570292 363334
rect 570528 363098 570612 363334
rect 570848 363098 570880 363334
rect 570260 363066 570880 363098
rect 585310 363654 585930 403098
rect 585310 363418 585342 363654
rect 585578 363418 585662 363654
rect 585898 363418 585930 363654
rect 585310 363334 585930 363418
rect 585310 363098 585342 363334
rect 585578 363098 585662 363334
rect 585898 363098 585930 363334
rect 7844 343654 8464 343686
rect 7844 343418 7876 343654
rect 8112 343418 8196 343654
rect 8432 343418 8464 343654
rect 7844 343334 8464 343418
rect 7844 343098 7876 343334
rect 8112 343098 8196 343334
rect 8432 343098 8464 343334
rect 7844 343066 8464 343098
rect 38000 343654 38620 343686
rect 38000 343418 38032 343654
rect 38268 343418 38352 343654
rect 38588 343418 38620 343654
rect 38000 343334 38620 343418
rect 38000 343098 38032 343334
rect 38268 343098 38352 343334
rect 38588 343098 38620 343334
rect 38000 343066 38620 343098
rect 74000 343654 74620 343686
rect 74000 343418 74032 343654
rect 74268 343418 74352 343654
rect 74588 343418 74620 343654
rect 74000 343334 74620 343418
rect 74000 343098 74032 343334
rect 74268 343098 74352 343334
rect 74588 343098 74620 343334
rect 74000 343066 74620 343098
rect 110000 343654 110620 343686
rect 110000 343418 110032 343654
rect 110268 343418 110352 343654
rect 110588 343418 110620 343654
rect 110000 343334 110620 343418
rect 110000 343098 110032 343334
rect 110268 343098 110352 343334
rect 110588 343098 110620 343334
rect 110000 343066 110620 343098
rect 146000 343654 146620 343686
rect 146000 343418 146032 343654
rect 146268 343418 146352 343654
rect 146588 343418 146620 343654
rect 146000 343334 146620 343418
rect 146000 343098 146032 343334
rect 146268 343098 146352 343334
rect 146588 343098 146620 343334
rect 146000 343066 146620 343098
rect 182000 343654 182620 343686
rect 182000 343418 182032 343654
rect 182268 343418 182352 343654
rect 182588 343418 182620 343654
rect 182000 343334 182620 343418
rect 182000 343098 182032 343334
rect 182268 343098 182352 343334
rect 182588 343098 182620 343334
rect 182000 343066 182620 343098
rect 218000 343654 218620 343686
rect 218000 343418 218032 343654
rect 218268 343418 218352 343654
rect 218588 343418 218620 343654
rect 218000 343334 218620 343418
rect 218000 343098 218032 343334
rect 218268 343098 218352 343334
rect 218588 343098 218620 343334
rect 218000 343066 218620 343098
rect 254000 343654 254620 343686
rect 254000 343418 254032 343654
rect 254268 343418 254352 343654
rect 254588 343418 254620 343654
rect 254000 343334 254620 343418
rect 254000 343098 254032 343334
rect 254268 343098 254352 343334
rect 254588 343098 254620 343334
rect 254000 343066 254620 343098
rect 290000 343654 290620 343686
rect 290000 343418 290032 343654
rect 290268 343418 290352 343654
rect 290588 343418 290620 343654
rect 290000 343334 290620 343418
rect 290000 343098 290032 343334
rect 290268 343098 290352 343334
rect 290588 343098 290620 343334
rect 290000 343066 290620 343098
rect 326000 343654 326620 343686
rect 326000 343418 326032 343654
rect 326268 343418 326352 343654
rect 326588 343418 326620 343654
rect 326000 343334 326620 343418
rect 326000 343098 326032 343334
rect 326268 343098 326352 343334
rect 326588 343098 326620 343334
rect 326000 343066 326620 343098
rect 362000 343654 362620 343686
rect 362000 343418 362032 343654
rect 362268 343418 362352 343654
rect 362588 343418 362620 343654
rect 362000 343334 362620 343418
rect 362000 343098 362032 343334
rect 362268 343098 362352 343334
rect 362588 343098 362620 343334
rect 362000 343066 362620 343098
rect 398000 343654 398620 343686
rect 398000 343418 398032 343654
rect 398268 343418 398352 343654
rect 398588 343418 398620 343654
rect 398000 343334 398620 343418
rect 398000 343098 398032 343334
rect 398268 343098 398352 343334
rect 398588 343098 398620 343334
rect 398000 343066 398620 343098
rect 434000 343654 434620 343686
rect 434000 343418 434032 343654
rect 434268 343418 434352 343654
rect 434588 343418 434620 343654
rect 434000 343334 434620 343418
rect 434000 343098 434032 343334
rect 434268 343098 434352 343334
rect 434588 343098 434620 343334
rect 434000 343066 434620 343098
rect 470000 343654 470620 343686
rect 470000 343418 470032 343654
rect 470268 343418 470352 343654
rect 470588 343418 470620 343654
rect 470000 343334 470620 343418
rect 470000 343098 470032 343334
rect 470268 343098 470352 343334
rect 470588 343098 470620 343334
rect 470000 343066 470620 343098
rect 506000 343654 506620 343686
rect 506000 343418 506032 343654
rect 506268 343418 506352 343654
rect 506588 343418 506620 343654
rect 506000 343334 506620 343418
rect 506000 343098 506032 343334
rect 506268 343098 506352 343334
rect 506588 343098 506620 343334
rect 506000 343066 506620 343098
rect 542000 343654 542620 343686
rect 542000 343418 542032 343654
rect 542268 343418 542352 343654
rect 542588 343418 542620 343654
rect 542000 343334 542620 343418
rect 542000 343098 542032 343334
rect 542268 343098 542352 343334
rect 542588 343098 542620 343334
rect 542000 343066 542620 343098
rect 571500 343654 572120 343686
rect 571500 343418 571532 343654
rect 571768 343418 571852 343654
rect 572088 343418 572120 343654
rect 571500 343334 572120 343418
rect 571500 343098 571532 343334
rect 571768 343098 571852 343334
rect 572088 343098 572120 343334
rect 571500 343066 572120 343098
rect -2006 323418 -1974 323654
rect -1738 323418 -1654 323654
rect -1418 323418 -1386 323654
rect -2006 323334 -1386 323418
rect -2006 323098 -1974 323334
rect -1738 323098 -1654 323334
rect -1418 323098 -1386 323334
rect -2006 283654 -1386 323098
rect 9084 323654 9704 323686
rect 9084 323418 9116 323654
rect 9352 323418 9436 323654
rect 9672 323418 9704 323654
rect 9084 323334 9704 323418
rect 9084 323098 9116 323334
rect 9352 323098 9436 323334
rect 9672 323098 9704 323334
rect 9084 323066 9704 323098
rect 56620 323654 57240 323686
rect 56620 323418 56652 323654
rect 56888 323418 56972 323654
rect 57208 323418 57240 323654
rect 56620 323334 57240 323418
rect 56620 323098 56652 323334
rect 56888 323098 56972 323334
rect 57208 323098 57240 323334
rect 56620 323066 57240 323098
rect 92620 323654 93240 323686
rect 92620 323418 92652 323654
rect 92888 323418 92972 323654
rect 93208 323418 93240 323654
rect 92620 323334 93240 323418
rect 92620 323098 92652 323334
rect 92888 323098 92972 323334
rect 93208 323098 93240 323334
rect 92620 323066 93240 323098
rect 128620 323654 129240 323686
rect 128620 323418 128652 323654
rect 128888 323418 128972 323654
rect 129208 323418 129240 323654
rect 128620 323334 129240 323418
rect 128620 323098 128652 323334
rect 128888 323098 128972 323334
rect 129208 323098 129240 323334
rect 128620 323066 129240 323098
rect 164620 323654 165240 323686
rect 164620 323418 164652 323654
rect 164888 323418 164972 323654
rect 165208 323418 165240 323654
rect 164620 323334 165240 323418
rect 164620 323098 164652 323334
rect 164888 323098 164972 323334
rect 165208 323098 165240 323334
rect 164620 323066 165240 323098
rect 200620 323654 201240 323686
rect 200620 323418 200652 323654
rect 200888 323418 200972 323654
rect 201208 323418 201240 323654
rect 200620 323334 201240 323418
rect 200620 323098 200652 323334
rect 200888 323098 200972 323334
rect 201208 323098 201240 323334
rect 200620 323066 201240 323098
rect 236620 323654 237240 323686
rect 236620 323418 236652 323654
rect 236888 323418 236972 323654
rect 237208 323418 237240 323654
rect 236620 323334 237240 323418
rect 236620 323098 236652 323334
rect 236888 323098 236972 323334
rect 237208 323098 237240 323334
rect 236620 323066 237240 323098
rect 272620 323654 273240 323686
rect 272620 323418 272652 323654
rect 272888 323418 272972 323654
rect 273208 323418 273240 323654
rect 272620 323334 273240 323418
rect 272620 323098 272652 323334
rect 272888 323098 272972 323334
rect 273208 323098 273240 323334
rect 272620 323066 273240 323098
rect 308620 323654 309240 323686
rect 308620 323418 308652 323654
rect 308888 323418 308972 323654
rect 309208 323418 309240 323654
rect 308620 323334 309240 323418
rect 308620 323098 308652 323334
rect 308888 323098 308972 323334
rect 309208 323098 309240 323334
rect 308620 323066 309240 323098
rect 344620 323654 345240 323686
rect 344620 323418 344652 323654
rect 344888 323418 344972 323654
rect 345208 323418 345240 323654
rect 344620 323334 345240 323418
rect 344620 323098 344652 323334
rect 344888 323098 344972 323334
rect 345208 323098 345240 323334
rect 344620 323066 345240 323098
rect 380620 323654 381240 323686
rect 380620 323418 380652 323654
rect 380888 323418 380972 323654
rect 381208 323418 381240 323654
rect 380620 323334 381240 323418
rect 380620 323098 380652 323334
rect 380888 323098 380972 323334
rect 381208 323098 381240 323334
rect 380620 323066 381240 323098
rect 416620 323654 417240 323686
rect 416620 323418 416652 323654
rect 416888 323418 416972 323654
rect 417208 323418 417240 323654
rect 416620 323334 417240 323418
rect 416620 323098 416652 323334
rect 416888 323098 416972 323334
rect 417208 323098 417240 323334
rect 416620 323066 417240 323098
rect 452620 323654 453240 323686
rect 452620 323418 452652 323654
rect 452888 323418 452972 323654
rect 453208 323418 453240 323654
rect 452620 323334 453240 323418
rect 452620 323098 452652 323334
rect 452888 323098 452972 323334
rect 453208 323098 453240 323334
rect 452620 323066 453240 323098
rect 488620 323654 489240 323686
rect 488620 323418 488652 323654
rect 488888 323418 488972 323654
rect 489208 323418 489240 323654
rect 488620 323334 489240 323418
rect 488620 323098 488652 323334
rect 488888 323098 488972 323334
rect 489208 323098 489240 323334
rect 488620 323066 489240 323098
rect 524620 323654 525240 323686
rect 524620 323418 524652 323654
rect 524888 323418 524972 323654
rect 525208 323418 525240 323654
rect 524620 323334 525240 323418
rect 524620 323098 524652 323334
rect 524888 323098 524972 323334
rect 525208 323098 525240 323334
rect 524620 323066 525240 323098
rect 560620 323654 561240 323686
rect 560620 323418 560652 323654
rect 560888 323418 560972 323654
rect 561208 323418 561240 323654
rect 560620 323334 561240 323418
rect 560620 323098 560652 323334
rect 560888 323098 560972 323334
rect 561208 323098 561240 323334
rect 560620 323066 561240 323098
rect 570260 323654 570880 323686
rect 570260 323418 570292 323654
rect 570528 323418 570612 323654
rect 570848 323418 570880 323654
rect 570260 323334 570880 323418
rect 570260 323098 570292 323334
rect 570528 323098 570612 323334
rect 570848 323098 570880 323334
rect 570260 323066 570880 323098
rect 585310 323654 585930 363098
rect 585310 323418 585342 323654
rect 585578 323418 585662 323654
rect 585898 323418 585930 323654
rect 585310 323334 585930 323418
rect 585310 323098 585342 323334
rect 585578 323098 585662 323334
rect 585898 323098 585930 323334
rect 7844 303654 8464 303686
rect 7844 303418 7876 303654
rect 8112 303418 8196 303654
rect 8432 303418 8464 303654
rect 7844 303334 8464 303418
rect 7844 303098 7876 303334
rect 8112 303098 8196 303334
rect 8432 303098 8464 303334
rect 7844 303066 8464 303098
rect 38000 303654 38620 303686
rect 38000 303418 38032 303654
rect 38268 303418 38352 303654
rect 38588 303418 38620 303654
rect 38000 303334 38620 303418
rect 38000 303098 38032 303334
rect 38268 303098 38352 303334
rect 38588 303098 38620 303334
rect 38000 303066 38620 303098
rect 74000 303654 74620 303686
rect 74000 303418 74032 303654
rect 74268 303418 74352 303654
rect 74588 303418 74620 303654
rect 74000 303334 74620 303418
rect 74000 303098 74032 303334
rect 74268 303098 74352 303334
rect 74588 303098 74620 303334
rect 74000 303066 74620 303098
rect 110000 303654 110620 303686
rect 110000 303418 110032 303654
rect 110268 303418 110352 303654
rect 110588 303418 110620 303654
rect 110000 303334 110620 303418
rect 110000 303098 110032 303334
rect 110268 303098 110352 303334
rect 110588 303098 110620 303334
rect 110000 303066 110620 303098
rect 146000 303654 146620 303686
rect 146000 303418 146032 303654
rect 146268 303418 146352 303654
rect 146588 303418 146620 303654
rect 146000 303334 146620 303418
rect 146000 303098 146032 303334
rect 146268 303098 146352 303334
rect 146588 303098 146620 303334
rect 146000 303066 146620 303098
rect 182000 303654 182620 303686
rect 182000 303418 182032 303654
rect 182268 303418 182352 303654
rect 182588 303418 182620 303654
rect 182000 303334 182620 303418
rect 182000 303098 182032 303334
rect 182268 303098 182352 303334
rect 182588 303098 182620 303334
rect 182000 303066 182620 303098
rect 218000 303654 218620 303686
rect 218000 303418 218032 303654
rect 218268 303418 218352 303654
rect 218588 303418 218620 303654
rect 218000 303334 218620 303418
rect 218000 303098 218032 303334
rect 218268 303098 218352 303334
rect 218588 303098 218620 303334
rect 218000 303066 218620 303098
rect 254000 303654 254620 303686
rect 254000 303418 254032 303654
rect 254268 303418 254352 303654
rect 254588 303418 254620 303654
rect 254000 303334 254620 303418
rect 254000 303098 254032 303334
rect 254268 303098 254352 303334
rect 254588 303098 254620 303334
rect 254000 303066 254620 303098
rect 290000 303654 290620 303686
rect 290000 303418 290032 303654
rect 290268 303418 290352 303654
rect 290588 303418 290620 303654
rect 290000 303334 290620 303418
rect 290000 303098 290032 303334
rect 290268 303098 290352 303334
rect 290588 303098 290620 303334
rect 290000 303066 290620 303098
rect 326000 303654 326620 303686
rect 326000 303418 326032 303654
rect 326268 303418 326352 303654
rect 326588 303418 326620 303654
rect 326000 303334 326620 303418
rect 326000 303098 326032 303334
rect 326268 303098 326352 303334
rect 326588 303098 326620 303334
rect 326000 303066 326620 303098
rect 362000 303654 362620 303686
rect 362000 303418 362032 303654
rect 362268 303418 362352 303654
rect 362588 303418 362620 303654
rect 362000 303334 362620 303418
rect 362000 303098 362032 303334
rect 362268 303098 362352 303334
rect 362588 303098 362620 303334
rect 362000 303066 362620 303098
rect 398000 303654 398620 303686
rect 398000 303418 398032 303654
rect 398268 303418 398352 303654
rect 398588 303418 398620 303654
rect 398000 303334 398620 303418
rect 398000 303098 398032 303334
rect 398268 303098 398352 303334
rect 398588 303098 398620 303334
rect 398000 303066 398620 303098
rect 434000 303654 434620 303686
rect 434000 303418 434032 303654
rect 434268 303418 434352 303654
rect 434588 303418 434620 303654
rect 434000 303334 434620 303418
rect 434000 303098 434032 303334
rect 434268 303098 434352 303334
rect 434588 303098 434620 303334
rect 434000 303066 434620 303098
rect 470000 303654 470620 303686
rect 470000 303418 470032 303654
rect 470268 303418 470352 303654
rect 470588 303418 470620 303654
rect 470000 303334 470620 303418
rect 470000 303098 470032 303334
rect 470268 303098 470352 303334
rect 470588 303098 470620 303334
rect 470000 303066 470620 303098
rect 506000 303654 506620 303686
rect 506000 303418 506032 303654
rect 506268 303418 506352 303654
rect 506588 303418 506620 303654
rect 506000 303334 506620 303418
rect 506000 303098 506032 303334
rect 506268 303098 506352 303334
rect 506588 303098 506620 303334
rect 506000 303066 506620 303098
rect 542000 303654 542620 303686
rect 542000 303418 542032 303654
rect 542268 303418 542352 303654
rect 542588 303418 542620 303654
rect 542000 303334 542620 303418
rect 542000 303098 542032 303334
rect 542268 303098 542352 303334
rect 542588 303098 542620 303334
rect 542000 303066 542620 303098
rect 571500 303654 572120 303686
rect 571500 303418 571532 303654
rect 571768 303418 571852 303654
rect 572088 303418 572120 303654
rect 571500 303334 572120 303418
rect 571500 303098 571532 303334
rect 571768 303098 571852 303334
rect 572088 303098 572120 303334
rect 571500 303066 572120 303098
rect -2006 283418 -1974 283654
rect -1738 283418 -1654 283654
rect -1418 283418 -1386 283654
rect -2006 283334 -1386 283418
rect -2006 283098 -1974 283334
rect -1738 283098 -1654 283334
rect -1418 283098 -1386 283334
rect -2006 243654 -1386 283098
rect 9084 283654 9704 283686
rect 9084 283418 9116 283654
rect 9352 283418 9436 283654
rect 9672 283418 9704 283654
rect 9084 283334 9704 283418
rect 9084 283098 9116 283334
rect 9352 283098 9436 283334
rect 9672 283098 9704 283334
rect 9084 283066 9704 283098
rect 56620 283654 57240 283686
rect 56620 283418 56652 283654
rect 56888 283418 56972 283654
rect 57208 283418 57240 283654
rect 56620 283334 57240 283418
rect 56620 283098 56652 283334
rect 56888 283098 56972 283334
rect 57208 283098 57240 283334
rect 56620 283066 57240 283098
rect 92620 283654 93240 283686
rect 92620 283418 92652 283654
rect 92888 283418 92972 283654
rect 93208 283418 93240 283654
rect 92620 283334 93240 283418
rect 92620 283098 92652 283334
rect 92888 283098 92972 283334
rect 93208 283098 93240 283334
rect 92620 283066 93240 283098
rect 128620 283654 129240 283686
rect 128620 283418 128652 283654
rect 128888 283418 128972 283654
rect 129208 283418 129240 283654
rect 128620 283334 129240 283418
rect 128620 283098 128652 283334
rect 128888 283098 128972 283334
rect 129208 283098 129240 283334
rect 128620 283066 129240 283098
rect 164620 283654 165240 283686
rect 164620 283418 164652 283654
rect 164888 283418 164972 283654
rect 165208 283418 165240 283654
rect 164620 283334 165240 283418
rect 164620 283098 164652 283334
rect 164888 283098 164972 283334
rect 165208 283098 165240 283334
rect 164620 283066 165240 283098
rect 200620 283654 201240 283686
rect 200620 283418 200652 283654
rect 200888 283418 200972 283654
rect 201208 283418 201240 283654
rect 200620 283334 201240 283418
rect 200620 283098 200652 283334
rect 200888 283098 200972 283334
rect 201208 283098 201240 283334
rect 200620 283066 201240 283098
rect 236620 283654 237240 283686
rect 236620 283418 236652 283654
rect 236888 283418 236972 283654
rect 237208 283418 237240 283654
rect 236620 283334 237240 283418
rect 236620 283098 236652 283334
rect 236888 283098 236972 283334
rect 237208 283098 237240 283334
rect 236620 283066 237240 283098
rect 272620 283654 273240 283686
rect 272620 283418 272652 283654
rect 272888 283418 272972 283654
rect 273208 283418 273240 283654
rect 272620 283334 273240 283418
rect 272620 283098 272652 283334
rect 272888 283098 272972 283334
rect 273208 283098 273240 283334
rect 272620 283066 273240 283098
rect 308620 283654 309240 283686
rect 308620 283418 308652 283654
rect 308888 283418 308972 283654
rect 309208 283418 309240 283654
rect 308620 283334 309240 283418
rect 308620 283098 308652 283334
rect 308888 283098 308972 283334
rect 309208 283098 309240 283334
rect 308620 283066 309240 283098
rect 344620 283654 345240 283686
rect 344620 283418 344652 283654
rect 344888 283418 344972 283654
rect 345208 283418 345240 283654
rect 344620 283334 345240 283418
rect 344620 283098 344652 283334
rect 344888 283098 344972 283334
rect 345208 283098 345240 283334
rect 344620 283066 345240 283098
rect 380620 283654 381240 283686
rect 380620 283418 380652 283654
rect 380888 283418 380972 283654
rect 381208 283418 381240 283654
rect 380620 283334 381240 283418
rect 380620 283098 380652 283334
rect 380888 283098 380972 283334
rect 381208 283098 381240 283334
rect 380620 283066 381240 283098
rect 416620 283654 417240 283686
rect 416620 283418 416652 283654
rect 416888 283418 416972 283654
rect 417208 283418 417240 283654
rect 416620 283334 417240 283418
rect 416620 283098 416652 283334
rect 416888 283098 416972 283334
rect 417208 283098 417240 283334
rect 416620 283066 417240 283098
rect 452620 283654 453240 283686
rect 452620 283418 452652 283654
rect 452888 283418 452972 283654
rect 453208 283418 453240 283654
rect 452620 283334 453240 283418
rect 452620 283098 452652 283334
rect 452888 283098 452972 283334
rect 453208 283098 453240 283334
rect 452620 283066 453240 283098
rect 488620 283654 489240 283686
rect 488620 283418 488652 283654
rect 488888 283418 488972 283654
rect 489208 283418 489240 283654
rect 488620 283334 489240 283418
rect 488620 283098 488652 283334
rect 488888 283098 488972 283334
rect 489208 283098 489240 283334
rect 488620 283066 489240 283098
rect 524620 283654 525240 283686
rect 524620 283418 524652 283654
rect 524888 283418 524972 283654
rect 525208 283418 525240 283654
rect 524620 283334 525240 283418
rect 524620 283098 524652 283334
rect 524888 283098 524972 283334
rect 525208 283098 525240 283334
rect 524620 283066 525240 283098
rect 560620 283654 561240 283686
rect 560620 283418 560652 283654
rect 560888 283418 560972 283654
rect 561208 283418 561240 283654
rect 560620 283334 561240 283418
rect 560620 283098 560652 283334
rect 560888 283098 560972 283334
rect 561208 283098 561240 283334
rect 560620 283066 561240 283098
rect 570260 283654 570880 283686
rect 570260 283418 570292 283654
rect 570528 283418 570612 283654
rect 570848 283418 570880 283654
rect 570260 283334 570880 283418
rect 570260 283098 570292 283334
rect 570528 283098 570612 283334
rect 570848 283098 570880 283334
rect 570260 283066 570880 283098
rect 585310 283654 585930 323098
rect 585310 283418 585342 283654
rect 585578 283418 585662 283654
rect 585898 283418 585930 283654
rect 585310 283334 585930 283418
rect 585310 283098 585342 283334
rect 585578 283098 585662 283334
rect 585898 283098 585930 283334
rect 7844 263654 8464 263686
rect 7844 263418 7876 263654
rect 8112 263418 8196 263654
rect 8432 263418 8464 263654
rect 7844 263334 8464 263418
rect 7844 263098 7876 263334
rect 8112 263098 8196 263334
rect 8432 263098 8464 263334
rect 7844 263066 8464 263098
rect 38000 263654 38620 263686
rect 38000 263418 38032 263654
rect 38268 263418 38352 263654
rect 38588 263418 38620 263654
rect 38000 263334 38620 263418
rect 38000 263098 38032 263334
rect 38268 263098 38352 263334
rect 38588 263098 38620 263334
rect 38000 263066 38620 263098
rect 74000 263654 74620 263686
rect 74000 263418 74032 263654
rect 74268 263418 74352 263654
rect 74588 263418 74620 263654
rect 74000 263334 74620 263418
rect 74000 263098 74032 263334
rect 74268 263098 74352 263334
rect 74588 263098 74620 263334
rect 74000 263066 74620 263098
rect 110000 263654 110620 263686
rect 110000 263418 110032 263654
rect 110268 263418 110352 263654
rect 110588 263418 110620 263654
rect 110000 263334 110620 263418
rect 110000 263098 110032 263334
rect 110268 263098 110352 263334
rect 110588 263098 110620 263334
rect 110000 263066 110620 263098
rect 146000 263654 146620 263686
rect 146000 263418 146032 263654
rect 146268 263418 146352 263654
rect 146588 263418 146620 263654
rect 146000 263334 146620 263418
rect 146000 263098 146032 263334
rect 146268 263098 146352 263334
rect 146588 263098 146620 263334
rect 146000 263066 146620 263098
rect 182000 263654 182620 263686
rect 182000 263418 182032 263654
rect 182268 263418 182352 263654
rect 182588 263418 182620 263654
rect 182000 263334 182620 263418
rect 182000 263098 182032 263334
rect 182268 263098 182352 263334
rect 182588 263098 182620 263334
rect 182000 263066 182620 263098
rect 218000 263654 218620 263686
rect 218000 263418 218032 263654
rect 218268 263418 218352 263654
rect 218588 263418 218620 263654
rect 218000 263334 218620 263418
rect 218000 263098 218032 263334
rect 218268 263098 218352 263334
rect 218588 263098 218620 263334
rect 218000 263066 218620 263098
rect 254000 263654 254620 263686
rect 254000 263418 254032 263654
rect 254268 263418 254352 263654
rect 254588 263418 254620 263654
rect 254000 263334 254620 263418
rect 254000 263098 254032 263334
rect 254268 263098 254352 263334
rect 254588 263098 254620 263334
rect 254000 263066 254620 263098
rect 290000 263654 290620 263686
rect 290000 263418 290032 263654
rect 290268 263418 290352 263654
rect 290588 263418 290620 263654
rect 290000 263334 290620 263418
rect 290000 263098 290032 263334
rect 290268 263098 290352 263334
rect 290588 263098 290620 263334
rect 290000 263066 290620 263098
rect 326000 263654 326620 263686
rect 326000 263418 326032 263654
rect 326268 263418 326352 263654
rect 326588 263418 326620 263654
rect 326000 263334 326620 263418
rect 326000 263098 326032 263334
rect 326268 263098 326352 263334
rect 326588 263098 326620 263334
rect 326000 263066 326620 263098
rect 362000 263654 362620 263686
rect 362000 263418 362032 263654
rect 362268 263418 362352 263654
rect 362588 263418 362620 263654
rect 362000 263334 362620 263418
rect 362000 263098 362032 263334
rect 362268 263098 362352 263334
rect 362588 263098 362620 263334
rect 362000 263066 362620 263098
rect 398000 263654 398620 263686
rect 398000 263418 398032 263654
rect 398268 263418 398352 263654
rect 398588 263418 398620 263654
rect 398000 263334 398620 263418
rect 398000 263098 398032 263334
rect 398268 263098 398352 263334
rect 398588 263098 398620 263334
rect 398000 263066 398620 263098
rect 434000 263654 434620 263686
rect 434000 263418 434032 263654
rect 434268 263418 434352 263654
rect 434588 263418 434620 263654
rect 434000 263334 434620 263418
rect 434000 263098 434032 263334
rect 434268 263098 434352 263334
rect 434588 263098 434620 263334
rect 434000 263066 434620 263098
rect 470000 263654 470620 263686
rect 470000 263418 470032 263654
rect 470268 263418 470352 263654
rect 470588 263418 470620 263654
rect 470000 263334 470620 263418
rect 470000 263098 470032 263334
rect 470268 263098 470352 263334
rect 470588 263098 470620 263334
rect 470000 263066 470620 263098
rect 506000 263654 506620 263686
rect 506000 263418 506032 263654
rect 506268 263418 506352 263654
rect 506588 263418 506620 263654
rect 506000 263334 506620 263418
rect 506000 263098 506032 263334
rect 506268 263098 506352 263334
rect 506588 263098 506620 263334
rect 506000 263066 506620 263098
rect 542000 263654 542620 263686
rect 542000 263418 542032 263654
rect 542268 263418 542352 263654
rect 542588 263418 542620 263654
rect 542000 263334 542620 263418
rect 542000 263098 542032 263334
rect 542268 263098 542352 263334
rect 542588 263098 542620 263334
rect 542000 263066 542620 263098
rect 571500 263654 572120 263686
rect 571500 263418 571532 263654
rect 571768 263418 571852 263654
rect 572088 263418 572120 263654
rect 571500 263334 572120 263418
rect 571500 263098 571532 263334
rect 571768 263098 571852 263334
rect 572088 263098 572120 263334
rect 571500 263066 572120 263098
rect -2006 243418 -1974 243654
rect -1738 243418 -1654 243654
rect -1418 243418 -1386 243654
rect -2006 243334 -1386 243418
rect -2006 243098 -1974 243334
rect -1738 243098 -1654 243334
rect -1418 243098 -1386 243334
rect -2006 203654 -1386 243098
rect 9084 243654 9704 243686
rect 9084 243418 9116 243654
rect 9352 243418 9436 243654
rect 9672 243418 9704 243654
rect 9084 243334 9704 243418
rect 9084 243098 9116 243334
rect 9352 243098 9436 243334
rect 9672 243098 9704 243334
rect 9084 243066 9704 243098
rect 56620 243654 57240 243686
rect 56620 243418 56652 243654
rect 56888 243418 56972 243654
rect 57208 243418 57240 243654
rect 56620 243334 57240 243418
rect 56620 243098 56652 243334
rect 56888 243098 56972 243334
rect 57208 243098 57240 243334
rect 56620 243066 57240 243098
rect 92620 243654 93240 243686
rect 92620 243418 92652 243654
rect 92888 243418 92972 243654
rect 93208 243418 93240 243654
rect 92620 243334 93240 243418
rect 92620 243098 92652 243334
rect 92888 243098 92972 243334
rect 93208 243098 93240 243334
rect 92620 243066 93240 243098
rect 128620 243654 129240 243686
rect 128620 243418 128652 243654
rect 128888 243418 128972 243654
rect 129208 243418 129240 243654
rect 128620 243334 129240 243418
rect 128620 243098 128652 243334
rect 128888 243098 128972 243334
rect 129208 243098 129240 243334
rect 128620 243066 129240 243098
rect 164620 243654 165240 243686
rect 164620 243418 164652 243654
rect 164888 243418 164972 243654
rect 165208 243418 165240 243654
rect 164620 243334 165240 243418
rect 164620 243098 164652 243334
rect 164888 243098 164972 243334
rect 165208 243098 165240 243334
rect 164620 243066 165240 243098
rect 200620 243654 201240 243686
rect 200620 243418 200652 243654
rect 200888 243418 200972 243654
rect 201208 243418 201240 243654
rect 200620 243334 201240 243418
rect 200620 243098 200652 243334
rect 200888 243098 200972 243334
rect 201208 243098 201240 243334
rect 200620 243066 201240 243098
rect 236620 243654 237240 243686
rect 236620 243418 236652 243654
rect 236888 243418 236972 243654
rect 237208 243418 237240 243654
rect 236620 243334 237240 243418
rect 236620 243098 236652 243334
rect 236888 243098 236972 243334
rect 237208 243098 237240 243334
rect 236620 243066 237240 243098
rect 272620 243654 273240 243686
rect 272620 243418 272652 243654
rect 272888 243418 272972 243654
rect 273208 243418 273240 243654
rect 272620 243334 273240 243418
rect 272620 243098 272652 243334
rect 272888 243098 272972 243334
rect 273208 243098 273240 243334
rect 272620 243066 273240 243098
rect 308620 243654 309240 243686
rect 308620 243418 308652 243654
rect 308888 243418 308972 243654
rect 309208 243418 309240 243654
rect 308620 243334 309240 243418
rect 308620 243098 308652 243334
rect 308888 243098 308972 243334
rect 309208 243098 309240 243334
rect 308620 243066 309240 243098
rect 344620 243654 345240 243686
rect 344620 243418 344652 243654
rect 344888 243418 344972 243654
rect 345208 243418 345240 243654
rect 344620 243334 345240 243418
rect 344620 243098 344652 243334
rect 344888 243098 344972 243334
rect 345208 243098 345240 243334
rect 344620 243066 345240 243098
rect 380620 243654 381240 243686
rect 380620 243418 380652 243654
rect 380888 243418 380972 243654
rect 381208 243418 381240 243654
rect 380620 243334 381240 243418
rect 380620 243098 380652 243334
rect 380888 243098 380972 243334
rect 381208 243098 381240 243334
rect 380620 243066 381240 243098
rect 416620 243654 417240 243686
rect 416620 243418 416652 243654
rect 416888 243418 416972 243654
rect 417208 243418 417240 243654
rect 416620 243334 417240 243418
rect 416620 243098 416652 243334
rect 416888 243098 416972 243334
rect 417208 243098 417240 243334
rect 416620 243066 417240 243098
rect 452620 243654 453240 243686
rect 452620 243418 452652 243654
rect 452888 243418 452972 243654
rect 453208 243418 453240 243654
rect 452620 243334 453240 243418
rect 452620 243098 452652 243334
rect 452888 243098 452972 243334
rect 453208 243098 453240 243334
rect 452620 243066 453240 243098
rect 488620 243654 489240 243686
rect 488620 243418 488652 243654
rect 488888 243418 488972 243654
rect 489208 243418 489240 243654
rect 488620 243334 489240 243418
rect 488620 243098 488652 243334
rect 488888 243098 488972 243334
rect 489208 243098 489240 243334
rect 488620 243066 489240 243098
rect 524620 243654 525240 243686
rect 524620 243418 524652 243654
rect 524888 243418 524972 243654
rect 525208 243418 525240 243654
rect 524620 243334 525240 243418
rect 524620 243098 524652 243334
rect 524888 243098 524972 243334
rect 525208 243098 525240 243334
rect 524620 243066 525240 243098
rect 560620 243654 561240 243686
rect 560620 243418 560652 243654
rect 560888 243418 560972 243654
rect 561208 243418 561240 243654
rect 560620 243334 561240 243418
rect 560620 243098 560652 243334
rect 560888 243098 560972 243334
rect 561208 243098 561240 243334
rect 560620 243066 561240 243098
rect 570260 243654 570880 243686
rect 570260 243418 570292 243654
rect 570528 243418 570612 243654
rect 570848 243418 570880 243654
rect 570260 243334 570880 243418
rect 570260 243098 570292 243334
rect 570528 243098 570612 243334
rect 570848 243098 570880 243334
rect 570260 243066 570880 243098
rect 585310 243654 585930 283098
rect 585310 243418 585342 243654
rect 585578 243418 585662 243654
rect 585898 243418 585930 243654
rect 585310 243334 585930 243418
rect 585310 243098 585342 243334
rect 585578 243098 585662 243334
rect 585898 243098 585930 243334
rect 7844 223654 8464 223686
rect 7844 223418 7876 223654
rect 8112 223418 8196 223654
rect 8432 223418 8464 223654
rect 7844 223334 8464 223418
rect 7844 223098 7876 223334
rect 8112 223098 8196 223334
rect 8432 223098 8464 223334
rect 7844 223066 8464 223098
rect 38000 223654 38620 223686
rect 38000 223418 38032 223654
rect 38268 223418 38352 223654
rect 38588 223418 38620 223654
rect 38000 223334 38620 223418
rect 38000 223098 38032 223334
rect 38268 223098 38352 223334
rect 38588 223098 38620 223334
rect 38000 223066 38620 223098
rect 74000 223654 74620 223686
rect 74000 223418 74032 223654
rect 74268 223418 74352 223654
rect 74588 223418 74620 223654
rect 74000 223334 74620 223418
rect 74000 223098 74032 223334
rect 74268 223098 74352 223334
rect 74588 223098 74620 223334
rect 74000 223066 74620 223098
rect 110000 223654 110620 223686
rect 110000 223418 110032 223654
rect 110268 223418 110352 223654
rect 110588 223418 110620 223654
rect 110000 223334 110620 223418
rect 110000 223098 110032 223334
rect 110268 223098 110352 223334
rect 110588 223098 110620 223334
rect 110000 223066 110620 223098
rect 146000 223654 146620 223686
rect 146000 223418 146032 223654
rect 146268 223418 146352 223654
rect 146588 223418 146620 223654
rect 146000 223334 146620 223418
rect 146000 223098 146032 223334
rect 146268 223098 146352 223334
rect 146588 223098 146620 223334
rect 146000 223066 146620 223098
rect 182000 223654 182620 223686
rect 182000 223418 182032 223654
rect 182268 223418 182352 223654
rect 182588 223418 182620 223654
rect 182000 223334 182620 223418
rect 182000 223098 182032 223334
rect 182268 223098 182352 223334
rect 182588 223098 182620 223334
rect 182000 223066 182620 223098
rect 218000 223654 218620 223686
rect 218000 223418 218032 223654
rect 218268 223418 218352 223654
rect 218588 223418 218620 223654
rect 218000 223334 218620 223418
rect 218000 223098 218032 223334
rect 218268 223098 218352 223334
rect 218588 223098 218620 223334
rect 218000 223066 218620 223098
rect 254000 223654 254620 223686
rect 254000 223418 254032 223654
rect 254268 223418 254352 223654
rect 254588 223418 254620 223654
rect 254000 223334 254620 223418
rect 254000 223098 254032 223334
rect 254268 223098 254352 223334
rect 254588 223098 254620 223334
rect 254000 223066 254620 223098
rect 290000 223654 290620 223686
rect 290000 223418 290032 223654
rect 290268 223418 290352 223654
rect 290588 223418 290620 223654
rect 290000 223334 290620 223418
rect 290000 223098 290032 223334
rect 290268 223098 290352 223334
rect 290588 223098 290620 223334
rect 290000 223066 290620 223098
rect 326000 223654 326620 223686
rect 326000 223418 326032 223654
rect 326268 223418 326352 223654
rect 326588 223418 326620 223654
rect 326000 223334 326620 223418
rect 326000 223098 326032 223334
rect 326268 223098 326352 223334
rect 326588 223098 326620 223334
rect 326000 223066 326620 223098
rect 362000 223654 362620 223686
rect 362000 223418 362032 223654
rect 362268 223418 362352 223654
rect 362588 223418 362620 223654
rect 362000 223334 362620 223418
rect 362000 223098 362032 223334
rect 362268 223098 362352 223334
rect 362588 223098 362620 223334
rect 362000 223066 362620 223098
rect 398000 223654 398620 223686
rect 398000 223418 398032 223654
rect 398268 223418 398352 223654
rect 398588 223418 398620 223654
rect 398000 223334 398620 223418
rect 398000 223098 398032 223334
rect 398268 223098 398352 223334
rect 398588 223098 398620 223334
rect 398000 223066 398620 223098
rect 434000 223654 434620 223686
rect 434000 223418 434032 223654
rect 434268 223418 434352 223654
rect 434588 223418 434620 223654
rect 434000 223334 434620 223418
rect 434000 223098 434032 223334
rect 434268 223098 434352 223334
rect 434588 223098 434620 223334
rect 434000 223066 434620 223098
rect 470000 223654 470620 223686
rect 470000 223418 470032 223654
rect 470268 223418 470352 223654
rect 470588 223418 470620 223654
rect 470000 223334 470620 223418
rect 470000 223098 470032 223334
rect 470268 223098 470352 223334
rect 470588 223098 470620 223334
rect 470000 223066 470620 223098
rect 506000 223654 506620 223686
rect 506000 223418 506032 223654
rect 506268 223418 506352 223654
rect 506588 223418 506620 223654
rect 506000 223334 506620 223418
rect 506000 223098 506032 223334
rect 506268 223098 506352 223334
rect 506588 223098 506620 223334
rect 506000 223066 506620 223098
rect 542000 223654 542620 223686
rect 542000 223418 542032 223654
rect 542268 223418 542352 223654
rect 542588 223418 542620 223654
rect 542000 223334 542620 223418
rect 542000 223098 542032 223334
rect 542268 223098 542352 223334
rect 542588 223098 542620 223334
rect 542000 223066 542620 223098
rect 571500 223654 572120 223686
rect 571500 223418 571532 223654
rect 571768 223418 571852 223654
rect 572088 223418 572120 223654
rect 571500 223334 572120 223418
rect 571500 223098 571532 223334
rect 571768 223098 571852 223334
rect 572088 223098 572120 223334
rect 571500 223066 572120 223098
rect -2006 203418 -1974 203654
rect -1738 203418 -1654 203654
rect -1418 203418 -1386 203654
rect -2006 203334 -1386 203418
rect -2006 203098 -1974 203334
rect -1738 203098 -1654 203334
rect -1418 203098 -1386 203334
rect -2006 163654 -1386 203098
rect 9084 203654 9704 203686
rect 9084 203418 9116 203654
rect 9352 203418 9436 203654
rect 9672 203418 9704 203654
rect 9084 203334 9704 203418
rect 9084 203098 9116 203334
rect 9352 203098 9436 203334
rect 9672 203098 9704 203334
rect 9084 203066 9704 203098
rect 56620 203654 57240 203686
rect 56620 203418 56652 203654
rect 56888 203418 56972 203654
rect 57208 203418 57240 203654
rect 56620 203334 57240 203418
rect 56620 203098 56652 203334
rect 56888 203098 56972 203334
rect 57208 203098 57240 203334
rect 56620 203066 57240 203098
rect 92620 203654 93240 203686
rect 92620 203418 92652 203654
rect 92888 203418 92972 203654
rect 93208 203418 93240 203654
rect 92620 203334 93240 203418
rect 92620 203098 92652 203334
rect 92888 203098 92972 203334
rect 93208 203098 93240 203334
rect 92620 203066 93240 203098
rect 128620 203654 129240 203686
rect 128620 203418 128652 203654
rect 128888 203418 128972 203654
rect 129208 203418 129240 203654
rect 128620 203334 129240 203418
rect 128620 203098 128652 203334
rect 128888 203098 128972 203334
rect 129208 203098 129240 203334
rect 128620 203066 129240 203098
rect 164620 203654 165240 203686
rect 164620 203418 164652 203654
rect 164888 203418 164972 203654
rect 165208 203418 165240 203654
rect 164620 203334 165240 203418
rect 164620 203098 164652 203334
rect 164888 203098 164972 203334
rect 165208 203098 165240 203334
rect 164620 203066 165240 203098
rect 200620 203654 201240 203686
rect 200620 203418 200652 203654
rect 200888 203418 200972 203654
rect 201208 203418 201240 203654
rect 200620 203334 201240 203418
rect 200620 203098 200652 203334
rect 200888 203098 200972 203334
rect 201208 203098 201240 203334
rect 200620 203066 201240 203098
rect 236620 203654 237240 203686
rect 236620 203418 236652 203654
rect 236888 203418 236972 203654
rect 237208 203418 237240 203654
rect 236620 203334 237240 203418
rect 236620 203098 236652 203334
rect 236888 203098 236972 203334
rect 237208 203098 237240 203334
rect 236620 203066 237240 203098
rect 272620 203654 273240 203686
rect 272620 203418 272652 203654
rect 272888 203418 272972 203654
rect 273208 203418 273240 203654
rect 272620 203334 273240 203418
rect 272620 203098 272652 203334
rect 272888 203098 272972 203334
rect 273208 203098 273240 203334
rect 272620 203066 273240 203098
rect 308620 203654 309240 203686
rect 308620 203418 308652 203654
rect 308888 203418 308972 203654
rect 309208 203418 309240 203654
rect 308620 203334 309240 203418
rect 308620 203098 308652 203334
rect 308888 203098 308972 203334
rect 309208 203098 309240 203334
rect 308620 203066 309240 203098
rect 344620 203654 345240 203686
rect 344620 203418 344652 203654
rect 344888 203418 344972 203654
rect 345208 203418 345240 203654
rect 344620 203334 345240 203418
rect 344620 203098 344652 203334
rect 344888 203098 344972 203334
rect 345208 203098 345240 203334
rect 344620 203066 345240 203098
rect 380620 203654 381240 203686
rect 380620 203418 380652 203654
rect 380888 203418 380972 203654
rect 381208 203418 381240 203654
rect 380620 203334 381240 203418
rect 380620 203098 380652 203334
rect 380888 203098 380972 203334
rect 381208 203098 381240 203334
rect 380620 203066 381240 203098
rect 416620 203654 417240 203686
rect 416620 203418 416652 203654
rect 416888 203418 416972 203654
rect 417208 203418 417240 203654
rect 416620 203334 417240 203418
rect 416620 203098 416652 203334
rect 416888 203098 416972 203334
rect 417208 203098 417240 203334
rect 416620 203066 417240 203098
rect 452620 203654 453240 203686
rect 452620 203418 452652 203654
rect 452888 203418 452972 203654
rect 453208 203418 453240 203654
rect 452620 203334 453240 203418
rect 452620 203098 452652 203334
rect 452888 203098 452972 203334
rect 453208 203098 453240 203334
rect 452620 203066 453240 203098
rect 488620 203654 489240 203686
rect 488620 203418 488652 203654
rect 488888 203418 488972 203654
rect 489208 203418 489240 203654
rect 488620 203334 489240 203418
rect 488620 203098 488652 203334
rect 488888 203098 488972 203334
rect 489208 203098 489240 203334
rect 488620 203066 489240 203098
rect 524620 203654 525240 203686
rect 524620 203418 524652 203654
rect 524888 203418 524972 203654
rect 525208 203418 525240 203654
rect 524620 203334 525240 203418
rect 524620 203098 524652 203334
rect 524888 203098 524972 203334
rect 525208 203098 525240 203334
rect 524620 203066 525240 203098
rect 560620 203654 561240 203686
rect 560620 203418 560652 203654
rect 560888 203418 560972 203654
rect 561208 203418 561240 203654
rect 560620 203334 561240 203418
rect 560620 203098 560652 203334
rect 560888 203098 560972 203334
rect 561208 203098 561240 203334
rect 560620 203066 561240 203098
rect 570260 203654 570880 203686
rect 570260 203418 570292 203654
rect 570528 203418 570612 203654
rect 570848 203418 570880 203654
rect 570260 203334 570880 203418
rect 570260 203098 570292 203334
rect 570528 203098 570612 203334
rect 570848 203098 570880 203334
rect 570260 203066 570880 203098
rect 585310 203654 585930 243098
rect 585310 203418 585342 203654
rect 585578 203418 585662 203654
rect 585898 203418 585930 203654
rect 585310 203334 585930 203418
rect 585310 203098 585342 203334
rect 585578 203098 585662 203334
rect 585898 203098 585930 203334
rect 7844 183654 8464 183686
rect 7844 183418 7876 183654
rect 8112 183418 8196 183654
rect 8432 183418 8464 183654
rect 7844 183334 8464 183418
rect 7844 183098 7876 183334
rect 8112 183098 8196 183334
rect 8432 183098 8464 183334
rect 7844 183066 8464 183098
rect 38000 183654 38620 183686
rect 38000 183418 38032 183654
rect 38268 183418 38352 183654
rect 38588 183418 38620 183654
rect 38000 183334 38620 183418
rect 38000 183098 38032 183334
rect 38268 183098 38352 183334
rect 38588 183098 38620 183334
rect 38000 183066 38620 183098
rect 60560 183654 60920 183686
rect 60560 183418 60622 183654
rect 60858 183418 60920 183654
rect 60560 183334 60920 183418
rect 60560 183098 60622 183334
rect 60858 183098 60920 183334
rect 60560 183066 60920 183098
rect 159036 183654 159396 183686
rect 159036 183418 159098 183654
rect 159334 183418 159396 183654
rect 159036 183334 159396 183418
rect 159036 183098 159098 183334
rect 159334 183098 159396 183334
rect 159036 183066 159396 183098
rect 182000 183654 182620 183686
rect 182000 183418 182032 183654
rect 182268 183418 182352 183654
rect 182588 183418 182620 183654
rect 182000 183334 182620 183418
rect 182000 183098 182032 183334
rect 182268 183098 182352 183334
rect 182588 183098 182620 183334
rect 182000 183066 182620 183098
rect 185560 183654 185920 183686
rect 185560 183418 185622 183654
rect 185858 183418 185920 183654
rect 185560 183334 185920 183418
rect 185560 183098 185622 183334
rect 185858 183098 185920 183334
rect 185560 183066 185920 183098
rect 284036 183654 284396 183686
rect 284036 183418 284098 183654
rect 284334 183418 284396 183654
rect 284036 183334 284396 183418
rect 284036 183098 284098 183334
rect 284334 183098 284396 183334
rect 284036 183066 284396 183098
rect 290000 183654 290620 183686
rect 290000 183418 290032 183654
rect 290268 183418 290352 183654
rect 290588 183418 290620 183654
rect 290000 183334 290620 183418
rect 290000 183098 290032 183334
rect 290268 183098 290352 183334
rect 290588 183098 290620 183334
rect 290000 183066 290620 183098
rect 310560 183654 310920 183686
rect 310560 183418 310622 183654
rect 310858 183418 310920 183654
rect 310560 183334 310920 183418
rect 310560 183098 310622 183334
rect 310858 183098 310920 183334
rect 310560 183066 310920 183098
rect 409036 183654 409396 183686
rect 409036 183418 409098 183654
rect 409334 183418 409396 183654
rect 409036 183334 409396 183418
rect 409036 183098 409098 183334
rect 409334 183098 409396 183334
rect 409036 183066 409396 183098
rect 434000 183654 434620 183686
rect 434000 183418 434032 183654
rect 434268 183418 434352 183654
rect 434588 183418 434620 183654
rect 434000 183334 434620 183418
rect 434000 183098 434032 183334
rect 434268 183098 434352 183334
rect 434588 183098 434620 183334
rect 434000 183066 434620 183098
rect 436560 183654 436920 183686
rect 436560 183418 436622 183654
rect 436858 183418 436920 183654
rect 436560 183334 436920 183418
rect 436560 183098 436622 183334
rect 436858 183098 436920 183334
rect 436560 183066 436920 183098
rect 535036 183654 535396 183686
rect 535036 183418 535098 183654
rect 535334 183418 535396 183654
rect 535036 183334 535396 183418
rect 535036 183098 535098 183334
rect 535334 183098 535396 183334
rect 535036 183066 535396 183098
rect 542000 183654 542620 183686
rect 542000 183418 542032 183654
rect 542268 183418 542352 183654
rect 542588 183418 542620 183654
rect 542000 183334 542620 183418
rect 542000 183098 542032 183334
rect 542268 183098 542352 183334
rect 542588 183098 542620 183334
rect 542000 183066 542620 183098
rect 571500 183654 572120 183686
rect 571500 183418 571532 183654
rect 571768 183418 571852 183654
rect 572088 183418 572120 183654
rect 571500 183334 572120 183418
rect 571500 183098 571532 183334
rect 571768 183098 571852 183334
rect 572088 183098 572120 183334
rect 571500 183066 572120 183098
rect -2006 163418 -1974 163654
rect -1738 163418 -1654 163654
rect -1418 163418 -1386 163654
rect -2006 163334 -1386 163418
rect -2006 163098 -1974 163334
rect -1738 163098 -1654 163334
rect -1418 163098 -1386 163334
rect -2006 123654 -1386 163098
rect 9084 163654 9704 163686
rect 9084 163418 9116 163654
rect 9352 163418 9436 163654
rect 9672 163418 9704 163654
rect 9084 163334 9704 163418
rect 9084 163098 9116 163334
rect 9352 163098 9436 163334
rect 9672 163098 9704 163334
rect 9084 163066 9704 163098
rect 56620 163654 57240 163686
rect 56620 163418 56652 163654
rect 56888 163418 56972 163654
rect 57208 163418 57240 163654
rect 56620 163334 57240 163418
rect 56620 163098 56652 163334
rect 56888 163098 56972 163334
rect 57208 163098 57240 163334
rect 56620 163066 57240 163098
rect 61280 163654 61640 163686
rect 61280 163418 61342 163654
rect 61578 163418 61640 163654
rect 61280 163334 61640 163418
rect 61280 163098 61342 163334
rect 61578 163098 61640 163334
rect 61280 163066 61640 163098
rect 158316 163654 158676 163686
rect 158316 163418 158378 163654
rect 158614 163418 158676 163654
rect 158316 163334 158676 163418
rect 158316 163098 158378 163334
rect 158614 163098 158676 163334
rect 158316 163066 158676 163098
rect 164620 163654 165240 163686
rect 164620 163418 164652 163654
rect 164888 163418 164972 163654
rect 165208 163418 165240 163654
rect 164620 163334 165240 163418
rect 164620 163098 164652 163334
rect 164888 163098 164972 163334
rect 165208 163098 165240 163334
rect 164620 163066 165240 163098
rect 186280 163654 186640 163686
rect 186280 163418 186342 163654
rect 186578 163418 186640 163654
rect 186280 163334 186640 163418
rect 186280 163098 186342 163334
rect 186578 163098 186640 163334
rect 186280 163066 186640 163098
rect 283316 163654 283676 163686
rect 283316 163418 283378 163654
rect 283614 163418 283676 163654
rect 283316 163334 283676 163418
rect 283316 163098 283378 163334
rect 283614 163098 283676 163334
rect 283316 163066 283676 163098
rect 308620 163654 309240 163686
rect 308620 163418 308652 163654
rect 308888 163418 308972 163654
rect 309208 163418 309240 163654
rect 308620 163334 309240 163418
rect 308620 163098 308652 163334
rect 308888 163098 308972 163334
rect 309208 163098 309240 163334
rect 308620 163066 309240 163098
rect 311280 163654 311640 163686
rect 311280 163418 311342 163654
rect 311578 163418 311640 163654
rect 311280 163334 311640 163418
rect 311280 163098 311342 163334
rect 311578 163098 311640 163334
rect 311280 163066 311640 163098
rect 408316 163654 408676 163686
rect 408316 163418 408378 163654
rect 408614 163418 408676 163654
rect 408316 163334 408676 163418
rect 408316 163098 408378 163334
rect 408614 163098 408676 163334
rect 408316 163066 408676 163098
rect 416620 163654 417240 163686
rect 416620 163418 416652 163654
rect 416888 163418 416972 163654
rect 417208 163418 417240 163654
rect 416620 163334 417240 163418
rect 416620 163098 416652 163334
rect 416888 163098 416972 163334
rect 417208 163098 417240 163334
rect 416620 163066 417240 163098
rect 437280 163654 437640 163686
rect 437280 163418 437342 163654
rect 437578 163418 437640 163654
rect 437280 163334 437640 163418
rect 437280 163098 437342 163334
rect 437578 163098 437640 163334
rect 437280 163066 437640 163098
rect 534316 163654 534676 163686
rect 534316 163418 534378 163654
rect 534614 163418 534676 163654
rect 534316 163334 534676 163418
rect 534316 163098 534378 163334
rect 534614 163098 534676 163334
rect 534316 163066 534676 163098
rect 560620 163654 561240 163686
rect 560620 163418 560652 163654
rect 560888 163418 560972 163654
rect 561208 163418 561240 163654
rect 560620 163334 561240 163418
rect 560620 163098 560652 163334
rect 560888 163098 560972 163334
rect 561208 163098 561240 163334
rect 560620 163066 561240 163098
rect 570260 163654 570880 163686
rect 570260 163418 570292 163654
rect 570528 163418 570612 163654
rect 570848 163418 570880 163654
rect 570260 163334 570880 163418
rect 570260 163098 570292 163334
rect 570528 163098 570612 163334
rect 570848 163098 570880 163334
rect 570260 163066 570880 163098
rect 585310 163654 585930 203098
rect 585310 163418 585342 163654
rect 585578 163418 585662 163654
rect 585898 163418 585930 163654
rect 585310 163334 585930 163418
rect 585310 163098 585342 163334
rect 585578 163098 585662 163334
rect 585898 163098 585930 163334
rect 7844 143654 8464 143686
rect 7844 143418 7876 143654
rect 8112 143418 8196 143654
rect 8432 143418 8464 143654
rect 7844 143334 8464 143418
rect 7844 143098 7876 143334
rect 8112 143098 8196 143334
rect 8432 143098 8464 143334
rect 7844 143066 8464 143098
rect 38000 143654 38620 143686
rect 38000 143418 38032 143654
rect 38268 143418 38352 143654
rect 38588 143418 38620 143654
rect 38000 143334 38620 143418
rect 38000 143098 38032 143334
rect 38268 143098 38352 143334
rect 38588 143098 38620 143334
rect 38000 143066 38620 143098
rect 60560 143654 60920 143686
rect 60560 143418 60622 143654
rect 60858 143418 60920 143654
rect 60560 143334 60920 143418
rect 60560 143098 60622 143334
rect 60858 143098 60920 143334
rect 60560 143066 60920 143098
rect 159036 143654 159396 143686
rect 159036 143418 159098 143654
rect 159334 143418 159396 143654
rect 159036 143334 159396 143418
rect 159036 143098 159098 143334
rect 159334 143098 159396 143334
rect 159036 143066 159396 143098
rect 182000 143654 182620 143686
rect 182000 143418 182032 143654
rect 182268 143418 182352 143654
rect 182588 143418 182620 143654
rect 182000 143334 182620 143418
rect 182000 143098 182032 143334
rect 182268 143098 182352 143334
rect 182588 143098 182620 143334
rect 182000 143066 182620 143098
rect 185560 143654 185920 143686
rect 185560 143418 185622 143654
rect 185858 143418 185920 143654
rect 185560 143334 185920 143418
rect 185560 143098 185622 143334
rect 185858 143098 185920 143334
rect 185560 143066 185920 143098
rect 284036 143654 284396 143686
rect 284036 143418 284098 143654
rect 284334 143418 284396 143654
rect 284036 143334 284396 143418
rect 284036 143098 284098 143334
rect 284334 143098 284396 143334
rect 284036 143066 284396 143098
rect 290000 143654 290620 143686
rect 290000 143418 290032 143654
rect 290268 143418 290352 143654
rect 290588 143418 290620 143654
rect 290000 143334 290620 143418
rect 290000 143098 290032 143334
rect 290268 143098 290352 143334
rect 290588 143098 290620 143334
rect 290000 143066 290620 143098
rect 310560 143654 310920 143686
rect 310560 143418 310622 143654
rect 310858 143418 310920 143654
rect 310560 143334 310920 143418
rect 310560 143098 310622 143334
rect 310858 143098 310920 143334
rect 310560 143066 310920 143098
rect 409036 143654 409396 143686
rect 409036 143418 409098 143654
rect 409334 143418 409396 143654
rect 409036 143334 409396 143418
rect 409036 143098 409098 143334
rect 409334 143098 409396 143334
rect 409036 143066 409396 143098
rect 434000 143654 434620 143686
rect 434000 143418 434032 143654
rect 434268 143418 434352 143654
rect 434588 143418 434620 143654
rect 434000 143334 434620 143418
rect 434000 143098 434032 143334
rect 434268 143098 434352 143334
rect 434588 143098 434620 143334
rect 434000 143066 434620 143098
rect 436560 143654 436920 143686
rect 436560 143418 436622 143654
rect 436858 143418 436920 143654
rect 436560 143334 436920 143418
rect 436560 143098 436622 143334
rect 436858 143098 436920 143334
rect 436560 143066 436920 143098
rect 535036 143654 535396 143686
rect 535036 143418 535098 143654
rect 535334 143418 535396 143654
rect 535036 143334 535396 143418
rect 535036 143098 535098 143334
rect 535334 143098 535396 143334
rect 535036 143066 535396 143098
rect 542000 143654 542620 143686
rect 542000 143418 542032 143654
rect 542268 143418 542352 143654
rect 542588 143418 542620 143654
rect 542000 143334 542620 143418
rect 542000 143098 542032 143334
rect 542268 143098 542352 143334
rect 542588 143098 542620 143334
rect 542000 143066 542620 143098
rect 571500 143654 572120 143686
rect 571500 143418 571532 143654
rect 571768 143418 571852 143654
rect 572088 143418 572120 143654
rect 571500 143334 572120 143418
rect 571500 143098 571532 143334
rect 571768 143098 571852 143334
rect 572088 143098 572120 143334
rect 571500 143066 572120 143098
rect -2006 123418 -1974 123654
rect -1738 123418 -1654 123654
rect -1418 123418 -1386 123654
rect -2006 123334 -1386 123418
rect -2006 123098 -1974 123334
rect -1738 123098 -1654 123334
rect -1418 123098 -1386 123334
rect -2006 83654 -1386 123098
rect 9084 123654 9704 123686
rect 9084 123418 9116 123654
rect 9352 123418 9436 123654
rect 9672 123418 9704 123654
rect 9084 123334 9704 123418
rect 9084 123098 9116 123334
rect 9352 123098 9436 123334
rect 9672 123098 9704 123334
rect 9084 123066 9704 123098
rect 56620 123654 57240 123686
rect 56620 123418 56652 123654
rect 56888 123418 56972 123654
rect 57208 123418 57240 123654
rect 56620 123334 57240 123418
rect 56620 123098 56652 123334
rect 56888 123098 56972 123334
rect 57208 123098 57240 123334
rect 56620 123066 57240 123098
rect 61280 123654 61640 123686
rect 61280 123418 61342 123654
rect 61578 123418 61640 123654
rect 61280 123334 61640 123418
rect 61280 123098 61342 123334
rect 61578 123098 61640 123334
rect 61280 123066 61640 123098
rect 158316 123654 158676 123686
rect 158316 123418 158378 123654
rect 158614 123418 158676 123654
rect 158316 123334 158676 123418
rect 158316 123098 158378 123334
rect 158614 123098 158676 123334
rect 158316 123066 158676 123098
rect 164620 123654 165240 123686
rect 164620 123418 164652 123654
rect 164888 123418 164972 123654
rect 165208 123418 165240 123654
rect 164620 123334 165240 123418
rect 164620 123098 164652 123334
rect 164888 123098 164972 123334
rect 165208 123098 165240 123334
rect 164620 123066 165240 123098
rect 186280 123654 186640 123686
rect 186280 123418 186342 123654
rect 186578 123418 186640 123654
rect 186280 123334 186640 123418
rect 186280 123098 186342 123334
rect 186578 123098 186640 123334
rect 186280 123066 186640 123098
rect 283316 123654 283676 123686
rect 283316 123418 283378 123654
rect 283614 123418 283676 123654
rect 283316 123334 283676 123418
rect 283316 123098 283378 123334
rect 283614 123098 283676 123334
rect 283316 123066 283676 123098
rect 308620 123654 309240 123686
rect 308620 123418 308652 123654
rect 308888 123418 308972 123654
rect 309208 123418 309240 123654
rect 308620 123334 309240 123418
rect 308620 123098 308652 123334
rect 308888 123098 308972 123334
rect 309208 123098 309240 123334
rect 308620 123066 309240 123098
rect 311280 123654 311640 123686
rect 311280 123418 311342 123654
rect 311578 123418 311640 123654
rect 311280 123334 311640 123418
rect 311280 123098 311342 123334
rect 311578 123098 311640 123334
rect 311280 123066 311640 123098
rect 408316 123654 408676 123686
rect 408316 123418 408378 123654
rect 408614 123418 408676 123654
rect 408316 123334 408676 123418
rect 408316 123098 408378 123334
rect 408614 123098 408676 123334
rect 408316 123066 408676 123098
rect 416620 123654 417240 123686
rect 416620 123418 416652 123654
rect 416888 123418 416972 123654
rect 417208 123418 417240 123654
rect 416620 123334 417240 123418
rect 416620 123098 416652 123334
rect 416888 123098 416972 123334
rect 417208 123098 417240 123334
rect 416620 123066 417240 123098
rect 437280 123654 437640 123686
rect 437280 123418 437342 123654
rect 437578 123418 437640 123654
rect 437280 123334 437640 123418
rect 437280 123098 437342 123334
rect 437578 123098 437640 123334
rect 437280 123066 437640 123098
rect 534316 123654 534676 123686
rect 534316 123418 534378 123654
rect 534614 123418 534676 123654
rect 534316 123334 534676 123418
rect 534316 123098 534378 123334
rect 534614 123098 534676 123334
rect 534316 123066 534676 123098
rect 560620 123654 561240 123686
rect 560620 123418 560652 123654
rect 560888 123418 560972 123654
rect 561208 123418 561240 123654
rect 560620 123334 561240 123418
rect 560620 123098 560652 123334
rect 560888 123098 560972 123334
rect 561208 123098 561240 123334
rect 560620 123066 561240 123098
rect 570260 123654 570880 123686
rect 570260 123418 570292 123654
rect 570528 123418 570612 123654
rect 570848 123418 570880 123654
rect 570260 123334 570880 123418
rect 570260 123098 570292 123334
rect 570528 123098 570612 123334
rect 570848 123098 570880 123334
rect 570260 123066 570880 123098
rect 585310 123654 585930 163098
rect 585310 123418 585342 123654
rect 585578 123418 585662 123654
rect 585898 123418 585930 123654
rect 585310 123334 585930 123418
rect 585310 123098 585342 123334
rect 585578 123098 585662 123334
rect 585898 123098 585930 123334
rect 7844 103654 8464 103686
rect 7844 103418 7876 103654
rect 8112 103418 8196 103654
rect 8432 103418 8464 103654
rect 7844 103334 8464 103418
rect 7844 103098 7876 103334
rect 8112 103098 8196 103334
rect 8432 103098 8464 103334
rect 7844 103066 8464 103098
rect 38000 103654 38620 103686
rect 38000 103418 38032 103654
rect 38268 103418 38352 103654
rect 38588 103418 38620 103654
rect 38000 103334 38620 103418
rect 38000 103098 38032 103334
rect 38268 103098 38352 103334
rect 38588 103098 38620 103334
rect 38000 103066 38620 103098
rect 74000 103654 74620 103686
rect 74000 103418 74032 103654
rect 74268 103418 74352 103654
rect 74588 103418 74620 103654
rect 74000 103334 74620 103418
rect 74000 103098 74032 103334
rect 74268 103098 74352 103334
rect 74588 103098 74620 103334
rect 74000 103066 74620 103098
rect 110000 103654 110620 103686
rect 110000 103418 110032 103654
rect 110268 103418 110352 103654
rect 110588 103418 110620 103654
rect 110000 103334 110620 103418
rect 110000 103098 110032 103334
rect 110268 103098 110352 103334
rect 110588 103098 110620 103334
rect 110000 103066 110620 103098
rect 146000 103654 146620 103686
rect 146000 103418 146032 103654
rect 146268 103418 146352 103654
rect 146588 103418 146620 103654
rect 146000 103334 146620 103418
rect 146000 103098 146032 103334
rect 146268 103098 146352 103334
rect 146588 103098 146620 103334
rect 146000 103066 146620 103098
rect 182000 103654 182620 103686
rect 182000 103418 182032 103654
rect 182268 103418 182352 103654
rect 182588 103418 182620 103654
rect 182000 103334 182620 103418
rect 182000 103098 182032 103334
rect 182268 103098 182352 103334
rect 182588 103098 182620 103334
rect 182000 103066 182620 103098
rect 218000 103654 218620 103686
rect 218000 103418 218032 103654
rect 218268 103418 218352 103654
rect 218588 103418 218620 103654
rect 218000 103334 218620 103418
rect 218000 103098 218032 103334
rect 218268 103098 218352 103334
rect 218588 103098 218620 103334
rect 218000 103066 218620 103098
rect 254000 103654 254620 103686
rect 254000 103418 254032 103654
rect 254268 103418 254352 103654
rect 254588 103418 254620 103654
rect 254000 103334 254620 103418
rect 254000 103098 254032 103334
rect 254268 103098 254352 103334
rect 254588 103098 254620 103334
rect 254000 103066 254620 103098
rect 290000 103654 290620 103686
rect 290000 103418 290032 103654
rect 290268 103418 290352 103654
rect 290588 103418 290620 103654
rect 290000 103334 290620 103418
rect 290000 103098 290032 103334
rect 290268 103098 290352 103334
rect 290588 103098 290620 103334
rect 290000 103066 290620 103098
rect 326000 103654 326620 103686
rect 326000 103418 326032 103654
rect 326268 103418 326352 103654
rect 326588 103418 326620 103654
rect 326000 103334 326620 103418
rect 326000 103098 326032 103334
rect 326268 103098 326352 103334
rect 326588 103098 326620 103334
rect 326000 103066 326620 103098
rect 362000 103654 362620 103686
rect 362000 103418 362032 103654
rect 362268 103418 362352 103654
rect 362588 103418 362620 103654
rect 362000 103334 362620 103418
rect 362000 103098 362032 103334
rect 362268 103098 362352 103334
rect 362588 103098 362620 103334
rect 362000 103066 362620 103098
rect 398000 103654 398620 103686
rect 398000 103418 398032 103654
rect 398268 103418 398352 103654
rect 398588 103418 398620 103654
rect 398000 103334 398620 103418
rect 398000 103098 398032 103334
rect 398268 103098 398352 103334
rect 398588 103098 398620 103334
rect 398000 103066 398620 103098
rect 434000 103654 434620 103686
rect 434000 103418 434032 103654
rect 434268 103418 434352 103654
rect 434588 103418 434620 103654
rect 434000 103334 434620 103418
rect 434000 103098 434032 103334
rect 434268 103098 434352 103334
rect 434588 103098 434620 103334
rect 434000 103066 434620 103098
rect 470000 103654 470620 103686
rect 470000 103418 470032 103654
rect 470268 103418 470352 103654
rect 470588 103418 470620 103654
rect 470000 103334 470620 103418
rect 470000 103098 470032 103334
rect 470268 103098 470352 103334
rect 470588 103098 470620 103334
rect 470000 103066 470620 103098
rect 506000 103654 506620 103686
rect 506000 103418 506032 103654
rect 506268 103418 506352 103654
rect 506588 103418 506620 103654
rect 506000 103334 506620 103418
rect 506000 103098 506032 103334
rect 506268 103098 506352 103334
rect 506588 103098 506620 103334
rect 506000 103066 506620 103098
rect 542000 103654 542620 103686
rect 542000 103418 542032 103654
rect 542268 103418 542352 103654
rect 542588 103418 542620 103654
rect 542000 103334 542620 103418
rect 542000 103098 542032 103334
rect 542268 103098 542352 103334
rect 542588 103098 542620 103334
rect 542000 103066 542620 103098
rect 571500 103654 572120 103686
rect 571500 103418 571532 103654
rect 571768 103418 571852 103654
rect 572088 103418 572120 103654
rect 571500 103334 572120 103418
rect 571500 103098 571532 103334
rect 571768 103098 571852 103334
rect 572088 103098 572120 103334
rect 571500 103066 572120 103098
rect -2006 83418 -1974 83654
rect -1738 83418 -1654 83654
rect -1418 83418 -1386 83654
rect -2006 83334 -1386 83418
rect -2006 83098 -1974 83334
rect -1738 83098 -1654 83334
rect -1418 83098 -1386 83334
rect -2006 43654 -1386 83098
rect 9084 83654 9704 83686
rect 9084 83418 9116 83654
rect 9352 83418 9436 83654
rect 9672 83418 9704 83654
rect 9084 83334 9704 83418
rect 9084 83098 9116 83334
rect 9352 83098 9436 83334
rect 9672 83098 9704 83334
rect 9084 83066 9704 83098
rect 56620 83654 57240 83686
rect 56620 83418 56652 83654
rect 56888 83418 56972 83654
rect 57208 83418 57240 83654
rect 56620 83334 57240 83418
rect 56620 83098 56652 83334
rect 56888 83098 56972 83334
rect 57208 83098 57240 83334
rect 56620 83066 57240 83098
rect 61280 83654 61640 83686
rect 61280 83418 61342 83654
rect 61578 83418 61640 83654
rect 61280 83334 61640 83418
rect 61280 83098 61342 83334
rect 61578 83098 61640 83334
rect 61280 83066 61640 83098
rect 158316 83654 158676 83686
rect 158316 83418 158378 83654
rect 158614 83418 158676 83654
rect 158316 83334 158676 83418
rect 158316 83098 158378 83334
rect 158614 83098 158676 83334
rect 158316 83066 158676 83098
rect 164620 83654 165240 83686
rect 164620 83418 164652 83654
rect 164888 83418 164972 83654
rect 165208 83418 165240 83654
rect 164620 83334 165240 83418
rect 164620 83098 164652 83334
rect 164888 83098 164972 83334
rect 165208 83098 165240 83334
rect 164620 83066 165240 83098
rect 186280 83654 186640 83686
rect 186280 83418 186342 83654
rect 186578 83418 186640 83654
rect 186280 83334 186640 83418
rect 186280 83098 186342 83334
rect 186578 83098 186640 83334
rect 186280 83066 186640 83098
rect 283316 83654 283676 83686
rect 283316 83418 283378 83654
rect 283614 83418 283676 83654
rect 283316 83334 283676 83418
rect 283316 83098 283378 83334
rect 283614 83098 283676 83334
rect 283316 83066 283676 83098
rect 308620 83654 309240 83686
rect 308620 83418 308652 83654
rect 308888 83418 308972 83654
rect 309208 83418 309240 83654
rect 308620 83334 309240 83418
rect 308620 83098 308652 83334
rect 308888 83098 308972 83334
rect 309208 83098 309240 83334
rect 308620 83066 309240 83098
rect 311280 83654 311640 83686
rect 311280 83418 311342 83654
rect 311578 83418 311640 83654
rect 311280 83334 311640 83418
rect 311280 83098 311342 83334
rect 311578 83098 311640 83334
rect 311280 83066 311640 83098
rect 408316 83654 408676 83686
rect 408316 83418 408378 83654
rect 408614 83418 408676 83654
rect 408316 83334 408676 83418
rect 408316 83098 408378 83334
rect 408614 83098 408676 83334
rect 408316 83066 408676 83098
rect 416620 83654 417240 83686
rect 416620 83418 416652 83654
rect 416888 83418 416972 83654
rect 417208 83418 417240 83654
rect 416620 83334 417240 83418
rect 416620 83098 416652 83334
rect 416888 83098 416972 83334
rect 417208 83098 417240 83334
rect 416620 83066 417240 83098
rect 437280 83654 437640 83686
rect 437280 83418 437342 83654
rect 437578 83418 437640 83654
rect 437280 83334 437640 83418
rect 437280 83098 437342 83334
rect 437578 83098 437640 83334
rect 437280 83066 437640 83098
rect 534316 83654 534676 83686
rect 534316 83418 534378 83654
rect 534614 83418 534676 83654
rect 534316 83334 534676 83418
rect 534316 83098 534378 83334
rect 534614 83098 534676 83334
rect 534316 83066 534676 83098
rect 560620 83654 561240 83686
rect 560620 83418 560652 83654
rect 560888 83418 560972 83654
rect 561208 83418 561240 83654
rect 560620 83334 561240 83418
rect 560620 83098 560652 83334
rect 560888 83098 560972 83334
rect 561208 83098 561240 83334
rect 560620 83066 561240 83098
rect 570260 83654 570880 83686
rect 570260 83418 570292 83654
rect 570528 83418 570612 83654
rect 570848 83418 570880 83654
rect 570260 83334 570880 83418
rect 570260 83098 570292 83334
rect 570528 83098 570612 83334
rect 570848 83098 570880 83334
rect 570260 83066 570880 83098
rect 585310 83654 585930 123098
rect 585310 83418 585342 83654
rect 585578 83418 585662 83654
rect 585898 83418 585930 83654
rect 585310 83334 585930 83418
rect 585310 83098 585342 83334
rect 585578 83098 585662 83334
rect 585898 83098 585930 83334
rect 7844 63654 8464 63686
rect 7844 63418 7876 63654
rect 8112 63418 8196 63654
rect 8432 63418 8464 63654
rect 7844 63334 8464 63418
rect 7844 63098 7876 63334
rect 8112 63098 8196 63334
rect 8432 63098 8464 63334
rect 7844 63066 8464 63098
rect 38000 63654 38620 63686
rect 38000 63418 38032 63654
rect 38268 63418 38352 63654
rect 38588 63418 38620 63654
rect 38000 63334 38620 63418
rect 38000 63098 38032 63334
rect 38268 63098 38352 63334
rect 38588 63098 38620 63334
rect 38000 63066 38620 63098
rect 60560 63654 60920 63686
rect 60560 63418 60622 63654
rect 60858 63418 60920 63654
rect 60560 63334 60920 63418
rect 60560 63098 60622 63334
rect 60858 63098 60920 63334
rect 60560 63066 60920 63098
rect 159036 63654 159396 63686
rect 159036 63418 159098 63654
rect 159334 63418 159396 63654
rect 159036 63334 159396 63418
rect 159036 63098 159098 63334
rect 159334 63098 159396 63334
rect 159036 63066 159396 63098
rect 182000 63654 182620 63686
rect 182000 63418 182032 63654
rect 182268 63418 182352 63654
rect 182588 63418 182620 63654
rect 182000 63334 182620 63418
rect 182000 63098 182032 63334
rect 182268 63098 182352 63334
rect 182588 63098 182620 63334
rect 182000 63066 182620 63098
rect 185560 63654 185920 63686
rect 185560 63418 185622 63654
rect 185858 63418 185920 63654
rect 185560 63334 185920 63418
rect 185560 63098 185622 63334
rect 185858 63098 185920 63334
rect 185560 63066 185920 63098
rect 284036 63654 284396 63686
rect 284036 63418 284098 63654
rect 284334 63418 284396 63654
rect 284036 63334 284396 63418
rect 284036 63098 284098 63334
rect 284334 63098 284396 63334
rect 284036 63066 284396 63098
rect 290000 63654 290620 63686
rect 290000 63418 290032 63654
rect 290268 63418 290352 63654
rect 290588 63418 290620 63654
rect 290000 63334 290620 63418
rect 290000 63098 290032 63334
rect 290268 63098 290352 63334
rect 290588 63098 290620 63334
rect 290000 63066 290620 63098
rect 310560 63654 310920 63686
rect 310560 63418 310622 63654
rect 310858 63418 310920 63654
rect 310560 63334 310920 63418
rect 310560 63098 310622 63334
rect 310858 63098 310920 63334
rect 310560 63066 310920 63098
rect 409036 63654 409396 63686
rect 409036 63418 409098 63654
rect 409334 63418 409396 63654
rect 409036 63334 409396 63418
rect 409036 63098 409098 63334
rect 409334 63098 409396 63334
rect 409036 63066 409396 63098
rect 434000 63654 434620 63686
rect 434000 63418 434032 63654
rect 434268 63418 434352 63654
rect 434588 63418 434620 63654
rect 434000 63334 434620 63418
rect 434000 63098 434032 63334
rect 434268 63098 434352 63334
rect 434588 63098 434620 63334
rect 434000 63066 434620 63098
rect 436560 63654 436920 63686
rect 436560 63418 436622 63654
rect 436858 63418 436920 63654
rect 436560 63334 436920 63418
rect 436560 63098 436622 63334
rect 436858 63098 436920 63334
rect 436560 63066 436920 63098
rect 535036 63654 535396 63686
rect 535036 63418 535098 63654
rect 535334 63418 535396 63654
rect 535036 63334 535396 63418
rect 535036 63098 535098 63334
rect 535334 63098 535396 63334
rect 535036 63066 535396 63098
rect 542000 63654 542620 63686
rect 542000 63418 542032 63654
rect 542268 63418 542352 63654
rect 542588 63418 542620 63654
rect 542000 63334 542620 63418
rect 542000 63098 542032 63334
rect 542268 63098 542352 63334
rect 542588 63098 542620 63334
rect 542000 63066 542620 63098
rect 571500 63654 572120 63686
rect 571500 63418 571532 63654
rect 571768 63418 571852 63654
rect 572088 63418 572120 63654
rect 571500 63334 572120 63418
rect 571500 63098 571532 63334
rect 571768 63098 571852 63334
rect 572088 63098 572120 63334
rect 571500 63066 572120 63098
rect -2006 43418 -1974 43654
rect -1738 43418 -1654 43654
rect -1418 43418 -1386 43654
rect -2006 43334 -1386 43418
rect -2006 43098 -1974 43334
rect -1738 43098 -1654 43334
rect -1418 43098 -1386 43334
rect -2006 3654 -1386 43098
rect 9084 43654 9704 43686
rect 9084 43418 9116 43654
rect 9352 43418 9436 43654
rect 9672 43418 9704 43654
rect 9084 43334 9704 43418
rect 9084 43098 9116 43334
rect 9352 43098 9436 43334
rect 9672 43098 9704 43334
rect 9084 43066 9704 43098
rect 56620 43654 57240 43686
rect 56620 43418 56652 43654
rect 56888 43418 56972 43654
rect 57208 43418 57240 43654
rect 56620 43334 57240 43418
rect 56620 43098 56652 43334
rect 56888 43098 56972 43334
rect 57208 43098 57240 43334
rect 56620 43066 57240 43098
rect 61280 43654 61640 43686
rect 61280 43418 61342 43654
rect 61578 43418 61640 43654
rect 61280 43334 61640 43418
rect 61280 43098 61342 43334
rect 61578 43098 61640 43334
rect 61280 43066 61640 43098
rect 158316 43654 158676 43686
rect 158316 43418 158378 43654
rect 158614 43418 158676 43654
rect 158316 43334 158676 43418
rect 158316 43098 158378 43334
rect 158614 43098 158676 43334
rect 158316 43066 158676 43098
rect 164620 43654 165240 43686
rect 164620 43418 164652 43654
rect 164888 43418 164972 43654
rect 165208 43418 165240 43654
rect 164620 43334 165240 43418
rect 164620 43098 164652 43334
rect 164888 43098 164972 43334
rect 165208 43098 165240 43334
rect 164620 43066 165240 43098
rect 186280 43654 186640 43686
rect 186280 43418 186342 43654
rect 186578 43418 186640 43654
rect 186280 43334 186640 43418
rect 186280 43098 186342 43334
rect 186578 43098 186640 43334
rect 186280 43066 186640 43098
rect 283316 43654 283676 43686
rect 283316 43418 283378 43654
rect 283614 43418 283676 43654
rect 283316 43334 283676 43418
rect 283316 43098 283378 43334
rect 283614 43098 283676 43334
rect 283316 43066 283676 43098
rect 308620 43654 309240 43686
rect 308620 43418 308652 43654
rect 308888 43418 308972 43654
rect 309208 43418 309240 43654
rect 308620 43334 309240 43418
rect 308620 43098 308652 43334
rect 308888 43098 308972 43334
rect 309208 43098 309240 43334
rect 308620 43066 309240 43098
rect 311280 43654 311640 43686
rect 311280 43418 311342 43654
rect 311578 43418 311640 43654
rect 311280 43334 311640 43418
rect 311280 43098 311342 43334
rect 311578 43098 311640 43334
rect 311280 43066 311640 43098
rect 408316 43654 408676 43686
rect 408316 43418 408378 43654
rect 408614 43418 408676 43654
rect 408316 43334 408676 43418
rect 408316 43098 408378 43334
rect 408614 43098 408676 43334
rect 408316 43066 408676 43098
rect 416620 43654 417240 43686
rect 416620 43418 416652 43654
rect 416888 43418 416972 43654
rect 417208 43418 417240 43654
rect 416620 43334 417240 43418
rect 416620 43098 416652 43334
rect 416888 43098 416972 43334
rect 417208 43098 417240 43334
rect 416620 43066 417240 43098
rect 437280 43654 437640 43686
rect 437280 43418 437342 43654
rect 437578 43418 437640 43654
rect 437280 43334 437640 43418
rect 437280 43098 437342 43334
rect 437578 43098 437640 43334
rect 437280 43066 437640 43098
rect 534316 43654 534676 43686
rect 534316 43418 534378 43654
rect 534614 43418 534676 43654
rect 534316 43334 534676 43418
rect 534316 43098 534378 43334
rect 534614 43098 534676 43334
rect 534316 43066 534676 43098
rect 560620 43654 561240 43686
rect 560620 43418 560652 43654
rect 560888 43418 560972 43654
rect 561208 43418 561240 43654
rect 560620 43334 561240 43418
rect 560620 43098 560652 43334
rect 560888 43098 560972 43334
rect 561208 43098 561240 43334
rect 560620 43066 561240 43098
rect 570260 43654 570880 43686
rect 570260 43418 570292 43654
rect 570528 43418 570612 43654
rect 570848 43418 570880 43654
rect 570260 43334 570880 43418
rect 570260 43098 570292 43334
rect 570528 43098 570612 43334
rect 570848 43098 570880 43334
rect 570260 43066 570880 43098
rect 585310 43654 585930 83098
rect 585310 43418 585342 43654
rect 585578 43418 585662 43654
rect 585898 43418 585930 43654
rect 585310 43334 585930 43418
rect 585310 43098 585342 43334
rect 585578 43098 585662 43334
rect 585898 43098 585930 43334
rect 7844 23654 8464 23686
rect 7844 23418 7876 23654
rect 8112 23418 8196 23654
rect 8432 23418 8464 23654
rect 7844 23334 8464 23418
rect 7844 23098 7876 23334
rect 8112 23098 8196 23334
rect 8432 23098 8464 23334
rect 7844 23066 8464 23098
rect 38000 23654 38620 23686
rect 38000 23418 38032 23654
rect 38268 23418 38352 23654
rect 38588 23418 38620 23654
rect 38000 23334 38620 23418
rect 38000 23098 38032 23334
rect 38268 23098 38352 23334
rect 38588 23098 38620 23334
rect 38000 23066 38620 23098
rect 60560 23654 60920 23686
rect 60560 23418 60622 23654
rect 60858 23418 60920 23654
rect 60560 23334 60920 23418
rect 60560 23098 60622 23334
rect 60858 23098 60920 23334
rect 60560 23066 60920 23098
rect 159036 23654 159396 23686
rect 159036 23418 159098 23654
rect 159334 23418 159396 23654
rect 159036 23334 159396 23418
rect 159036 23098 159098 23334
rect 159334 23098 159396 23334
rect 159036 23066 159396 23098
rect 182000 23654 182620 23686
rect 182000 23418 182032 23654
rect 182268 23418 182352 23654
rect 182588 23418 182620 23654
rect 182000 23334 182620 23418
rect 182000 23098 182032 23334
rect 182268 23098 182352 23334
rect 182588 23098 182620 23334
rect 182000 23066 182620 23098
rect 185560 23654 185920 23686
rect 185560 23418 185622 23654
rect 185858 23418 185920 23654
rect 185560 23334 185920 23418
rect 185560 23098 185622 23334
rect 185858 23098 185920 23334
rect 185560 23066 185920 23098
rect 284036 23654 284396 23686
rect 284036 23418 284098 23654
rect 284334 23418 284396 23654
rect 284036 23334 284396 23418
rect 284036 23098 284098 23334
rect 284334 23098 284396 23334
rect 284036 23066 284396 23098
rect 290000 23654 290620 23686
rect 290000 23418 290032 23654
rect 290268 23418 290352 23654
rect 290588 23418 290620 23654
rect 290000 23334 290620 23418
rect 290000 23098 290032 23334
rect 290268 23098 290352 23334
rect 290588 23098 290620 23334
rect 290000 23066 290620 23098
rect 310560 23654 310920 23686
rect 310560 23418 310622 23654
rect 310858 23418 310920 23654
rect 310560 23334 310920 23418
rect 310560 23098 310622 23334
rect 310858 23098 310920 23334
rect 310560 23066 310920 23098
rect 409036 23654 409396 23686
rect 409036 23418 409098 23654
rect 409334 23418 409396 23654
rect 409036 23334 409396 23418
rect 409036 23098 409098 23334
rect 409334 23098 409396 23334
rect 409036 23066 409396 23098
rect 434000 23654 434620 23686
rect 434000 23418 434032 23654
rect 434268 23418 434352 23654
rect 434588 23418 434620 23654
rect 434000 23334 434620 23418
rect 434000 23098 434032 23334
rect 434268 23098 434352 23334
rect 434588 23098 434620 23334
rect 434000 23066 434620 23098
rect 436560 23654 436920 23686
rect 436560 23418 436622 23654
rect 436858 23418 436920 23654
rect 436560 23334 436920 23418
rect 436560 23098 436622 23334
rect 436858 23098 436920 23334
rect 436560 23066 436920 23098
rect 535036 23654 535396 23686
rect 535036 23418 535098 23654
rect 535334 23418 535396 23654
rect 535036 23334 535396 23418
rect 535036 23098 535098 23334
rect 535334 23098 535396 23334
rect 535036 23066 535396 23098
rect 542000 23654 542620 23686
rect 542000 23418 542032 23654
rect 542268 23418 542352 23654
rect 542588 23418 542620 23654
rect 542000 23334 542620 23418
rect 542000 23098 542032 23334
rect 542268 23098 542352 23334
rect 542588 23098 542620 23334
rect 542000 23066 542620 23098
rect 571500 23654 572120 23686
rect 571500 23418 571532 23654
rect 571768 23418 571852 23654
rect 572088 23418 572120 23654
rect 571500 23334 572120 23418
rect 571500 23098 571532 23334
rect 571768 23098 571852 23334
rect 572088 23098 572120 23334
rect 571500 23066 572120 23098
rect -2006 3418 -1974 3654
rect -1738 3418 -1654 3654
rect -1418 3418 -1386 3654
rect -2006 3334 -1386 3418
rect -2006 3098 -1974 3334
rect -1738 3098 -1654 3334
rect -1418 3098 -1386 3334
rect -2006 -346 -1386 3098
rect 585310 3654 585930 43098
rect 585310 3418 585342 3654
rect 585578 3418 585662 3654
rect 585898 3418 585930 3654
rect 585310 3334 585930 3418
rect 585310 3098 585342 3334
rect 585578 3098 585662 3334
rect 585898 3098 585930 3334
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1994 -346 2614 2000
rect 1994 -582 2026 -346
rect 2262 -582 2346 -346
rect 2582 -582 2614 -346
rect 1994 -666 2614 -582
rect 1994 -902 2026 -666
rect 2262 -902 2346 -666
rect 2582 -902 2614 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1994 -1894 2614 -902
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5714 -2266 6334 2000
rect 5714 -2502 5746 -2266
rect 5982 -2502 6066 -2266
rect 6302 -2502 6334 -2266
rect 5714 -2586 6334 -2502
rect 5714 -2822 5746 -2586
rect 5982 -2822 6066 -2586
rect 6302 -2822 6334 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5714 -3814 6334 -2822
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9434 -4186 10054 2000
rect 9434 -4422 9466 -4186
rect 9702 -4422 9786 -4186
rect 10022 -4422 10054 -4186
rect 9434 -4506 10054 -4422
rect 9434 -4742 9466 -4506
rect 9702 -4742 9786 -4506
rect 10022 -4742 10054 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9434 -5734 10054 -4742
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 13154 -6106 13774 2000
rect 21994 -1306 22614 2000
rect 21994 -1542 22026 -1306
rect 22262 -1542 22346 -1306
rect 22582 -1542 22614 -1306
rect 21994 -1626 22614 -1542
rect 21994 -1862 22026 -1626
rect 22262 -1862 22346 -1626
rect 22582 -1862 22614 -1626
rect 21994 -1894 22614 -1862
rect 25714 -3226 26334 2000
rect 25714 -3462 25746 -3226
rect 25982 -3462 26066 -3226
rect 26302 -3462 26334 -3226
rect 25714 -3546 26334 -3462
rect 25714 -3782 25746 -3546
rect 25982 -3782 26066 -3546
rect 26302 -3782 26334 -3546
rect 25714 -3814 26334 -3782
rect 29434 -5146 30054 2000
rect 29434 -5382 29466 -5146
rect 29702 -5382 29786 -5146
rect 30022 -5382 30054 -5146
rect 29434 -5466 30054 -5382
rect 29434 -5702 29466 -5466
rect 29702 -5702 29786 -5466
rect 30022 -5702 30054 -5466
rect 29434 -5734 30054 -5702
rect 13154 -6342 13186 -6106
rect 13422 -6342 13506 -6106
rect 13742 -6342 13774 -6106
rect 13154 -6426 13774 -6342
rect 13154 -6662 13186 -6426
rect 13422 -6662 13506 -6426
rect 13742 -6662 13774 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 13154 -7654 13774 -6662
rect 33154 -7066 33774 2000
rect 41994 -346 42614 2000
rect 41994 -582 42026 -346
rect 42262 -582 42346 -346
rect 42582 -582 42614 -346
rect 41994 -666 42614 -582
rect 41994 -902 42026 -666
rect 42262 -902 42346 -666
rect 42582 -902 42614 -666
rect 41994 -1894 42614 -902
rect 45714 -2266 46334 2000
rect 45714 -2502 45746 -2266
rect 45982 -2502 46066 -2266
rect 46302 -2502 46334 -2266
rect 45714 -2586 46334 -2502
rect 45714 -2822 45746 -2586
rect 45982 -2822 46066 -2586
rect 46302 -2822 46334 -2586
rect 45714 -3814 46334 -2822
rect 49434 -4186 50054 2000
rect 49434 -4422 49466 -4186
rect 49702 -4422 49786 -4186
rect 50022 -4422 50054 -4186
rect 49434 -4506 50054 -4422
rect 49434 -4742 49466 -4506
rect 49702 -4742 49786 -4506
rect 50022 -4742 50054 -4506
rect 49434 -5734 50054 -4742
rect 33154 -7302 33186 -7066
rect 33422 -7302 33506 -7066
rect 33742 -7302 33774 -7066
rect 33154 -7386 33774 -7302
rect 33154 -7622 33186 -7386
rect 33422 -7622 33506 -7386
rect 33742 -7622 33774 -7386
rect 33154 -7654 33774 -7622
rect 53154 -6106 53774 2000
rect 61994 -1306 62614 2000
rect 61994 -1542 62026 -1306
rect 62262 -1542 62346 -1306
rect 62582 -1542 62614 -1306
rect 61994 -1626 62614 -1542
rect 61994 -1862 62026 -1626
rect 62262 -1862 62346 -1626
rect 62582 -1862 62614 -1626
rect 61994 -1894 62614 -1862
rect 65714 -3226 66334 2000
rect 65714 -3462 65746 -3226
rect 65982 -3462 66066 -3226
rect 66302 -3462 66334 -3226
rect 65714 -3546 66334 -3462
rect 65714 -3782 65746 -3546
rect 65982 -3782 66066 -3546
rect 66302 -3782 66334 -3546
rect 65714 -3814 66334 -3782
rect 69434 -5146 70054 2000
rect 69434 -5382 69466 -5146
rect 69702 -5382 69786 -5146
rect 70022 -5382 70054 -5146
rect 69434 -5466 70054 -5382
rect 69434 -5702 69466 -5466
rect 69702 -5702 69786 -5466
rect 70022 -5702 70054 -5466
rect 69434 -5734 70054 -5702
rect 53154 -6342 53186 -6106
rect 53422 -6342 53506 -6106
rect 53742 -6342 53774 -6106
rect 53154 -6426 53774 -6342
rect 53154 -6662 53186 -6426
rect 53422 -6662 53506 -6426
rect 53742 -6662 53774 -6426
rect 53154 -7654 53774 -6662
rect 73154 -7066 73774 2000
rect 81994 -346 82614 2000
rect 81994 -582 82026 -346
rect 82262 -582 82346 -346
rect 82582 -582 82614 -346
rect 81994 -666 82614 -582
rect 81994 -902 82026 -666
rect 82262 -902 82346 -666
rect 82582 -902 82614 -666
rect 81994 -1894 82614 -902
rect 85714 -2266 86334 2000
rect 85714 -2502 85746 -2266
rect 85982 -2502 86066 -2266
rect 86302 -2502 86334 -2266
rect 85714 -2586 86334 -2502
rect 85714 -2822 85746 -2586
rect 85982 -2822 86066 -2586
rect 86302 -2822 86334 -2586
rect 85714 -3814 86334 -2822
rect 89434 -4186 90054 2000
rect 89434 -4422 89466 -4186
rect 89702 -4422 89786 -4186
rect 90022 -4422 90054 -4186
rect 89434 -4506 90054 -4422
rect 89434 -4742 89466 -4506
rect 89702 -4742 89786 -4506
rect 90022 -4742 90054 -4506
rect 89434 -5734 90054 -4742
rect 73154 -7302 73186 -7066
rect 73422 -7302 73506 -7066
rect 73742 -7302 73774 -7066
rect 73154 -7386 73774 -7302
rect 73154 -7622 73186 -7386
rect 73422 -7622 73506 -7386
rect 73742 -7622 73774 -7386
rect 73154 -7654 73774 -7622
rect 93154 -6106 93774 2000
rect 101994 -1306 102614 2000
rect 101994 -1542 102026 -1306
rect 102262 -1542 102346 -1306
rect 102582 -1542 102614 -1306
rect 101994 -1626 102614 -1542
rect 101994 -1862 102026 -1626
rect 102262 -1862 102346 -1626
rect 102582 -1862 102614 -1626
rect 101994 -1894 102614 -1862
rect 105714 -3226 106334 2000
rect 105714 -3462 105746 -3226
rect 105982 -3462 106066 -3226
rect 106302 -3462 106334 -3226
rect 105714 -3546 106334 -3462
rect 105714 -3782 105746 -3546
rect 105982 -3782 106066 -3546
rect 106302 -3782 106334 -3546
rect 105714 -3814 106334 -3782
rect 109434 -5146 110054 2000
rect 109434 -5382 109466 -5146
rect 109702 -5382 109786 -5146
rect 110022 -5382 110054 -5146
rect 109434 -5466 110054 -5382
rect 109434 -5702 109466 -5466
rect 109702 -5702 109786 -5466
rect 110022 -5702 110054 -5466
rect 109434 -5734 110054 -5702
rect 93154 -6342 93186 -6106
rect 93422 -6342 93506 -6106
rect 93742 -6342 93774 -6106
rect 93154 -6426 93774 -6342
rect 93154 -6662 93186 -6426
rect 93422 -6662 93506 -6426
rect 93742 -6662 93774 -6426
rect 93154 -7654 93774 -6662
rect 113154 -7066 113774 2000
rect 121994 -346 122614 2000
rect 121994 -582 122026 -346
rect 122262 -582 122346 -346
rect 122582 -582 122614 -346
rect 121994 -666 122614 -582
rect 121994 -902 122026 -666
rect 122262 -902 122346 -666
rect 122582 -902 122614 -666
rect 121994 -1894 122614 -902
rect 125714 -2266 126334 2000
rect 125714 -2502 125746 -2266
rect 125982 -2502 126066 -2266
rect 126302 -2502 126334 -2266
rect 125714 -2586 126334 -2502
rect 125714 -2822 125746 -2586
rect 125982 -2822 126066 -2586
rect 126302 -2822 126334 -2586
rect 125714 -3814 126334 -2822
rect 129434 -4186 130054 2000
rect 129434 -4422 129466 -4186
rect 129702 -4422 129786 -4186
rect 130022 -4422 130054 -4186
rect 129434 -4506 130054 -4422
rect 129434 -4742 129466 -4506
rect 129702 -4742 129786 -4506
rect 130022 -4742 130054 -4506
rect 129434 -5734 130054 -4742
rect 113154 -7302 113186 -7066
rect 113422 -7302 113506 -7066
rect 113742 -7302 113774 -7066
rect 113154 -7386 113774 -7302
rect 113154 -7622 113186 -7386
rect 113422 -7622 113506 -7386
rect 113742 -7622 113774 -7386
rect 113154 -7654 113774 -7622
rect 133154 -6106 133774 2000
rect 141994 -1306 142614 2000
rect 141994 -1542 142026 -1306
rect 142262 -1542 142346 -1306
rect 142582 -1542 142614 -1306
rect 141994 -1626 142614 -1542
rect 141994 -1862 142026 -1626
rect 142262 -1862 142346 -1626
rect 142582 -1862 142614 -1626
rect 141994 -1894 142614 -1862
rect 145714 -3226 146334 2000
rect 145714 -3462 145746 -3226
rect 145982 -3462 146066 -3226
rect 146302 -3462 146334 -3226
rect 145714 -3546 146334 -3462
rect 145714 -3782 145746 -3546
rect 145982 -3782 146066 -3546
rect 146302 -3782 146334 -3546
rect 145714 -3814 146334 -3782
rect 149434 -5146 150054 2000
rect 149434 -5382 149466 -5146
rect 149702 -5382 149786 -5146
rect 150022 -5382 150054 -5146
rect 149434 -5466 150054 -5382
rect 149434 -5702 149466 -5466
rect 149702 -5702 149786 -5466
rect 150022 -5702 150054 -5466
rect 149434 -5734 150054 -5702
rect 133154 -6342 133186 -6106
rect 133422 -6342 133506 -6106
rect 133742 -6342 133774 -6106
rect 133154 -6426 133774 -6342
rect 133154 -6662 133186 -6426
rect 133422 -6662 133506 -6426
rect 133742 -6662 133774 -6426
rect 133154 -7654 133774 -6662
rect 153154 -7066 153774 2000
rect 161994 -346 162614 2000
rect 161994 -582 162026 -346
rect 162262 -582 162346 -346
rect 162582 -582 162614 -346
rect 161994 -666 162614 -582
rect 161994 -902 162026 -666
rect 162262 -902 162346 -666
rect 162582 -902 162614 -666
rect 161994 -1894 162614 -902
rect 165714 -2266 166334 2000
rect 165714 -2502 165746 -2266
rect 165982 -2502 166066 -2266
rect 166302 -2502 166334 -2266
rect 165714 -2586 166334 -2502
rect 165714 -2822 165746 -2586
rect 165982 -2822 166066 -2586
rect 166302 -2822 166334 -2586
rect 165714 -3814 166334 -2822
rect 169434 -4186 170054 2000
rect 169434 -4422 169466 -4186
rect 169702 -4422 169786 -4186
rect 170022 -4422 170054 -4186
rect 169434 -4506 170054 -4422
rect 169434 -4742 169466 -4506
rect 169702 -4742 169786 -4506
rect 170022 -4742 170054 -4506
rect 169434 -5734 170054 -4742
rect 153154 -7302 153186 -7066
rect 153422 -7302 153506 -7066
rect 153742 -7302 153774 -7066
rect 153154 -7386 153774 -7302
rect 153154 -7622 153186 -7386
rect 153422 -7622 153506 -7386
rect 153742 -7622 153774 -7386
rect 153154 -7654 153774 -7622
rect 173154 -6106 173774 2000
rect 181994 -1306 182614 2000
rect 181994 -1542 182026 -1306
rect 182262 -1542 182346 -1306
rect 182582 -1542 182614 -1306
rect 181994 -1626 182614 -1542
rect 181994 -1862 182026 -1626
rect 182262 -1862 182346 -1626
rect 182582 -1862 182614 -1626
rect 181994 -1894 182614 -1862
rect 185714 -3226 186334 2000
rect 185714 -3462 185746 -3226
rect 185982 -3462 186066 -3226
rect 186302 -3462 186334 -3226
rect 185714 -3546 186334 -3462
rect 185714 -3782 185746 -3546
rect 185982 -3782 186066 -3546
rect 186302 -3782 186334 -3546
rect 185714 -3814 186334 -3782
rect 189434 -5146 190054 2000
rect 189434 -5382 189466 -5146
rect 189702 -5382 189786 -5146
rect 190022 -5382 190054 -5146
rect 189434 -5466 190054 -5382
rect 189434 -5702 189466 -5466
rect 189702 -5702 189786 -5466
rect 190022 -5702 190054 -5466
rect 189434 -5734 190054 -5702
rect 173154 -6342 173186 -6106
rect 173422 -6342 173506 -6106
rect 173742 -6342 173774 -6106
rect 173154 -6426 173774 -6342
rect 173154 -6662 173186 -6426
rect 173422 -6662 173506 -6426
rect 173742 -6662 173774 -6426
rect 173154 -7654 173774 -6662
rect 193154 -7066 193774 2000
rect 201994 -346 202614 2000
rect 201994 -582 202026 -346
rect 202262 -582 202346 -346
rect 202582 -582 202614 -346
rect 201994 -666 202614 -582
rect 201994 -902 202026 -666
rect 202262 -902 202346 -666
rect 202582 -902 202614 -666
rect 201994 -1894 202614 -902
rect 205714 -2266 206334 2000
rect 205714 -2502 205746 -2266
rect 205982 -2502 206066 -2266
rect 206302 -2502 206334 -2266
rect 205714 -2586 206334 -2502
rect 205714 -2822 205746 -2586
rect 205982 -2822 206066 -2586
rect 206302 -2822 206334 -2586
rect 205714 -3814 206334 -2822
rect 209434 -4186 210054 2000
rect 209434 -4422 209466 -4186
rect 209702 -4422 209786 -4186
rect 210022 -4422 210054 -4186
rect 209434 -4506 210054 -4422
rect 209434 -4742 209466 -4506
rect 209702 -4742 209786 -4506
rect 210022 -4742 210054 -4506
rect 209434 -5734 210054 -4742
rect 193154 -7302 193186 -7066
rect 193422 -7302 193506 -7066
rect 193742 -7302 193774 -7066
rect 193154 -7386 193774 -7302
rect 193154 -7622 193186 -7386
rect 193422 -7622 193506 -7386
rect 193742 -7622 193774 -7386
rect 193154 -7654 193774 -7622
rect 213154 -6106 213774 2000
rect 221994 -1306 222614 2000
rect 221994 -1542 222026 -1306
rect 222262 -1542 222346 -1306
rect 222582 -1542 222614 -1306
rect 221994 -1626 222614 -1542
rect 221994 -1862 222026 -1626
rect 222262 -1862 222346 -1626
rect 222582 -1862 222614 -1626
rect 221994 -1894 222614 -1862
rect 225714 -3226 226334 2000
rect 225714 -3462 225746 -3226
rect 225982 -3462 226066 -3226
rect 226302 -3462 226334 -3226
rect 225714 -3546 226334 -3462
rect 225714 -3782 225746 -3546
rect 225982 -3782 226066 -3546
rect 226302 -3782 226334 -3546
rect 225714 -3814 226334 -3782
rect 229434 -5146 230054 2000
rect 229434 -5382 229466 -5146
rect 229702 -5382 229786 -5146
rect 230022 -5382 230054 -5146
rect 229434 -5466 230054 -5382
rect 229434 -5702 229466 -5466
rect 229702 -5702 229786 -5466
rect 230022 -5702 230054 -5466
rect 229434 -5734 230054 -5702
rect 213154 -6342 213186 -6106
rect 213422 -6342 213506 -6106
rect 213742 -6342 213774 -6106
rect 213154 -6426 213774 -6342
rect 213154 -6662 213186 -6426
rect 213422 -6662 213506 -6426
rect 213742 -6662 213774 -6426
rect 213154 -7654 213774 -6662
rect 233154 -7066 233774 2000
rect 241994 -346 242614 2000
rect 241994 -582 242026 -346
rect 242262 -582 242346 -346
rect 242582 -582 242614 -346
rect 241994 -666 242614 -582
rect 241994 -902 242026 -666
rect 242262 -902 242346 -666
rect 242582 -902 242614 -666
rect 241994 -1894 242614 -902
rect 245714 -2266 246334 2000
rect 245714 -2502 245746 -2266
rect 245982 -2502 246066 -2266
rect 246302 -2502 246334 -2266
rect 245714 -2586 246334 -2502
rect 245714 -2822 245746 -2586
rect 245982 -2822 246066 -2586
rect 246302 -2822 246334 -2586
rect 245714 -3814 246334 -2822
rect 249434 -4186 250054 2000
rect 249434 -4422 249466 -4186
rect 249702 -4422 249786 -4186
rect 250022 -4422 250054 -4186
rect 249434 -4506 250054 -4422
rect 249434 -4742 249466 -4506
rect 249702 -4742 249786 -4506
rect 250022 -4742 250054 -4506
rect 249434 -5734 250054 -4742
rect 233154 -7302 233186 -7066
rect 233422 -7302 233506 -7066
rect 233742 -7302 233774 -7066
rect 233154 -7386 233774 -7302
rect 233154 -7622 233186 -7386
rect 233422 -7622 233506 -7386
rect 233742 -7622 233774 -7386
rect 233154 -7654 233774 -7622
rect 253154 -6106 253774 2000
rect 261994 -1306 262614 2000
rect 261994 -1542 262026 -1306
rect 262262 -1542 262346 -1306
rect 262582 -1542 262614 -1306
rect 261994 -1626 262614 -1542
rect 261994 -1862 262026 -1626
rect 262262 -1862 262346 -1626
rect 262582 -1862 262614 -1626
rect 261994 -1894 262614 -1862
rect 265714 -3226 266334 2000
rect 265714 -3462 265746 -3226
rect 265982 -3462 266066 -3226
rect 266302 -3462 266334 -3226
rect 265714 -3546 266334 -3462
rect 265714 -3782 265746 -3546
rect 265982 -3782 266066 -3546
rect 266302 -3782 266334 -3546
rect 265714 -3814 266334 -3782
rect 269434 -5146 270054 2000
rect 269434 -5382 269466 -5146
rect 269702 -5382 269786 -5146
rect 270022 -5382 270054 -5146
rect 269434 -5466 270054 -5382
rect 269434 -5702 269466 -5466
rect 269702 -5702 269786 -5466
rect 270022 -5702 270054 -5466
rect 269434 -5734 270054 -5702
rect 253154 -6342 253186 -6106
rect 253422 -6342 253506 -6106
rect 253742 -6342 253774 -6106
rect 253154 -6426 253774 -6342
rect 253154 -6662 253186 -6426
rect 253422 -6662 253506 -6426
rect 253742 -6662 253774 -6426
rect 253154 -7654 253774 -6662
rect 273154 -7066 273774 2000
rect 281994 -346 282614 2000
rect 281994 -582 282026 -346
rect 282262 -582 282346 -346
rect 282582 -582 282614 -346
rect 281994 -666 282614 -582
rect 281994 -902 282026 -666
rect 282262 -902 282346 -666
rect 282582 -902 282614 -666
rect 281994 -1894 282614 -902
rect 285714 -2266 286334 2000
rect 285714 -2502 285746 -2266
rect 285982 -2502 286066 -2266
rect 286302 -2502 286334 -2266
rect 285714 -2586 286334 -2502
rect 285714 -2822 285746 -2586
rect 285982 -2822 286066 -2586
rect 286302 -2822 286334 -2586
rect 285714 -3814 286334 -2822
rect 289434 -4186 290054 2000
rect 289434 -4422 289466 -4186
rect 289702 -4422 289786 -4186
rect 290022 -4422 290054 -4186
rect 289434 -4506 290054 -4422
rect 289434 -4742 289466 -4506
rect 289702 -4742 289786 -4506
rect 290022 -4742 290054 -4506
rect 289434 -5734 290054 -4742
rect 273154 -7302 273186 -7066
rect 273422 -7302 273506 -7066
rect 273742 -7302 273774 -7066
rect 273154 -7386 273774 -7302
rect 273154 -7622 273186 -7386
rect 273422 -7622 273506 -7386
rect 273742 -7622 273774 -7386
rect 273154 -7654 273774 -7622
rect 293154 -6106 293774 2000
rect 301994 -1306 302614 2000
rect 301994 -1542 302026 -1306
rect 302262 -1542 302346 -1306
rect 302582 -1542 302614 -1306
rect 301994 -1626 302614 -1542
rect 301994 -1862 302026 -1626
rect 302262 -1862 302346 -1626
rect 302582 -1862 302614 -1626
rect 301994 -1894 302614 -1862
rect 305714 -3226 306334 2000
rect 305714 -3462 305746 -3226
rect 305982 -3462 306066 -3226
rect 306302 -3462 306334 -3226
rect 305714 -3546 306334 -3462
rect 305714 -3782 305746 -3546
rect 305982 -3782 306066 -3546
rect 306302 -3782 306334 -3546
rect 305714 -3814 306334 -3782
rect 309434 -5146 310054 2000
rect 309434 -5382 309466 -5146
rect 309702 -5382 309786 -5146
rect 310022 -5382 310054 -5146
rect 309434 -5466 310054 -5382
rect 309434 -5702 309466 -5466
rect 309702 -5702 309786 -5466
rect 310022 -5702 310054 -5466
rect 309434 -5734 310054 -5702
rect 293154 -6342 293186 -6106
rect 293422 -6342 293506 -6106
rect 293742 -6342 293774 -6106
rect 293154 -6426 293774 -6342
rect 293154 -6662 293186 -6426
rect 293422 -6662 293506 -6426
rect 293742 -6662 293774 -6426
rect 293154 -7654 293774 -6662
rect 313154 -7066 313774 2000
rect 321994 -346 322614 2000
rect 321994 -582 322026 -346
rect 322262 -582 322346 -346
rect 322582 -582 322614 -346
rect 321994 -666 322614 -582
rect 321994 -902 322026 -666
rect 322262 -902 322346 -666
rect 322582 -902 322614 -666
rect 321994 -1894 322614 -902
rect 325714 -2266 326334 2000
rect 325714 -2502 325746 -2266
rect 325982 -2502 326066 -2266
rect 326302 -2502 326334 -2266
rect 325714 -2586 326334 -2502
rect 325714 -2822 325746 -2586
rect 325982 -2822 326066 -2586
rect 326302 -2822 326334 -2586
rect 325714 -3814 326334 -2822
rect 329434 -4186 330054 2000
rect 329434 -4422 329466 -4186
rect 329702 -4422 329786 -4186
rect 330022 -4422 330054 -4186
rect 329434 -4506 330054 -4422
rect 329434 -4742 329466 -4506
rect 329702 -4742 329786 -4506
rect 330022 -4742 330054 -4506
rect 329434 -5734 330054 -4742
rect 313154 -7302 313186 -7066
rect 313422 -7302 313506 -7066
rect 313742 -7302 313774 -7066
rect 313154 -7386 313774 -7302
rect 313154 -7622 313186 -7386
rect 313422 -7622 313506 -7386
rect 313742 -7622 313774 -7386
rect 313154 -7654 313774 -7622
rect 333154 -6106 333774 2000
rect 341994 -1306 342614 2000
rect 341994 -1542 342026 -1306
rect 342262 -1542 342346 -1306
rect 342582 -1542 342614 -1306
rect 341994 -1626 342614 -1542
rect 341994 -1862 342026 -1626
rect 342262 -1862 342346 -1626
rect 342582 -1862 342614 -1626
rect 341994 -1894 342614 -1862
rect 345714 -3226 346334 2000
rect 345714 -3462 345746 -3226
rect 345982 -3462 346066 -3226
rect 346302 -3462 346334 -3226
rect 345714 -3546 346334 -3462
rect 345714 -3782 345746 -3546
rect 345982 -3782 346066 -3546
rect 346302 -3782 346334 -3546
rect 345714 -3814 346334 -3782
rect 349434 -5146 350054 2000
rect 349434 -5382 349466 -5146
rect 349702 -5382 349786 -5146
rect 350022 -5382 350054 -5146
rect 349434 -5466 350054 -5382
rect 349434 -5702 349466 -5466
rect 349702 -5702 349786 -5466
rect 350022 -5702 350054 -5466
rect 349434 -5734 350054 -5702
rect 333154 -6342 333186 -6106
rect 333422 -6342 333506 -6106
rect 333742 -6342 333774 -6106
rect 333154 -6426 333774 -6342
rect 333154 -6662 333186 -6426
rect 333422 -6662 333506 -6426
rect 333742 -6662 333774 -6426
rect 333154 -7654 333774 -6662
rect 353154 -7066 353774 2000
rect 361994 -346 362614 2000
rect 361994 -582 362026 -346
rect 362262 -582 362346 -346
rect 362582 -582 362614 -346
rect 361994 -666 362614 -582
rect 361994 -902 362026 -666
rect 362262 -902 362346 -666
rect 362582 -902 362614 -666
rect 361994 -1894 362614 -902
rect 365714 -2266 366334 2000
rect 365714 -2502 365746 -2266
rect 365982 -2502 366066 -2266
rect 366302 -2502 366334 -2266
rect 365714 -2586 366334 -2502
rect 365714 -2822 365746 -2586
rect 365982 -2822 366066 -2586
rect 366302 -2822 366334 -2586
rect 365714 -3814 366334 -2822
rect 369434 -4186 370054 2000
rect 369434 -4422 369466 -4186
rect 369702 -4422 369786 -4186
rect 370022 -4422 370054 -4186
rect 369434 -4506 370054 -4422
rect 369434 -4742 369466 -4506
rect 369702 -4742 369786 -4506
rect 370022 -4742 370054 -4506
rect 369434 -5734 370054 -4742
rect 353154 -7302 353186 -7066
rect 353422 -7302 353506 -7066
rect 353742 -7302 353774 -7066
rect 353154 -7386 353774 -7302
rect 353154 -7622 353186 -7386
rect 353422 -7622 353506 -7386
rect 353742 -7622 353774 -7386
rect 353154 -7654 353774 -7622
rect 373154 -6106 373774 2000
rect 381994 -1306 382614 2000
rect 381994 -1542 382026 -1306
rect 382262 -1542 382346 -1306
rect 382582 -1542 382614 -1306
rect 381994 -1626 382614 -1542
rect 381994 -1862 382026 -1626
rect 382262 -1862 382346 -1626
rect 382582 -1862 382614 -1626
rect 381994 -1894 382614 -1862
rect 385714 -3226 386334 2000
rect 385714 -3462 385746 -3226
rect 385982 -3462 386066 -3226
rect 386302 -3462 386334 -3226
rect 385714 -3546 386334 -3462
rect 385714 -3782 385746 -3546
rect 385982 -3782 386066 -3546
rect 386302 -3782 386334 -3546
rect 385714 -3814 386334 -3782
rect 389434 -5146 390054 2000
rect 389434 -5382 389466 -5146
rect 389702 -5382 389786 -5146
rect 390022 -5382 390054 -5146
rect 389434 -5466 390054 -5382
rect 389434 -5702 389466 -5466
rect 389702 -5702 389786 -5466
rect 390022 -5702 390054 -5466
rect 389434 -5734 390054 -5702
rect 373154 -6342 373186 -6106
rect 373422 -6342 373506 -6106
rect 373742 -6342 373774 -6106
rect 373154 -6426 373774 -6342
rect 373154 -6662 373186 -6426
rect 373422 -6662 373506 -6426
rect 373742 -6662 373774 -6426
rect 373154 -7654 373774 -6662
rect 393154 -7066 393774 2000
rect 401994 -346 402614 2000
rect 401994 -582 402026 -346
rect 402262 -582 402346 -346
rect 402582 -582 402614 -346
rect 401994 -666 402614 -582
rect 401994 -902 402026 -666
rect 402262 -902 402346 -666
rect 402582 -902 402614 -666
rect 401994 -1894 402614 -902
rect 405714 -2266 406334 2000
rect 405714 -2502 405746 -2266
rect 405982 -2502 406066 -2266
rect 406302 -2502 406334 -2266
rect 405714 -2586 406334 -2502
rect 405714 -2822 405746 -2586
rect 405982 -2822 406066 -2586
rect 406302 -2822 406334 -2586
rect 405714 -3814 406334 -2822
rect 409434 -4186 410054 2000
rect 409434 -4422 409466 -4186
rect 409702 -4422 409786 -4186
rect 410022 -4422 410054 -4186
rect 409434 -4506 410054 -4422
rect 409434 -4742 409466 -4506
rect 409702 -4742 409786 -4506
rect 410022 -4742 410054 -4506
rect 409434 -5734 410054 -4742
rect 393154 -7302 393186 -7066
rect 393422 -7302 393506 -7066
rect 393742 -7302 393774 -7066
rect 393154 -7386 393774 -7302
rect 393154 -7622 393186 -7386
rect 393422 -7622 393506 -7386
rect 393742 -7622 393774 -7386
rect 393154 -7654 393774 -7622
rect 413154 -6106 413774 2000
rect 421994 -1306 422614 2000
rect 421994 -1542 422026 -1306
rect 422262 -1542 422346 -1306
rect 422582 -1542 422614 -1306
rect 421994 -1626 422614 -1542
rect 421994 -1862 422026 -1626
rect 422262 -1862 422346 -1626
rect 422582 -1862 422614 -1626
rect 421994 -1894 422614 -1862
rect 425714 -3226 426334 2000
rect 425714 -3462 425746 -3226
rect 425982 -3462 426066 -3226
rect 426302 -3462 426334 -3226
rect 425714 -3546 426334 -3462
rect 425714 -3782 425746 -3546
rect 425982 -3782 426066 -3546
rect 426302 -3782 426334 -3546
rect 425714 -3814 426334 -3782
rect 429434 -5146 430054 2000
rect 429434 -5382 429466 -5146
rect 429702 -5382 429786 -5146
rect 430022 -5382 430054 -5146
rect 429434 -5466 430054 -5382
rect 429434 -5702 429466 -5466
rect 429702 -5702 429786 -5466
rect 430022 -5702 430054 -5466
rect 429434 -5734 430054 -5702
rect 413154 -6342 413186 -6106
rect 413422 -6342 413506 -6106
rect 413742 -6342 413774 -6106
rect 413154 -6426 413774 -6342
rect 413154 -6662 413186 -6426
rect 413422 -6662 413506 -6426
rect 413742 -6662 413774 -6426
rect 413154 -7654 413774 -6662
rect 433154 -7066 433774 2000
rect 441994 -346 442614 2000
rect 441994 -582 442026 -346
rect 442262 -582 442346 -346
rect 442582 -582 442614 -346
rect 441994 -666 442614 -582
rect 441994 -902 442026 -666
rect 442262 -902 442346 -666
rect 442582 -902 442614 -666
rect 441994 -1894 442614 -902
rect 445714 -2266 446334 2000
rect 445714 -2502 445746 -2266
rect 445982 -2502 446066 -2266
rect 446302 -2502 446334 -2266
rect 445714 -2586 446334 -2502
rect 445714 -2822 445746 -2586
rect 445982 -2822 446066 -2586
rect 446302 -2822 446334 -2586
rect 445714 -3814 446334 -2822
rect 449434 -4186 450054 2000
rect 449434 -4422 449466 -4186
rect 449702 -4422 449786 -4186
rect 450022 -4422 450054 -4186
rect 449434 -4506 450054 -4422
rect 449434 -4742 449466 -4506
rect 449702 -4742 449786 -4506
rect 450022 -4742 450054 -4506
rect 449434 -5734 450054 -4742
rect 433154 -7302 433186 -7066
rect 433422 -7302 433506 -7066
rect 433742 -7302 433774 -7066
rect 433154 -7386 433774 -7302
rect 433154 -7622 433186 -7386
rect 433422 -7622 433506 -7386
rect 433742 -7622 433774 -7386
rect 433154 -7654 433774 -7622
rect 453154 -6106 453774 2000
rect 461994 -1306 462614 2000
rect 461994 -1542 462026 -1306
rect 462262 -1542 462346 -1306
rect 462582 -1542 462614 -1306
rect 461994 -1626 462614 -1542
rect 461994 -1862 462026 -1626
rect 462262 -1862 462346 -1626
rect 462582 -1862 462614 -1626
rect 461994 -1894 462614 -1862
rect 465714 -3226 466334 2000
rect 465714 -3462 465746 -3226
rect 465982 -3462 466066 -3226
rect 466302 -3462 466334 -3226
rect 465714 -3546 466334 -3462
rect 465714 -3782 465746 -3546
rect 465982 -3782 466066 -3546
rect 466302 -3782 466334 -3546
rect 465714 -3814 466334 -3782
rect 469434 -5146 470054 2000
rect 469434 -5382 469466 -5146
rect 469702 -5382 469786 -5146
rect 470022 -5382 470054 -5146
rect 469434 -5466 470054 -5382
rect 469434 -5702 469466 -5466
rect 469702 -5702 469786 -5466
rect 470022 -5702 470054 -5466
rect 469434 -5734 470054 -5702
rect 453154 -6342 453186 -6106
rect 453422 -6342 453506 -6106
rect 453742 -6342 453774 -6106
rect 453154 -6426 453774 -6342
rect 453154 -6662 453186 -6426
rect 453422 -6662 453506 -6426
rect 453742 -6662 453774 -6426
rect 453154 -7654 453774 -6662
rect 473154 -7066 473774 2000
rect 481994 -346 482614 2000
rect 481994 -582 482026 -346
rect 482262 -582 482346 -346
rect 482582 -582 482614 -346
rect 481994 -666 482614 -582
rect 481994 -902 482026 -666
rect 482262 -902 482346 -666
rect 482582 -902 482614 -666
rect 481994 -1894 482614 -902
rect 485714 -2266 486334 2000
rect 485714 -2502 485746 -2266
rect 485982 -2502 486066 -2266
rect 486302 -2502 486334 -2266
rect 485714 -2586 486334 -2502
rect 485714 -2822 485746 -2586
rect 485982 -2822 486066 -2586
rect 486302 -2822 486334 -2586
rect 485714 -3814 486334 -2822
rect 489434 -4186 490054 2000
rect 489434 -4422 489466 -4186
rect 489702 -4422 489786 -4186
rect 490022 -4422 490054 -4186
rect 489434 -4506 490054 -4422
rect 489434 -4742 489466 -4506
rect 489702 -4742 489786 -4506
rect 490022 -4742 490054 -4506
rect 489434 -5734 490054 -4742
rect 473154 -7302 473186 -7066
rect 473422 -7302 473506 -7066
rect 473742 -7302 473774 -7066
rect 473154 -7386 473774 -7302
rect 473154 -7622 473186 -7386
rect 473422 -7622 473506 -7386
rect 473742 -7622 473774 -7386
rect 473154 -7654 473774 -7622
rect 493154 -6106 493774 2000
rect 501994 -1306 502614 2000
rect 501994 -1542 502026 -1306
rect 502262 -1542 502346 -1306
rect 502582 -1542 502614 -1306
rect 501994 -1626 502614 -1542
rect 501994 -1862 502026 -1626
rect 502262 -1862 502346 -1626
rect 502582 -1862 502614 -1626
rect 501994 -1894 502614 -1862
rect 505714 -3226 506334 2000
rect 505714 -3462 505746 -3226
rect 505982 -3462 506066 -3226
rect 506302 -3462 506334 -3226
rect 505714 -3546 506334 -3462
rect 505714 -3782 505746 -3546
rect 505982 -3782 506066 -3546
rect 506302 -3782 506334 -3546
rect 505714 -3814 506334 -3782
rect 509434 -5146 510054 2000
rect 509434 -5382 509466 -5146
rect 509702 -5382 509786 -5146
rect 510022 -5382 510054 -5146
rect 509434 -5466 510054 -5382
rect 509434 -5702 509466 -5466
rect 509702 -5702 509786 -5466
rect 510022 -5702 510054 -5466
rect 509434 -5734 510054 -5702
rect 493154 -6342 493186 -6106
rect 493422 -6342 493506 -6106
rect 493742 -6342 493774 -6106
rect 493154 -6426 493774 -6342
rect 493154 -6662 493186 -6426
rect 493422 -6662 493506 -6426
rect 493742 -6662 493774 -6426
rect 493154 -7654 493774 -6662
rect 513154 -7066 513774 2000
rect 521994 -346 522614 2000
rect 521994 -582 522026 -346
rect 522262 -582 522346 -346
rect 522582 -582 522614 -346
rect 521994 -666 522614 -582
rect 521994 -902 522026 -666
rect 522262 -902 522346 -666
rect 522582 -902 522614 -666
rect 521994 -1894 522614 -902
rect 525714 -2266 526334 2000
rect 525714 -2502 525746 -2266
rect 525982 -2502 526066 -2266
rect 526302 -2502 526334 -2266
rect 525714 -2586 526334 -2502
rect 525714 -2822 525746 -2586
rect 525982 -2822 526066 -2586
rect 526302 -2822 526334 -2586
rect 525714 -3814 526334 -2822
rect 529434 -4186 530054 2000
rect 529434 -4422 529466 -4186
rect 529702 -4422 529786 -4186
rect 530022 -4422 530054 -4186
rect 529434 -4506 530054 -4422
rect 529434 -4742 529466 -4506
rect 529702 -4742 529786 -4506
rect 530022 -4742 530054 -4506
rect 529434 -5734 530054 -4742
rect 513154 -7302 513186 -7066
rect 513422 -7302 513506 -7066
rect 513742 -7302 513774 -7066
rect 513154 -7386 513774 -7302
rect 513154 -7622 513186 -7386
rect 513422 -7622 513506 -7386
rect 513742 -7622 513774 -7386
rect 513154 -7654 513774 -7622
rect 533154 -6106 533774 2000
rect 541994 -1306 542614 2000
rect 541994 -1542 542026 -1306
rect 542262 -1542 542346 -1306
rect 542582 -1542 542614 -1306
rect 541994 -1626 542614 -1542
rect 541994 -1862 542026 -1626
rect 542262 -1862 542346 -1626
rect 542582 -1862 542614 -1626
rect 541994 -1894 542614 -1862
rect 545714 -3226 546334 2000
rect 545714 -3462 545746 -3226
rect 545982 -3462 546066 -3226
rect 546302 -3462 546334 -3226
rect 545714 -3546 546334 -3462
rect 545714 -3782 545746 -3546
rect 545982 -3782 546066 -3546
rect 546302 -3782 546334 -3546
rect 545714 -3814 546334 -3782
rect 549434 -5146 550054 2000
rect 549434 -5382 549466 -5146
rect 549702 -5382 549786 -5146
rect 550022 -5382 550054 -5146
rect 549434 -5466 550054 -5382
rect 549434 -5702 549466 -5466
rect 549702 -5702 549786 -5466
rect 550022 -5702 550054 -5466
rect 549434 -5734 550054 -5702
rect 533154 -6342 533186 -6106
rect 533422 -6342 533506 -6106
rect 533742 -6342 533774 -6106
rect 533154 -6426 533774 -6342
rect 533154 -6662 533186 -6426
rect 533422 -6662 533506 -6426
rect 533742 -6662 533774 -6426
rect 533154 -7654 533774 -6662
rect 553154 -7066 553774 2000
rect 561994 -346 562614 2000
rect 561994 -582 562026 -346
rect 562262 -582 562346 -346
rect 562582 -582 562614 -346
rect 561994 -666 562614 -582
rect 561994 -902 562026 -666
rect 562262 -902 562346 -666
rect 562582 -902 562614 -666
rect 561994 -1894 562614 -902
rect 565714 -2266 566334 2000
rect 565714 -2502 565746 -2266
rect 565982 -2502 566066 -2266
rect 566302 -2502 566334 -2266
rect 565714 -2586 566334 -2502
rect 565714 -2822 565746 -2586
rect 565982 -2822 566066 -2586
rect 566302 -2822 566334 -2586
rect 565714 -3814 566334 -2822
rect 569434 -4186 570054 2000
rect 569434 -4422 569466 -4186
rect 569702 -4422 569786 -4186
rect 570022 -4422 570054 -4186
rect 569434 -4506 570054 -4422
rect 569434 -4742 569466 -4506
rect 569702 -4742 569786 -4506
rect 570022 -4742 570054 -4506
rect 569434 -5734 570054 -4742
rect 553154 -7302 553186 -7066
rect 553422 -7302 553506 -7066
rect 553742 -7302 553774 -7066
rect 553154 -7386 553774 -7302
rect 553154 -7622 553186 -7386
rect 553422 -7622 553506 -7386
rect 553742 -7622 553774 -7386
rect 553154 -7654 553774 -7622
rect 573154 -6106 573774 2000
rect 585310 -346 585930 3098
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 663654 586890 705242
rect 586270 663418 586302 663654
rect 586538 663418 586622 663654
rect 586858 663418 586890 663654
rect 586270 663334 586890 663418
rect 586270 663098 586302 663334
rect 586538 663098 586622 663334
rect 586858 663098 586890 663334
rect 586270 623654 586890 663098
rect 586270 623418 586302 623654
rect 586538 623418 586622 623654
rect 586858 623418 586890 623654
rect 586270 623334 586890 623418
rect 586270 623098 586302 623334
rect 586538 623098 586622 623334
rect 586858 623098 586890 623334
rect 586270 583654 586890 623098
rect 586270 583418 586302 583654
rect 586538 583418 586622 583654
rect 586858 583418 586890 583654
rect 586270 583334 586890 583418
rect 586270 583098 586302 583334
rect 586538 583098 586622 583334
rect 586858 583098 586890 583334
rect 586270 543654 586890 583098
rect 586270 543418 586302 543654
rect 586538 543418 586622 543654
rect 586858 543418 586890 543654
rect 586270 543334 586890 543418
rect 586270 543098 586302 543334
rect 586538 543098 586622 543334
rect 586858 543098 586890 543334
rect 586270 503654 586890 543098
rect 586270 503418 586302 503654
rect 586538 503418 586622 503654
rect 586858 503418 586890 503654
rect 586270 503334 586890 503418
rect 586270 503098 586302 503334
rect 586538 503098 586622 503334
rect 586858 503098 586890 503334
rect 586270 463654 586890 503098
rect 586270 463418 586302 463654
rect 586538 463418 586622 463654
rect 586858 463418 586890 463654
rect 586270 463334 586890 463418
rect 586270 463098 586302 463334
rect 586538 463098 586622 463334
rect 586858 463098 586890 463334
rect 586270 423654 586890 463098
rect 586270 423418 586302 423654
rect 586538 423418 586622 423654
rect 586858 423418 586890 423654
rect 586270 423334 586890 423418
rect 586270 423098 586302 423334
rect 586538 423098 586622 423334
rect 586858 423098 586890 423334
rect 586270 383654 586890 423098
rect 586270 383418 586302 383654
rect 586538 383418 586622 383654
rect 586858 383418 586890 383654
rect 586270 383334 586890 383418
rect 586270 383098 586302 383334
rect 586538 383098 586622 383334
rect 586858 383098 586890 383334
rect 586270 343654 586890 383098
rect 586270 343418 586302 343654
rect 586538 343418 586622 343654
rect 586858 343418 586890 343654
rect 586270 343334 586890 343418
rect 586270 343098 586302 343334
rect 586538 343098 586622 343334
rect 586858 343098 586890 343334
rect 586270 303654 586890 343098
rect 586270 303418 586302 303654
rect 586538 303418 586622 303654
rect 586858 303418 586890 303654
rect 586270 303334 586890 303418
rect 586270 303098 586302 303334
rect 586538 303098 586622 303334
rect 586858 303098 586890 303334
rect 586270 263654 586890 303098
rect 586270 263418 586302 263654
rect 586538 263418 586622 263654
rect 586858 263418 586890 263654
rect 586270 263334 586890 263418
rect 586270 263098 586302 263334
rect 586538 263098 586622 263334
rect 586858 263098 586890 263334
rect 586270 223654 586890 263098
rect 586270 223418 586302 223654
rect 586538 223418 586622 223654
rect 586858 223418 586890 223654
rect 586270 223334 586890 223418
rect 586270 223098 586302 223334
rect 586538 223098 586622 223334
rect 586858 223098 586890 223334
rect 586270 183654 586890 223098
rect 586270 183418 586302 183654
rect 586538 183418 586622 183654
rect 586858 183418 586890 183654
rect 586270 183334 586890 183418
rect 586270 183098 586302 183334
rect 586538 183098 586622 183334
rect 586858 183098 586890 183334
rect 586270 143654 586890 183098
rect 586270 143418 586302 143654
rect 586538 143418 586622 143654
rect 586858 143418 586890 143654
rect 586270 143334 586890 143418
rect 586270 143098 586302 143334
rect 586538 143098 586622 143334
rect 586858 143098 586890 143334
rect 586270 103654 586890 143098
rect 586270 103418 586302 103654
rect 586538 103418 586622 103654
rect 586858 103418 586890 103654
rect 586270 103334 586890 103418
rect 586270 103098 586302 103334
rect 586538 103098 586622 103334
rect 586858 103098 586890 103334
rect 586270 63654 586890 103098
rect 586270 63418 586302 63654
rect 586538 63418 586622 63654
rect 586858 63418 586890 63654
rect 586270 63334 586890 63418
rect 586270 63098 586302 63334
rect 586538 63098 586622 63334
rect 586858 63098 586890 63334
rect 586270 23654 586890 63098
rect 586270 23418 586302 23654
rect 586538 23418 586622 23654
rect 586858 23418 586890 23654
rect 586270 23334 586890 23418
rect 586270 23098 586302 23334
rect 586538 23098 586622 23334
rect 586858 23098 586890 23334
rect 586270 -1306 586890 23098
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 687374 587850 706202
rect 587230 687138 587262 687374
rect 587498 687138 587582 687374
rect 587818 687138 587850 687374
rect 587230 687054 587850 687138
rect 587230 686818 587262 687054
rect 587498 686818 587582 687054
rect 587818 686818 587850 687054
rect 587230 647374 587850 686818
rect 587230 647138 587262 647374
rect 587498 647138 587582 647374
rect 587818 647138 587850 647374
rect 587230 647054 587850 647138
rect 587230 646818 587262 647054
rect 587498 646818 587582 647054
rect 587818 646818 587850 647054
rect 587230 607374 587850 646818
rect 587230 607138 587262 607374
rect 587498 607138 587582 607374
rect 587818 607138 587850 607374
rect 587230 607054 587850 607138
rect 587230 606818 587262 607054
rect 587498 606818 587582 607054
rect 587818 606818 587850 607054
rect 587230 567374 587850 606818
rect 587230 567138 587262 567374
rect 587498 567138 587582 567374
rect 587818 567138 587850 567374
rect 587230 567054 587850 567138
rect 587230 566818 587262 567054
rect 587498 566818 587582 567054
rect 587818 566818 587850 567054
rect 587230 527374 587850 566818
rect 587230 527138 587262 527374
rect 587498 527138 587582 527374
rect 587818 527138 587850 527374
rect 587230 527054 587850 527138
rect 587230 526818 587262 527054
rect 587498 526818 587582 527054
rect 587818 526818 587850 527054
rect 587230 487374 587850 526818
rect 587230 487138 587262 487374
rect 587498 487138 587582 487374
rect 587818 487138 587850 487374
rect 587230 487054 587850 487138
rect 587230 486818 587262 487054
rect 587498 486818 587582 487054
rect 587818 486818 587850 487054
rect 587230 447374 587850 486818
rect 587230 447138 587262 447374
rect 587498 447138 587582 447374
rect 587818 447138 587850 447374
rect 587230 447054 587850 447138
rect 587230 446818 587262 447054
rect 587498 446818 587582 447054
rect 587818 446818 587850 447054
rect 587230 407374 587850 446818
rect 587230 407138 587262 407374
rect 587498 407138 587582 407374
rect 587818 407138 587850 407374
rect 587230 407054 587850 407138
rect 587230 406818 587262 407054
rect 587498 406818 587582 407054
rect 587818 406818 587850 407054
rect 587230 367374 587850 406818
rect 587230 367138 587262 367374
rect 587498 367138 587582 367374
rect 587818 367138 587850 367374
rect 587230 367054 587850 367138
rect 587230 366818 587262 367054
rect 587498 366818 587582 367054
rect 587818 366818 587850 367054
rect 587230 327374 587850 366818
rect 587230 327138 587262 327374
rect 587498 327138 587582 327374
rect 587818 327138 587850 327374
rect 587230 327054 587850 327138
rect 587230 326818 587262 327054
rect 587498 326818 587582 327054
rect 587818 326818 587850 327054
rect 587230 287374 587850 326818
rect 587230 287138 587262 287374
rect 587498 287138 587582 287374
rect 587818 287138 587850 287374
rect 587230 287054 587850 287138
rect 587230 286818 587262 287054
rect 587498 286818 587582 287054
rect 587818 286818 587850 287054
rect 587230 247374 587850 286818
rect 587230 247138 587262 247374
rect 587498 247138 587582 247374
rect 587818 247138 587850 247374
rect 587230 247054 587850 247138
rect 587230 246818 587262 247054
rect 587498 246818 587582 247054
rect 587818 246818 587850 247054
rect 587230 207374 587850 246818
rect 587230 207138 587262 207374
rect 587498 207138 587582 207374
rect 587818 207138 587850 207374
rect 587230 207054 587850 207138
rect 587230 206818 587262 207054
rect 587498 206818 587582 207054
rect 587818 206818 587850 207054
rect 587230 167374 587850 206818
rect 587230 167138 587262 167374
rect 587498 167138 587582 167374
rect 587818 167138 587850 167374
rect 587230 167054 587850 167138
rect 587230 166818 587262 167054
rect 587498 166818 587582 167054
rect 587818 166818 587850 167054
rect 587230 127374 587850 166818
rect 587230 127138 587262 127374
rect 587498 127138 587582 127374
rect 587818 127138 587850 127374
rect 587230 127054 587850 127138
rect 587230 126818 587262 127054
rect 587498 126818 587582 127054
rect 587818 126818 587850 127054
rect 587230 87374 587850 126818
rect 587230 87138 587262 87374
rect 587498 87138 587582 87374
rect 587818 87138 587850 87374
rect 587230 87054 587850 87138
rect 587230 86818 587262 87054
rect 587498 86818 587582 87054
rect 587818 86818 587850 87054
rect 587230 47374 587850 86818
rect 587230 47138 587262 47374
rect 587498 47138 587582 47374
rect 587818 47138 587850 47374
rect 587230 47054 587850 47138
rect 587230 46818 587262 47054
rect 587498 46818 587582 47054
rect 587818 46818 587850 47054
rect 587230 7374 587850 46818
rect 587230 7138 587262 7374
rect 587498 7138 587582 7374
rect 587818 7138 587850 7374
rect 587230 7054 587850 7138
rect 587230 6818 587262 7054
rect 587498 6818 587582 7054
rect 587818 6818 587850 7054
rect 587230 -2266 587850 6818
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 667374 588810 707162
rect 588190 667138 588222 667374
rect 588458 667138 588542 667374
rect 588778 667138 588810 667374
rect 588190 667054 588810 667138
rect 588190 666818 588222 667054
rect 588458 666818 588542 667054
rect 588778 666818 588810 667054
rect 588190 627374 588810 666818
rect 588190 627138 588222 627374
rect 588458 627138 588542 627374
rect 588778 627138 588810 627374
rect 588190 627054 588810 627138
rect 588190 626818 588222 627054
rect 588458 626818 588542 627054
rect 588778 626818 588810 627054
rect 588190 587374 588810 626818
rect 588190 587138 588222 587374
rect 588458 587138 588542 587374
rect 588778 587138 588810 587374
rect 588190 587054 588810 587138
rect 588190 586818 588222 587054
rect 588458 586818 588542 587054
rect 588778 586818 588810 587054
rect 588190 547374 588810 586818
rect 588190 547138 588222 547374
rect 588458 547138 588542 547374
rect 588778 547138 588810 547374
rect 588190 547054 588810 547138
rect 588190 546818 588222 547054
rect 588458 546818 588542 547054
rect 588778 546818 588810 547054
rect 588190 507374 588810 546818
rect 588190 507138 588222 507374
rect 588458 507138 588542 507374
rect 588778 507138 588810 507374
rect 588190 507054 588810 507138
rect 588190 506818 588222 507054
rect 588458 506818 588542 507054
rect 588778 506818 588810 507054
rect 588190 467374 588810 506818
rect 588190 467138 588222 467374
rect 588458 467138 588542 467374
rect 588778 467138 588810 467374
rect 588190 467054 588810 467138
rect 588190 466818 588222 467054
rect 588458 466818 588542 467054
rect 588778 466818 588810 467054
rect 588190 427374 588810 466818
rect 588190 427138 588222 427374
rect 588458 427138 588542 427374
rect 588778 427138 588810 427374
rect 588190 427054 588810 427138
rect 588190 426818 588222 427054
rect 588458 426818 588542 427054
rect 588778 426818 588810 427054
rect 588190 387374 588810 426818
rect 588190 387138 588222 387374
rect 588458 387138 588542 387374
rect 588778 387138 588810 387374
rect 588190 387054 588810 387138
rect 588190 386818 588222 387054
rect 588458 386818 588542 387054
rect 588778 386818 588810 387054
rect 588190 347374 588810 386818
rect 588190 347138 588222 347374
rect 588458 347138 588542 347374
rect 588778 347138 588810 347374
rect 588190 347054 588810 347138
rect 588190 346818 588222 347054
rect 588458 346818 588542 347054
rect 588778 346818 588810 347054
rect 588190 307374 588810 346818
rect 588190 307138 588222 307374
rect 588458 307138 588542 307374
rect 588778 307138 588810 307374
rect 588190 307054 588810 307138
rect 588190 306818 588222 307054
rect 588458 306818 588542 307054
rect 588778 306818 588810 307054
rect 588190 267374 588810 306818
rect 588190 267138 588222 267374
rect 588458 267138 588542 267374
rect 588778 267138 588810 267374
rect 588190 267054 588810 267138
rect 588190 266818 588222 267054
rect 588458 266818 588542 267054
rect 588778 266818 588810 267054
rect 588190 227374 588810 266818
rect 588190 227138 588222 227374
rect 588458 227138 588542 227374
rect 588778 227138 588810 227374
rect 588190 227054 588810 227138
rect 588190 226818 588222 227054
rect 588458 226818 588542 227054
rect 588778 226818 588810 227054
rect 588190 187374 588810 226818
rect 588190 187138 588222 187374
rect 588458 187138 588542 187374
rect 588778 187138 588810 187374
rect 588190 187054 588810 187138
rect 588190 186818 588222 187054
rect 588458 186818 588542 187054
rect 588778 186818 588810 187054
rect 588190 147374 588810 186818
rect 588190 147138 588222 147374
rect 588458 147138 588542 147374
rect 588778 147138 588810 147374
rect 588190 147054 588810 147138
rect 588190 146818 588222 147054
rect 588458 146818 588542 147054
rect 588778 146818 588810 147054
rect 588190 107374 588810 146818
rect 588190 107138 588222 107374
rect 588458 107138 588542 107374
rect 588778 107138 588810 107374
rect 588190 107054 588810 107138
rect 588190 106818 588222 107054
rect 588458 106818 588542 107054
rect 588778 106818 588810 107054
rect 588190 67374 588810 106818
rect 588190 67138 588222 67374
rect 588458 67138 588542 67374
rect 588778 67138 588810 67374
rect 588190 67054 588810 67138
rect 588190 66818 588222 67054
rect 588458 66818 588542 67054
rect 588778 66818 588810 67054
rect 588190 27374 588810 66818
rect 588190 27138 588222 27374
rect 588458 27138 588542 27374
rect 588778 27138 588810 27374
rect 588190 27054 588810 27138
rect 588190 26818 588222 27054
rect 588458 26818 588542 27054
rect 588778 26818 588810 27054
rect 588190 -3226 588810 26818
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 691094 589770 708122
rect 589150 690858 589182 691094
rect 589418 690858 589502 691094
rect 589738 690858 589770 691094
rect 589150 690774 589770 690858
rect 589150 690538 589182 690774
rect 589418 690538 589502 690774
rect 589738 690538 589770 690774
rect 589150 651094 589770 690538
rect 589150 650858 589182 651094
rect 589418 650858 589502 651094
rect 589738 650858 589770 651094
rect 589150 650774 589770 650858
rect 589150 650538 589182 650774
rect 589418 650538 589502 650774
rect 589738 650538 589770 650774
rect 589150 611094 589770 650538
rect 589150 610858 589182 611094
rect 589418 610858 589502 611094
rect 589738 610858 589770 611094
rect 589150 610774 589770 610858
rect 589150 610538 589182 610774
rect 589418 610538 589502 610774
rect 589738 610538 589770 610774
rect 589150 571094 589770 610538
rect 589150 570858 589182 571094
rect 589418 570858 589502 571094
rect 589738 570858 589770 571094
rect 589150 570774 589770 570858
rect 589150 570538 589182 570774
rect 589418 570538 589502 570774
rect 589738 570538 589770 570774
rect 589150 531094 589770 570538
rect 589150 530858 589182 531094
rect 589418 530858 589502 531094
rect 589738 530858 589770 531094
rect 589150 530774 589770 530858
rect 589150 530538 589182 530774
rect 589418 530538 589502 530774
rect 589738 530538 589770 530774
rect 589150 491094 589770 530538
rect 589150 490858 589182 491094
rect 589418 490858 589502 491094
rect 589738 490858 589770 491094
rect 589150 490774 589770 490858
rect 589150 490538 589182 490774
rect 589418 490538 589502 490774
rect 589738 490538 589770 490774
rect 589150 451094 589770 490538
rect 589150 450858 589182 451094
rect 589418 450858 589502 451094
rect 589738 450858 589770 451094
rect 589150 450774 589770 450858
rect 589150 450538 589182 450774
rect 589418 450538 589502 450774
rect 589738 450538 589770 450774
rect 589150 411094 589770 450538
rect 589150 410858 589182 411094
rect 589418 410858 589502 411094
rect 589738 410858 589770 411094
rect 589150 410774 589770 410858
rect 589150 410538 589182 410774
rect 589418 410538 589502 410774
rect 589738 410538 589770 410774
rect 589150 371094 589770 410538
rect 589150 370858 589182 371094
rect 589418 370858 589502 371094
rect 589738 370858 589770 371094
rect 589150 370774 589770 370858
rect 589150 370538 589182 370774
rect 589418 370538 589502 370774
rect 589738 370538 589770 370774
rect 589150 331094 589770 370538
rect 589150 330858 589182 331094
rect 589418 330858 589502 331094
rect 589738 330858 589770 331094
rect 589150 330774 589770 330858
rect 589150 330538 589182 330774
rect 589418 330538 589502 330774
rect 589738 330538 589770 330774
rect 589150 291094 589770 330538
rect 589150 290858 589182 291094
rect 589418 290858 589502 291094
rect 589738 290858 589770 291094
rect 589150 290774 589770 290858
rect 589150 290538 589182 290774
rect 589418 290538 589502 290774
rect 589738 290538 589770 290774
rect 589150 251094 589770 290538
rect 589150 250858 589182 251094
rect 589418 250858 589502 251094
rect 589738 250858 589770 251094
rect 589150 250774 589770 250858
rect 589150 250538 589182 250774
rect 589418 250538 589502 250774
rect 589738 250538 589770 250774
rect 589150 211094 589770 250538
rect 589150 210858 589182 211094
rect 589418 210858 589502 211094
rect 589738 210858 589770 211094
rect 589150 210774 589770 210858
rect 589150 210538 589182 210774
rect 589418 210538 589502 210774
rect 589738 210538 589770 210774
rect 589150 171094 589770 210538
rect 589150 170858 589182 171094
rect 589418 170858 589502 171094
rect 589738 170858 589770 171094
rect 589150 170774 589770 170858
rect 589150 170538 589182 170774
rect 589418 170538 589502 170774
rect 589738 170538 589770 170774
rect 589150 131094 589770 170538
rect 589150 130858 589182 131094
rect 589418 130858 589502 131094
rect 589738 130858 589770 131094
rect 589150 130774 589770 130858
rect 589150 130538 589182 130774
rect 589418 130538 589502 130774
rect 589738 130538 589770 130774
rect 589150 91094 589770 130538
rect 589150 90858 589182 91094
rect 589418 90858 589502 91094
rect 589738 90858 589770 91094
rect 589150 90774 589770 90858
rect 589150 90538 589182 90774
rect 589418 90538 589502 90774
rect 589738 90538 589770 90774
rect 589150 51094 589770 90538
rect 589150 50858 589182 51094
rect 589418 50858 589502 51094
rect 589738 50858 589770 51094
rect 589150 50774 589770 50858
rect 589150 50538 589182 50774
rect 589418 50538 589502 50774
rect 589738 50538 589770 50774
rect 589150 11094 589770 50538
rect 589150 10858 589182 11094
rect 589418 10858 589502 11094
rect 589738 10858 589770 11094
rect 589150 10774 589770 10858
rect 589150 10538 589182 10774
rect 589418 10538 589502 10774
rect 589738 10538 589770 10774
rect 589150 -4186 589770 10538
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 671094 590730 709082
rect 590110 670858 590142 671094
rect 590378 670858 590462 671094
rect 590698 670858 590730 671094
rect 590110 670774 590730 670858
rect 590110 670538 590142 670774
rect 590378 670538 590462 670774
rect 590698 670538 590730 670774
rect 590110 631094 590730 670538
rect 590110 630858 590142 631094
rect 590378 630858 590462 631094
rect 590698 630858 590730 631094
rect 590110 630774 590730 630858
rect 590110 630538 590142 630774
rect 590378 630538 590462 630774
rect 590698 630538 590730 630774
rect 590110 591094 590730 630538
rect 590110 590858 590142 591094
rect 590378 590858 590462 591094
rect 590698 590858 590730 591094
rect 590110 590774 590730 590858
rect 590110 590538 590142 590774
rect 590378 590538 590462 590774
rect 590698 590538 590730 590774
rect 590110 551094 590730 590538
rect 590110 550858 590142 551094
rect 590378 550858 590462 551094
rect 590698 550858 590730 551094
rect 590110 550774 590730 550858
rect 590110 550538 590142 550774
rect 590378 550538 590462 550774
rect 590698 550538 590730 550774
rect 590110 511094 590730 550538
rect 590110 510858 590142 511094
rect 590378 510858 590462 511094
rect 590698 510858 590730 511094
rect 590110 510774 590730 510858
rect 590110 510538 590142 510774
rect 590378 510538 590462 510774
rect 590698 510538 590730 510774
rect 590110 471094 590730 510538
rect 590110 470858 590142 471094
rect 590378 470858 590462 471094
rect 590698 470858 590730 471094
rect 590110 470774 590730 470858
rect 590110 470538 590142 470774
rect 590378 470538 590462 470774
rect 590698 470538 590730 470774
rect 590110 431094 590730 470538
rect 590110 430858 590142 431094
rect 590378 430858 590462 431094
rect 590698 430858 590730 431094
rect 590110 430774 590730 430858
rect 590110 430538 590142 430774
rect 590378 430538 590462 430774
rect 590698 430538 590730 430774
rect 590110 391094 590730 430538
rect 590110 390858 590142 391094
rect 590378 390858 590462 391094
rect 590698 390858 590730 391094
rect 590110 390774 590730 390858
rect 590110 390538 590142 390774
rect 590378 390538 590462 390774
rect 590698 390538 590730 390774
rect 590110 351094 590730 390538
rect 590110 350858 590142 351094
rect 590378 350858 590462 351094
rect 590698 350858 590730 351094
rect 590110 350774 590730 350858
rect 590110 350538 590142 350774
rect 590378 350538 590462 350774
rect 590698 350538 590730 350774
rect 590110 311094 590730 350538
rect 590110 310858 590142 311094
rect 590378 310858 590462 311094
rect 590698 310858 590730 311094
rect 590110 310774 590730 310858
rect 590110 310538 590142 310774
rect 590378 310538 590462 310774
rect 590698 310538 590730 310774
rect 590110 271094 590730 310538
rect 590110 270858 590142 271094
rect 590378 270858 590462 271094
rect 590698 270858 590730 271094
rect 590110 270774 590730 270858
rect 590110 270538 590142 270774
rect 590378 270538 590462 270774
rect 590698 270538 590730 270774
rect 590110 231094 590730 270538
rect 590110 230858 590142 231094
rect 590378 230858 590462 231094
rect 590698 230858 590730 231094
rect 590110 230774 590730 230858
rect 590110 230538 590142 230774
rect 590378 230538 590462 230774
rect 590698 230538 590730 230774
rect 590110 191094 590730 230538
rect 590110 190858 590142 191094
rect 590378 190858 590462 191094
rect 590698 190858 590730 191094
rect 590110 190774 590730 190858
rect 590110 190538 590142 190774
rect 590378 190538 590462 190774
rect 590698 190538 590730 190774
rect 590110 151094 590730 190538
rect 590110 150858 590142 151094
rect 590378 150858 590462 151094
rect 590698 150858 590730 151094
rect 590110 150774 590730 150858
rect 590110 150538 590142 150774
rect 590378 150538 590462 150774
rect 590698 150538 590730 150774
rect 590110 111094 590730 150538
rect 590110 110858 590142 111094
rect 590378 110858 590462 111094
rect 590698 110858 590730 111094
rect 590110 110774 590730 110858
rect 590110 110538 590142 110774
rect 590378 110538 590462 110774
rect 590698 110538 590730 110774
rect 590110 71094 590730 110538
rect 590110 70858 590142 71094
rect 590378 70858 590462 71094
rect 590698 70858 590730 71094
rect 590110 70774 590730 70858
rect 590110 70538 590142 70774
rect 590378 70538 590462 70774
rect 590698 70538 590730 70774
rect 590110 31094 590730 70538
rect 590110 30858 590142 31094
rect 590378 30858 590462 31094
rect 590698 30858 590730 31094
rect 590110 30774 590730 30858
rect 590110 30538 590142 30774
rect 590378 30538 590462 30774
rect 590698 30538 590730 30774
rect 590110 -5146 590730 30538
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 694814 591690 710042
rect 591070 694578 591102 694814
rect 591338 694578 591422 694814
rect 591658 694578 591690 694814
rect 591070 694494 591690 694578
rect 591070 694258 591102 694494
rect 591338 694258 591422 694494
rect 591658 694258 591690 694494
rect 591070 654814 591690 694258
rect 591070 654578 591102 654814
rect 591338 654578 591422 654814
rect 591658 654578 591690 654814
rect 591070 654494 591690 654578
rect 591070 654258 591102 654494
rect 591338 654258 591422 654494
rect 591658 654258 591690 654494
rect 591070 614814 591690 654258
rect 591070 614578 591102 614814
rect 591338 614578 591422 614814
rect 591658 614578 591690 614814
rect 591070 614494 591690 614578
rect 591070 614258 591102 614494
rect 591338 614258 591422 614494
rect 591658 614258 591690 614494
rect 591070 574814 591690 614258
rect 591070 574578 591102 574814
rect 591338 574578 591422 574814
rect 591658 574578 591690 574814
rect 591070 574494 591690 574578
rect 591070 574258 591102 574494
rect 591338 574258 591422 574494
rect 591658 574258 591690 574494
rect 591070 534814 591690 574258
rect 591070 534578 591102 534814
rect 591338 534578 591422 534814
rect 591658 534578 591690 534814
rect 591070 534494 591690 534578
rect 591070 534258 591102 534494
rect 591338 534258 591422 534494
rect 591658 534258 591690 534494
rect 591070 494814 591690 534258
rect 591070 494578 591102 494814
rect 591338 494578 591422 494814
rect 591658 494578 591690 494814
rect 591070 494494 591690 494578
rect 591070 494258 591102 494494
rect 591338 494258 591422 494494
rect 591658 494258 591690 494494
rect 591070 454814 591690 494258
rect 591070 454578 591102 454814
rect 591338 454578 591422 454814
rect 591658 454578 591690 454814
rect 591070 454494 591690 454578
rect 591070 454258 591102 454494
rect 591338 454258 591422 454494
rect 591658 454258 591690 454494
rect 591070 414814 591690 454258
rect 591070 414578 591102 414814
rect 591338 414578 591422 414814
rect 591658 414578 591690 414814
rect 591070 414494 591690 414578
rect 591070 414258 591102 414494
rect 591338 414258 591422 414494
rect 591658 414258 591690 414494
rect 591070 374814 591690 414258
rect 591070 374578 591102 374814
rect 591338 374578 591422 374814
rect 591658 374578 591690 374814
rect 591070 374494 591690 374578
rect 591070 374258 591102 374494
rect 591338 374258 591422 374494
rect 591658 374258 591690 374494
rect 591070 334814 591690 374258
rect 591070 334578 591102 334814
rect 591338 334578 591422 334814
rect 591658 334578 591690 334814
rect 591070 334494 591690 334578
rect 591070 334258 591102 334494
rect 591338 334258 591422 334494
rect 591658 334258 591690 334494
rect 591070 294814 591690 334258
rect 591070 294578 591102 294814
rect 591338 294578 591422 294814
rect 591658 294578 591690 294814
rect 591070 294494 591690 294578
rect 591070 294258 591102 294494
rect 591338 294258 591422 294494
rect 591658 294258 591690 294494
rect 591070 254814 591690 294258
rect 591070 254578 591102 254814
rect 591338 254578 591422 254814
rect 591658 254578 591690 254814
rect 591070 254494 591690 254578
rect 591070 254258 591102 254494
rect 591338 254258 591422 254494
rect 591658 254258 591690 254494
rect 591070 214814 591690 254258
rect 591070 214578 591102 214814
rect 591338 214578 591422 214814
rect 591658 214578 591690 214814
rect 591070 214494 591690 214578
rect 591070 214258 591102 214494
rect 591338 214258 591422 214494
rect 591658 214258 591690 214494
rect 591070 174814 591690 214258
rect 591070 174578 591102 174814
rect 591338 174578 591422 174814
rect 591658 174578 591690 174814
rect 591070 174494 591690 174578
rect 591070 174258 591102 174494
rect 591338 174258 591422 174494
rect 591658 174258 591690 174494
rect 591070 134814 591690 174258
rect 591070 134578 591102 134814
rect 591338 134578 591422 134814
rect 591658 134578 591690 134814
rect 591070 134494 591690 134578
rect 591070 134258 591102 134494
rect 591338 134258 591422 134494
rect 591658 134258 591690 134494
rect 591070 94814 591690 134258
rect 591070 94578 591102 94814
rect 591338 94578 591422 94814
rect 591658 94578 591690 94814
rect 591070 94494 591690 94578
rect 591070 94258 591102 94494
rect 591338 94258 591422 94494
rect 591658 94258 591690 94494
rect 591070 54814 591690 94258
rect 591070 54578 591102 54814
rect 591338 54578 591422 54814
rect 591658 54578 591690 54814
rect 591070 54494 591690 54578
rect 591070 54258 591102 54494
rect 591338 54258 591422 54494
rect 591658 54258 591690 54494
rect 591070 14814 591690 54258
rect 591070 14578 591102 14814
rect 591338 14578 591422 14814
rect 591658 14578 591690 14814
rect 591070 14494 591690 14578
rect 591070 14258 591102 14494
rect 591338 14258 591422 14494
rect 591658 14258 591690 14494
rect 573154 -6342 573186 -6106
rect 573422 -6342 573506 -6106
rect 573742 -6342 573774 -6106
rect 573154 -6426 573774 -6342
rect 573154 -6662 573186 -6426
rect 573422 -6662 573506 -6426
rect 573742 -6662 573774 -6426
rect 573154 -7654 573774 -6662
rect 591070 -6106 591690 14258
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 674814 592650 711002
rect 592030 674578 592062 674814
rect 592298 674578 592382 674814
rect 592618 674578 592650 674814
rect 592030 674494 592650 674578
rect 592030 674258 592062 674494
rect 592298 674258 592382 674494
rect 592618 674258 592650 674494
rect 592030 634814 592650 674258
rect 592030 634578 592062 634814
rect 592298 634578 592382 634814
rect 592618 634578 592650 634814
rect 592030 634494 592650 634578
rect 592030 634258 592062 634494
rect 592298 634258 592382 634494
rect 592618 634258 592650 634494
rect 592030 594814 592650 634258
rect 592030 594578 592062 594814
rect 592298 594578 592382 594814
rect 592618 594578 592650 594814
rect 592030 594494 592650 594578
rect 592030 594258 592062 594494
rect 592298 594258 592382 594494
rect 592618 594258 592650 594494
rect 592030 554814 592650 594258
rect 592030 554578 592062 554814
rect 592298 554578 592382 554814
rect 592618 554578 592650 554814
rect 592030 554494 592650 554578
rect 592030 554258 592062 554494
rect 592298 554258 592382 554494
rect 592618 554258 592650 554494
rect 592030 514814 592650 554258
rect 592030 514578 592062 514814
rect 592298 514578 592382 514814
rect 592618 514578 592650 514814
rect 592030 514494 592650 514578
rect 592030 514258 592062 514494
rect 592298 514258 592382 514494
rect 592618 514258 592650 514494
rect 592030 474814 592650 514258
rect 592030 474578 592062 474814
rect 592298 474578 592382 474814
rect 592618 474578 592650 474814
rect 592030 474494 592650 474578
rect 592030 474258 592062 474494
rect 592298 474258 592382 474494
rect 592618 474258 592650 474494
rect 592030 434814 592650 474258
rect 592030 434578 592062 434814
rect 592298 434578 592382 434814
rect 592618 434578 592650 434814
rect 592030 434494 592650 434578
rect 592030 434258 592062 434494
rect 592298 434258 592382 434494
rect 592618 434258 592650 434494
rect 592030 394814 592650 434258
rect 592030 394578 592062 394814
rect 592298 394578 592382 394814
rect 592618 394578 592650 394814
rect 592030 394494 592650 394578
rect 592030 394258 592062 394494
rect 592298 394258 592382 394494
rect 592618 394258 592650 394494
rect 592030 354814 592650 394258
rect 592030 354578 592062 354814
rect 592298 354578 592382 354814
rect 592618 354578 592650 354814
rect 592030 354494 592650 354578
rect 592030 354258 592062 354494
rect 592298 354258 592382 354494
rect 592618 354258 592650 354494
rect 592030 314814 592650 354258
rect 592030 314578 592062 314814
rect 592298 314578 592382 314814
rect 592618 314578 592650 314814
rect 592030 314494 592650 314578
rect 592030 314258 592062 314494
rect 592298 314258 592382 314494
rect 592618 314258 592650 314494
rect 592030 274814 592650 314258
rect 592030 274578 592062 274814
rect 592298 274578 592382 274814
rect 592618 274578 592650 274814
rect 592030 274494 592650 274578
rect 592030 274258 592062 274494
rect 592298 274258 592382 274494
rect 592618 274258 592650 274494
rect 592030 234814 592650 274258
rect 592030 234578 592062 234814
rect 592298 234578 592382 234814
rect 592618 234578 592650 234814
rect 592030 234494 592650 234578
rect 592030 234258 592062 234494
rect 592298 234258 592382 234494
rect 592618 234258 592650 234494
rect 592030 194814 592650 234258
rect 592030 194578 592062 194814
rect 592298 194578 592382 194814
rect 592618 194578 592650 194814
rect 592030 194494 592650 194578
rect 592030 194258 592062 194494
rect 592298 194258 592382 194494
rect 592618 194258 592650 194494
rect 592030 154814 592650 194258
rect 592030 154578 592062 154814
rect 592298 154578 592382 154814
rect 592618 154578 592650 154814
rect 592030 154494 592650 154578
rect 592030 154258 592062 154494
rect 592298 154258 592382 154494
rect 592618 154258 592650 154494
rect 592030 114814 592650 154258
rect 592030 114578 592062 114814
rect 592298 114578 592382 114814
rect 592618 114578 592650 114814
rect 592030 114494 592650 114578
rect 592030 114258 592062 114494
rect 592298 114258 592382 114494
rect 592618 114258 592650 114494
rect 592030 74814 592650 114258
rect 592030 74578 592062 74814
rect 592298 74578 592382 74814
rect 592618 74578 592650 74814
rect 592030 74494 592650 74578
rect 592030 74258 592062 74494
rect 592298 74258 592382 74494
rect 592618 74258 592650 74494
rect 592030 34814 592650 74258
rect 592030 34578 592062 34814
rect 592298 34578 592382 34814
rect 592618 34578 592650 34814
rect 592030 34494 592650 34578
rect 592030 34258 592062 34494
rect 592298 34258 592382 34494
rect 592618 34258 592650 34494
rect 592030 -7066 592650 34258
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 674578 -8458 674814
rect -8374 674578 -8138 674814
rect -8694 674258 -8458 674494
rect -8374 674258 -8138 674494
rect -8694 634578 -8458 634814
rect -8374 634578 -8138 634814
rect -8694 634258 -8458 634494
rect -8374 634258 -8138 634494
rect -8694 594578 -8458 594814
rect -8374 594578 -8138 594814
rect -8694 594258 -8458 594494
rect -8374 594258 -8138 594494
rect -8694 554578 -8458 554814
rect -8374 554578 -8138 554814
rect -8694 554258 -8458 554494
rect -8374 554258 -8138 554494
rect -8694 514578 -8458 514814
rect -8374 514578 -8138 514814
rect -8694 514258 -8458 514494
rect -8374 514258 -8138 514494
rect -8694 474578 -8458 474814
rect -8374 474578 -8138 474814
rect -8694 474258 -8458 474494
rect -8374 474258 -8138 474494
rect -8694 434578 -8458 434814
rect -8374 434578 -8138 434814
rect -8694 434258 -8458 434494
rect -8374 434258 -8138 434494
rect -8694 394578 -8458 394814
rect -8374 394578 -8138 394814
rect -8694 394258 -8458 394494
rect -8374 394258 -8138 394494
rect -8694 354578 -8458 354814
rect -8374 354578 -8138 354814
rect -8694 354258 -8458 354494
rect -8374 354258 -8138 354494
rect -8694 314578 -8458 314814
rect -8374 314578 -8138 314814
rect -8694 314258 -8458 314494
rect -8374 314258 -8138 314494
rect -8694 274578 -8458 274814
rect -8374 274578 -8138 274814
rect -8694 274258 -8458 274494
rect -8374 274258 -8138 274494
rect -8694 234578 -8458 234814
rect -8374 234578 -8138 234814
rect -8694 234258 -8458 234494
rect -8374 234258 -8138 234494
rect -8694 194578 -8458 194814
rect -8374 194578 -8138 194814
rect -8694 194258 -8458 194494
rect -8374 194258 -8138 194494
rect -8694 154578 -8458 154814
rect -8374 154578 -8138 154814
rect -8694 154258 -8458 154494
rect -8374 154258 -8138 154494
rect -8694 114578 -8458 114814
rect -8374 114578 -8138 114814
rect -8694 114258 -8458 114494
rect -8374 114258 -8138 114494
rect -8694 74578 -8458 74814
rect -8374 74578 -8138 74814
rect -8694 74258 -8458 74494
rect -8374 74258 -8138 74494
rect -8694 34578 -8458 34814
rect -8374 34578 -8138 34814
rect -8694 34258 -8458 34494
rect -8374 34258 -8138 34494
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 13186 710362 13422 710598
rect 13506 710362 13742 710598
rect 13186 710042 13422 710278
rect 13506 710042 13742 710278
rect -7734 694578 -7498 694814
rect -7414 694578 -7178 694814
rect -7734 694258 -7498 694494
rect -7414 694258 -7178 694494
rect -7734 654578 -7498 654814
rect -7414 654578 -7178 654814
rect -7734 654258 -7498 654494
rect -7414 654258 -7178 654494
rect -7734 614578 -7498 614814
rect -7414 614578 -7178 614814
rect -7734 614258 -7498 614494
rect -7414 614258 -7178 614494
rect -7734 574578 -7498 574814
rect -7414 574578 -7178 574814
rect -7734 574258 -7498 574494
rect -7414 574258 -7178 574494
rect -7734 534578 -7498 534814
rect -7414 534578 -7178 534814
rect -7734 534258 -7498 534494
rect -7414 534258 -7178 534494
rect -7734 494578 -7498 494814
rect -7414 494578 -7178 494814
rect -7734 494258 -7498 494494
rect -7414 494258 -7178 494494
rect -7734 454578 -7498 454814
rect -7414 454578 -7178 454814
rect -7734 454258 -7498 454494
rect -7414 454258 -7178 454494
rect -7734 414578 -7498 414814
rect -7414 414578 -7178 414814
rect -7734 414258 -7498 414494
rect -7414 414258 -7178 414494
rect -7734 374578 -7498 374814
rect -7414 374578 -7178 374814
rect -7734 374258 -7498 374494
rect -7414 374258 -7178 374494
rect -7734 334578 -7498 334814
rect -7414 334578 -7178 334814
rect -7734 334258 -7498 334494
rect -7414 334258 -7178 334494
rect -7734 294578 -7498 294814
rect -7414 294578 -7178 294814
rect -7734 294258 -7498 294494
rect -7414 294258 -7178 294494
rect -7734 254578 -7498 254814
rect -7414 254578 -7178 254814
rect -7734 254258 -7498 254494
rect -7414 254258 -7178 254494
rect -7734 214578 -7498 214814
rect -7414 214578 -7178 214814
rect -7734 214258 -7498 214494
rect -7414 214258 -7178 214494
rect -7734 174578 -7498 174814
rect -7414 174578 -7178 174814
rect -7734 174258 -7498 174494
rect -7414 174258 -7178 174494
rect -7734 134578 -7498 134814
rect -7414 134578 -7178 134814
rect -7734 134258 -7498 134494
rect -7414 134258 -7178 134494
rect -7734 94578 -7498 94814
rect -7414 94578 -7178 94814
rect -7734 94258 -7498 94494
rect -7414 94258 -7178 94494
rect -7734 54578 -7498 54814
rect -7414 54578 -7178 54814
rect -7734 54258 -7498 54494
rect -7414 54258 -7178 54494
rect -7734 14578 -7498 14814
rect -7414 14578 -7178 14814
rect -7734 14258 -7498 14494
rect -7414 14258 -7178 14494
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 670858 -6538 671094
rect -6454 670858 -6218 671094
rect -6774 670538 -6538 670774
rect -6454 670538 -6218 670774
rect -6774 630858 -6538 631094
rect -6454 630858 -6218 631094
rect -6774 630538 -6538 630774
rect -6454 630538 -6218 630774
rect -6774 590858 -6538 591094
rect -6454 590858 -6218 591094
rect -6774 590538 -6538 590774
rect -6454 590538 -6218 590774
rect -6774 550858 -6538 551094
rect -6454 550858 -6218 551094
rect -6774 550538 -6538 550774
rect -6454 550538 -6218 550774
rect -6774 510858 -6538 511094
rect -6454 510858 -6218 511094
rect -6774 510538 -6538 510774
rect -6454 510538 -6218 510774
rect -6774 470858 -6538 471094
rect -6454 470858 -6218 471094
rect -6774 470538 -6538 470774
rect -6454 470538 -6218 470774
rect -6774 430858 -6538 431094
rect -6454 430858 -6218 431094
rect -6774 430538 -6538 430774
rect -6454 430538 -6218 430774
rect -6774 390858 -6538 391094
rect -6454 390858 -6218 391094
rect -6774 390538 -6538 390774
rect -6454 390538 -6218 390774
rect -6774 350858 -6538 351094
rect -6454 350858 -6218 351094
rect -6774 350538 -6538 350774
rect -6454 350538 -6218 350774
rect -6774 310858 -6538 311094
rect -6454 310858 -6218 311094
rect -6774 310538 -6538 310774
rect -6454 310538 -6218 310774
rect -6774 270858 -6538 271094
rect -6454 270858 -6218 271094
rect -6774 270538 -6538 270774
rect -6454 270538 -6218 270774
rect -6774 230858 -6538 231094
rect -6454 230858 -6218 231094
rect -6774 230538 -6538 230774
rect -6454 230538 -6218 230774
rect -6774 190858 -6538 191094
rect -6454 190858 -6218 191094
rect -6774 190538 -6538 190774
rect -6454 190538 -6218 190774
rect -6774 150858 -6538 151094
rect -6454 150858 -6218 151094
rect -6774 150538 -6538 150774
rect -6454 150538 -6218 150774
rect -6774 110858 -6538 111094
rect -6454 110858 -6218 111094
rect -6774 110538 -6538 110774
rect -6454 110538 -6218 110774
rect -6774 70858 -6538 71094
rect -6454 70858 -6218 71094
rect -6774 70538 -6538 70774
rect -6454 70538 -6218 70774
rect -6774 30858 -6538 31094
rect -6454 30858 -6218 31094
rect -6774 30538 -6538 30774
rect -6454 30538 -6218 30774
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9466 708442 9702 708678
rect 9786 708442 10022 708678
rect 9466 708122 9702 708358
rect 9786 708122 10022 708358
rect -5814 690858 -5578 691094
rect -5494 690858 -5258 691094
rect -5814 690538 -5578 690774
rect -5494 690538 -5258 690774
rect -5814 650858 -5578 651094
rect -5494 650858 -5258 651094
rect -5814 650538 -5578 650774
rect -5494 650538 -5258 650774
rect -5814 610858 -5578 611094
rect -5494 610858 -5258 611094
rect -5814 610538 -5578 610774
rect -5494 610538 -5258 610774
rect -5814 570858 -5578 571094
rect -5494 570858 -5258 571094
rect -5814 570538 -5578 570774
rect -5494 570538 -5258 570774
rect -5814 530858 -5578 531094
rect -5494 530858 -5258 531094
rect -5814 530538 -5578 530774
rect -5494 530538 -5258 530774
rect -5814 490858 -5578 491094
rect -5494 490858 -5258 491094
rect -5814 490538 -5578 490774
rect -5494 490538 -5258 490774
rect -5814 450858 -5578 451094
rect -5494 450858 -5258 451094
rect -5814 450538 -5578 450774
rect -5494 450538 -5258 450774
rect -5814 410858 -5578 411094
rect -5494 410858 -5258 411094
rect -5814 410538 -5578 410774
rect -5494 410538 -5258 410774
rect -5814 370858 -5578 371094
rect -5494 370858 -5258 371094
rect -5814 370538 -5578 370774
rect -5494 370538 -5258 370774
rect -5814 330858 -5578 331094
rect -5494 330858 -5258 331094
rect -5814 330538 -5578 330774
rect -5494 330538 -5258 330774
rect -5814 290858 -5578 291094
rect -5494 290858 -5258 291094
rect -5814 290538 -5578 290774
rect -5494 290538 -5258 290774
rect -5814 250858 -5578 251094
rect -5494 250858 -5258 251094
rect -5814 250538 -5578 250774
rect -5494 250538 -5258 250774
rect -5814 210858 -5578 211094
rect -5494 210858 -5258 211094
rect -5814 210538 -5578 210774
rect -5494 210538 -5258 210774
rect -5814 170858 -5578 171094
rect -5494 170858 -5258 171094
rect -5814 170538 -5578 170774
rect -5494 170538 -5258 170774
rect -5814 130858 -5578 131094
rect -5494 130858 -5258 131094
rect -5814 130538 -5578 130774
rect -5494 130538 -5258 130774
rect -5814 90858 -5578 91094
rect -5494 90858 -5258 91094
rect -5814 90538 -5578 90774
rect -5494 90538 -5258 90774
rect -5814 50858 -5578 51094
rect -5494 50858 -5258 51094
rect -5814 50538 -5578 50774
rect -5494 50538 -5258 50774
rect -5814 10858 -5578 11094
rect -5494 10858 -5258 11094
rect -5814 10538 -5578 10774
rect -5494 10538 -5258 10774
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 667138 -4618 667374
rect -4534 667138 -4298 667374
rect -4854 666818 -4618 667054
rect -4534 666818 -4298 667054
rect -4854 627138 -4618 627374
rect -4534 627138 -4298 627374
rect -4854 626818 -4618 627054
rect -4534 626818 -4298 627054
rect -4854 587138 -4618 587374
rect -4534 587138 -4298 587374
rect -4854 586818 -4618 587054
rect -4534 586818 -4298 587054
rect -4854 547138 -4618 547374
rect -4534 547138 -4298 547374
rect -4854 546818 -4618 547054
rect -4534 546818 -4298 547054
rect -4854 507138 -4618 507374
rect -4534 507138 -4298 507374
rect -4854 506818 -4618 507054
rect -4534 506818 -4298 507054
rect -4854 467138 -4618 467374
rect -4534 467138 -4298 467374
rect -4854 466818 -4618 467054
rect -4534 466818 -4298 467054
rect -4854 427138 -4618 427374
rect -4534 427138 -4298 427374
rect -4854 426818 -4618 427054
rect -4534 426818 -4298 427054
rect -4854 387138 -4618 387374
rect -4534 387138 -4298 387374
rect -4854 386818 -4618 387054
rect -4534 386818 -4298 387054
rect -4854 347138 -4618 347374
rect -4534 347138 -4298 347374
rect -4854 346818 -4618 347054
rect -4534 346818 -4298 347054
rect -4854 307138 -4618 307374
rect -4534 307138 -4298 307374
rect -4854 306818 -4618 307054
rect -4534 306818 -4298 307054
rect -4854 267138 -4618 267374
rect -4534 267138 -4298 267374
rect -4854 266818 -4618 267054
rect -4534 266818 -4298 267054
rect -4854 227138 -4618 227374
rect -4534 227138 -4298 227374
rect -4854 226818 -4618 227054
rect -4534 226818 -4298 227054
rect -4854 187138 -4618 187374
rect -4534 187138 -4298 187374
rect -4854 186818 -4618 187054
rect -4534 186818 -4298 187054
rect -4854 147138 -4618 147374
rect -4534 147138 -4298 147374
rect -4854 146818 -4618 147054
rect -4534 146818 -4298 147054
rect -4854 107138 -4618 107374
rect -4534 107138 -4298 107374
rect -4854 106818 -4618 107054
rect -4534 106818 -4298 107054
rect -4854 67138 -4618 67374
rect -4534 67138 -4298 67374
rect -4854 66818 -4618 67054
rect -4534 66818 -4298 67054
rect -4854 27138 -4618 27374
rect -4534 27138 -4298 27374
rect -4854 26818 -4618 27054
rect -4534 26818 -4298 27054
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5746 706522 5982 706758
rect 6066 706522 6302 706758
rect 5746 706202 5982 706438
rect 6066 706202 6302 706438
rect -3894 687138 -3658 687374
rect -3574 687138 -3338 687374
rect -3894 686818 -3658 687054
rect -3574 686818 -3338 687054
rect -3894 647138 -3658 647374
rect -3574 647138 -3338 647374
rect -3894 646818 -3658 647054
rect -3574 646818 -3338 647054
rect -3894 607138 -3658 607374
rect -3574 607138 -3338 607374
rect -3894 606818 -3658 607054
rect -3574 606818 -3338 607054
rect -3894 567138 -3658 567374
rect -3574 567138 -3338 567374
rect -3894 566818 -3658 567054
rect -3574 566818 -3338 567054
rect -3894 527138 -3658 527374
rect -3574 527138 -3338 527374
rect -3894 526818 -3658 527054
rect -3574 526818 -3338 527054
rect -3894 487138 -3658 487374
rect -3574 487138 -3338 487374
rect -3894 486818 -3658 487054
rect -3574 486818 -3338 487054
rect -3894 447138 -3658 447374
rect -3574 447138 -3338 447374
rect -3894 446818 -3658 447054
rect -3574 446818 -3338 447054
rect -3894 407138 -3658 407374
rect -3574 407138 -3338 407374
rect -3894 406818 -3658 407054
rect -3574 406818 -3338 407054
rect -3894 367138 -3658 367374
rect -3574 367138 -3338 367374
rect -3894 366818 -3658 367054
rect -3574 366818 -3338 367054
rect -3894 327138 -3658 327374
rect -3574 327138 -3338 327374
rect -3894 326818 -3658 327054
rect -3574 326818 -3338 327054
rect -3894 287138 -3658 287374
rect -3574 287138 -3338 287374
rect -3894 286818 -3658 287054
rect -3574 286818 -3338 287054
rect -3894 247138 -3658 247374
rect -3574 247138 -3338 247374
rect -3894 246818 -3658 247054
rect -3574 246818 -3338 247054
rect -3894 207138 -3658 207374
rect -3574 207138 -3338 207374
rect -3894 206818 -3658 207054
rect -3574 206818 -3338 207054
rect -3894 167138 -3658 167374
rect -3574 167138 -3338 167374
rect -3894 166818 -3658 167054
rect -3574 166818 -3338 167054
rect -3894 127138 -3658 127374
rect -3574 127138 -3338 127374
rect -3894 126818 -3658 127054
rect -3574 126818 -3338 127054
rect -3894 87138 -3658 87374
rect -3574 87138 -3338 87374
rect -3894 86818 -3658 87054
rect -3574 86818 -3338 87054
rect -3894 47138 -3658 47374
rect -3574 47138 -3338 47374
rect -3894 46818 -3658 47054
rect -3574 46818 -3338 47054
rect -3894 7138 -3658 7374
rect -3574 7138 -3338 7374
rect -3894 6818 -3658 7054
rect -3574 6818 -3338 7054
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 663418 -2698 663654
rect -2614 663418 -2378 663654
rect -2934 663098 -2698 663334
rect -2614 663098 -2378 663334
rect -2934 623418 -2698 623654
rect -2614 623418 -2378 623654
rect -2934 623098 -2698 623334
rect -2614 623098 -2378 623334
rect -2934 583418 -2698 583654
rect -2614 583418 -2378 583654
rect -2934 583098 -2698 583334
rect -2614 583098 -2378 583334
rect -2934 543418 -2698 543654
rect -2614 543418 -2378 543654
rect -2934 543098 -2698 543334
rect -2614 543098 -2378 543334
rect -2934 503418 -2698 503654
rect -2614 503418 -2378 503654
rect -2934 503098 -2698 503334
rect -2614 503098 -2378 503334
rect -2934 463418 -2698 463654
rect -2614 463418 -2378 463654
rect -2934 463098 -2698 463334
rect -2614 463098 -2378 463334
rect -2934 423418 -2698 423654
rect -2614 423418 -2378 423654
rect -2934 423098 -2698 423334
rect -2614 423098 -2378 423334
rect -2934 383418 -2698 383654
rect -2614 383418 -2378 383654
rect -2934 383098 -2698 383334
rect -2614 383098 -2378 383334
rect -2934 343418 -2698 343654
rect -2614 343418 -2378 343654
rect -2934 343098 -2698 343334
rect -2614 343098 -2378 343334
rect -2934 303418 -2698 303654
rect -2614 303418 -2378 303654
rect -2934 303098 -2698 303334
rect -2614 303098 -2378 303334
rect -2934 263418 -2698 263654
rect -2614 263418 -2378 263654
rect -2934 263098 -2698 263334
rect -2614 263098 -2378 263334
rect -2934 223418 -2698 223654
rect -2614 223418 -2378 223654
rect -2934 223098 -2698 223334
rect -2614 223098 -2378 223334
rect -2934 183418 -2698 183654
rect -2614 183418 -2378 183654
rect -2934 183098 -2698 183334
rect -2614 183098 -2378 183334
rect -2934 143418 -2698 143654
rect -2614 143418 -2378 143654
rect -2934 143098 -2698 143334
rect -2614 143098 -2378 143334
rect -2934 103418 -2698 103654
rect -2614 103418 -2378 103654
rect -2934 103098 -2698 103334
rect -2614 103098 -2378 103334
rect -2934 63418 -2698 63654
rect -2614 63418 -2378 63654
rect -2934 63098 -2698 63334
rect -2614 63098 -2378 63334
rect -2934 23418 -2698 23654
rect -2614 23418 -2378 23654
rect -2934 23098 -2698 23334
rect -2614 23098 -2378 23334
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect 2026 704602 2262 704838
rect 2346 704602 2582 704838
rect 2026 704282 2262 704518
rect 2346 704282 2582 704518
rect 33186 711322 33422 711558
rect 33506 711322 33742 711558
rect 33186 711002 33422 711238
rect 33506 711002 33742 711238
rect 29466 709402 29702 709638
rect 29786 709402 30022 709638
rect 29466 709082 29702 709318
rect 29786 709082 30022 709318
rect 25746 707482 25982 707718
rect 26066 707482 26302 707718
rect 25746 707162 25982 707398
rect 26066 707162 26302 707398
rect 22026 705562 22262 705798
rect 22346 705562 22582 705798
rect 22026 705242 22262 705478
rect 22346 705242 22582 705478
rect 53186 710362 53422 710598
rect 53506 710362 53742 710598
rect 53186 710042 53422 710278
rect 53506 710042 53742 710278
rect 49466 708442 49702 708678
rect 49786 708442 50022 708678
rect 49466 708122 49702 708358
rect 49786 708122 50022 708358
rect 45746 706522 45982 706758
rect 46066 706522 46302 706758
rect 45746 706202 45982 706438
rect 46066 706202 46302 706438
rect 42026 704602 42262 704838
rect 42346 704602 42582 704838
rect 42026 704282 42262 704518
rect 42346 704282 42582 704518
rect 73186 711322 73422 711558
rect 73506 711322 73742 711558
rect 73186 711002 73422 711238
rect 73506 711002 73742 711238
rect 69466 709402 69702 709638
rect 69786 709402 70022 709638
rect 69466 709082 69702 709318
rect 69786 709082 70022 709318
rect 65746 707482 65982 707718
rect 66066 707482 66302 707718
rect 65746 707162 65982 707398
rect 66066 707162 66302 707398
rect 62026 705562 62262 705798
rect 62346 705562 62582 705798
rect 62026 705242 62262 705478
rect 62346 705242 62582 705478
rect 93186 710362 93422 710598
rect 93506 710362 93742 710598
rect 93186 710042 93422 710278
rect 93506 710042 93742 710278
rect 89466 708442 89702 708678
rect 89786 708442 90022 708678
rect 89466 708122 89702 708358
rect 89786 708122 90022 708358
rect 85746 706522 85982 706758
rect 86066 706522 86302 706758
rect 85746 706202 85982 706438
rect 86066 706202 86302 706438
rect 82026 704602 82262 704838
rect 82346 704602 82582 704838
rect 82026 704282 82262 704518
rect 82346 704282 82582 704518
rect 113186 711322 113422 711558
rect 113506 711322 113742 711558
rect 113186 711002 113422 711238
rect 113506 711002 113742 711238
rect 109466 709402 109702 709638
rect 109786 709402 110022 709638
rect 109466 709082 109702 709318
rect 109786 709082 110022 709318
rect 105746 707482 105982 707718
rect 106066 707482 106302 707718
rect 105746 707162 105982 707398
rect 106066 707162 106302 707398
rect 102026 705562 102262 705798
rect 102346 705562 102582 705798
rect 102026 705242 102262 705478
rect 102346 705242 102582 705478
rect 133186 710362 133422 710598
rect 133506 710362 133742 710598
rect 133186 710042 133422 710278
rect 133506 710042 133742 710278
rect 129466 708442 129702 708678
rect 129786 708442 130022 708678
rect 129466 708122 129702 708358
rect 129786 708122 130022 708358
rect 125746 706522 125982 706758
rect 126066 706522 126302 706758
rect 125746 706202 125982 706438
rect 126066 706202 126302 706438
rect 122026 704602 122262 704838
rect 122346 704602 122582 704838
rect 122026 704282 122262 704518
rect 122346 704282 122582 704518
rect 153186 711322 153422 711558
rect 153506 711322 153742 711558
rect 153186 711002 153422 711238
rect 153506 711002 153742 711238
rect 149466 709402 149702 709638
rect 149786 709402 150022 709638
rect 149466 709082 149702 709318
rect 149786 709082 150022 709318
rect 145746 707482 145982 707718
rect 146066 707482 146302 707718
rect 145746 707162 145982 707398
rect 146066 707162 146302 707398
rect 142026 705562 142262 705798
rect 142346 705562 142582 705798
rect 142026 705242 142262 705478
rect 142346 705242 142582 705478
rect 173186 710362 173422 710598
rect 173506 710362 173742 710598
rect 173186 710042 173422 710278
rect 173506 710042 173742 710278
rect 169466 708442 169702 708678
rect 169786 708442 170022 708678
rect 169466 708122 169702 708358
rect 169786 708122 170022 708358
rect 165746 706522 165982 706758
rect 166066 706522 166302 706758
rect 165746 706202 165982 706438
rect 166066 706202 166302 706438
rect 162026 704602 162262 704838
rect 162346 704602 162582 704838
rect 162026 704282 162262 704518
rect 162346 704282 162582 704518
rect 193186 711322 193422 711558
rect 193506 711322 193742 711558
rect 193186 711002 193422 711238
rect 193506 711002 193742 711238
rect 189466 709402 189702 709638
rect 189786 709402 190022 709638
rect 189466 709082 189702 709318
rect 189786 709082 190022 709318
rect 185746 707482 185982 707718
rect 186066 707482 186302 707718
rect 185746 707162 185982 707398
rect 186066 707162 186302 707398
rect 182026 705562 182262 705798
rect 182346 705562 182582 705798
rect 182026 705242 182262 705478
rect 182346 705242 182582 705478
rect 213186 710362 213422 710598
rect 213506 710362 213742 710598
rect 213186 710042 213422 710278
rect 213506 710042 213742 710278
rect 209466 708442 209702 708678
rect 209786 708442 210022 708678
rect 209466 708122 209702 708358
rect 209786 708122 210022 708358
rect 205746 706522 205982 706758
rect 206066 706522 206302 706758
rect 205746 706202 205982 706438
rect 206066 706202 206302 706438
rect 202026 704602 202262 704838
rect 202346 704602 202582 704838
rect 202026 704282 202262 704518
rect 202346 704282 202582 704518
rect 233186 711322 233422 711558
rect 233506 711322 233742 711558
rect 233186 711002 233422 711238
rect 233506 711002 233742 711238
rect 229466 709402 229702 709638
rect 229786 709402 230022 709638
rect 229466 709082 229702 709318
rect 229786 709082 230022 709318
rect 225746 707482 225982 707718
rect 226066 707482 226302 707718
rect 225746 707162 225982 707398
rect 226066 707162 226302 707398
rect 222026 705562 222262 705798
rect 222346 705562 222582 705798
rect 222026 705242 222262 705478
rect 222346 705242 222582 705478
rect 253186 710362 253422 710598
rect 253506 710362 253742 710598
rect 253186 710042 253422 710278
rect 253506 710042 253742 710278
rect 249466 708442 249702 708678
rect 249786 708442 250022 708678
rect 249466 708122 249702 708358
rect 249786 708122 250022 708358
rect 245746 706522 245982 706758
rect 246066 706522 246302 706758
rect 245746 706202 245982 706438
rect 246066 706202 246302 706438
rect 242026 704602 242262 704838
rect 242346 704602 242582 704838
rect 242026 704282 242262 704518
rect 242346 704282 242582 704518
rect 273186 711322 273422 711558
rect 273506 711322 273742 711558
rect 273186 711002 273422 711238
rect 273506 711002 273742 711238
rect 269466 709402 269702 709638
rect 269786 709402 270022 709638
rect 269466 709082 269702 709318
rect 269786 709082 270022 709318
rect 265746 707482 265982 707718
rect 266066 707482 266302 707718
rect 265746 707162 265982 707398
rect 266066 707162 266302 707398
rect 262026 705562 262262 705798
rect 262346 705562 262582 705798
rect 262026 705242 262262 705478
rect 262346 705242 262582 705478
rect 293186 710362 293422 710598
rect 293506 710362 293742 710598
rect 293186 710042 293422 710278
rect 293506 710042 293742 710278
rect 289466 708442 289702 708678
rect 289786 708442 290022 708678
rect 289466 708122 289702 708358
rect 289786 708122 290022 708358
rect 285746 706522 285982 706758
rect 286066 706522 286302 706758
rect 285746 706202 285982 706438
rect 286066 706202 286302 706438
rect 282026 704602 282262 704838
rect 282346 704602 282582 704838
rect 282026 704282 282262 704518
rect 282346 704282 282582 704518
rect 313186 711322 313422 711558
rect 313506 711322 313742 711558
rect 313186 711002 313422 711238
rect 313506 711002 313742 711238
rect 309466 709402 309702 709638
rect 309786 709402 310022 709638
rect 309466 709082 309702 709318
rect 309786 709082 310022 709318
rect 305746 707482 305982 707718
rect 306066 707482 306302 707718
rect 305746 707162 305982 707398
rect 306066 707162 306302 707398
rect 302026 705562 302262 705798
rect 302346 705562 302582 705798
rect 302026 705242 302262 705478
rect 302346 705242 302582 705478
rect 333186 710362 333422 710598
rect 333506 710362 333742 710598
rect 333186 710042 333422 710278
rect 333506 710042 333742 710278
rect 329466 708442 329702 708678
rect 329786 708442 330022 708678
rect 329466 708122 329702 708358
rect 329786 708122 330022 708358
rect 325746 706522 325982 706758
rect 326066 706522 326302 706758
rect 325746 706202 325982 706438
rect 326066 706202 326302 706438
rect 322026 704602 322262 704838
rect 322346 704602 322582 704838
rect 322026 704282 322262 704518
rect 322346 704282 322582 704518
rect 353186 711322 353422 711558
rect 353506 711322 353742 711558
rect 353186 711002 353422 711238
rect 353506 711002 353742 711238
rect 349466 709402 349702 709638
rect 349786 709402 350022 709638
rect 349466 709082 349702 709318
rect 349786 709082 350022 709318
rect 345746 707482 345982 707718
rect 346066 707482 346302 707718
rect 345746 707162 345982 707398
rect 346066 707162 346302 707398
rect 342026 705562 342262 705798
rect 342346 705562 342582 705798
rect 342026 705242 342262 705478
rect 342346 705242 342582 705478
rect 373186 710362 373422 710598
rect 373506 710362 373742 710598
rect 373186 710042 373422 710278
rect 373506 710042 373742 710278
rect 369466 708442 369702 708678
rect 369786 708442 370022 708678
rect 369466 708122 369702 708358
rect 369786 708122 370022 708358
rect 365746 706522 365982 706758
rect 366066 706522 366302 706758
rect 365746 706202 365982 706438
rect 366066 706202 366302 706438
rect 362026 704602 362262 704838
rect 362346 704602 362582 704838
rect 362026 704282 362262 704518
rect 362346 704282 362582 704518
rect 393186 711322 393422 711558
rect 393506 711322 393742 711558
rect 393186 711002 393422 711238
rect 393506 711002 393742 711238
rect 389466 709402 389702 709638
rect 389786 709402 390022 709638
rect 389466 709082 389702 709318
rect 389786 709082 390022 709318
rect 385746 707482 385982 707718
rect 386066 707482 386302 707718
rect 385746 707162 385982 707398
rect 386066 707162 386302 707398
rect 382026 705562 382262 705798
rect 382346 705562 382582 705798
rect 382026 705242 382262 705478
rect 382346 705242 382582 705478
rect 413186 710362 413422 710598
rect 413506 710362 413742 710598
rect 413186 710042 413422 710278
rect 413506 710042 413742 710278
rect 409466 708442 409702 708678
rect 409786 708442 410022 708678
rect 409466 708122 409702 708358
rect 409786 708122 410022 708358
rect 405746 706522 405982 706758
rect 406066 706522 406302 706758
rect 405746 706202 405982 706438
rect 406066 706202 406302 706438
rect 402026 704602 402262 704838
rect 402346 704602 402582 704838
rect 402026 704282 402262 704518
rect 402346 704282 402582 704518
rect 433186 711322 433422 711558
rect 433506 711322 433742 711558
rect 433186 711002 433422 711238
rect 433506 711002 433742 711238
rect 429466 709402 429702 709638
rect 429786 709402 430022 709638
rect 429466 709082 429702 709318
rect 429786 709082 430022 709318
rect 425746 707482 425982 707718
rect 426066 707482 426302 707718
rect 425746 707162 425982 707398
rect 426066 707162 426302 707398
rect 422026 705562 422262 705798
rect 422346 705562 422582 705798
rect 422026 705242 422262 705478
rect 422346 705242 422582 705478
rect 453186 710362 453422 710598
rect 453506 710362 453742 710598
rect 453186 710042 453422 710278
rect 453506 710042 453742 710278
rect 449466 708442 449702 708678
rect 449786 708442 450022 708678
rect 449466 708122 449702 708358
rect 449786 708122 450022 708358
rect 445746 706522 445982 706758
rect 446066 706522 446302 706758
rect 445746 706202 445982 706438
rect 446066 706202 446302 706438
rect 442026 704602 442262 704838
rect 442346 704602 442582 704838
rect 442026 704282 442262 704518
rect 442346 704282 442582 704518
rect 473186 711322 473422 711558
rect 473506 711322 473742 711558
rect 473186 711002 473422 711238
rect 473506 711002 473742 711238
rect 469466 709402 469702 709638
rect 469786 709402 470022 709638
rect 469466 709082 469702 709318
rect 469786 709082 470022 709318
rect 465746 707482 465982 707718
rect 466066 707482 466302 707718
rect 465746 707162 465982 707398
rect 466066 707162 466302 707398
rect 462026 705562 462262 705798
rect 462346 705562 462582 705798
rect 462026 705242 462262 705478
rect 462346 705242 462582 705478
rect 493186 710362 493422 710598
rect 493506 710362 493742 710598
rect 493186 710042 493422 710278
rect 493506 710042 493742 710278
rect 489466 708442 489702 708678
rect 489786 708442 490022 708678
rect 489466 708122 489702 708358
rect 489786 708122 490022 708358
rect 485746 706522 485982 706758
rect 486066 706522 486302 706758
rect 485746 706202 485982 706438
rect 486066 706202 486302 706438
rect 482026 704602 482262 704838
rect 482346 704602 482582 704838
rect 482026 704282 482262 704518
rect 482346 704282 482582 704518
rect 513186 711322 513422 711558
rect 513506 711322 513742 711558
rect 513186 711002 513422 711238
rect 513506 711002 513742 711238
rect 509466 709402 509702 709638
rect 509786 709402 510022 709638
rect 509466 709082 509702 709318
rect 509786 709082 510022 709318
rect 505746 707482 505982 707718
rect 506066 707482 506302 707718
rect 505746 707162 505982 707398
rect 506066 707162 506302 707398
rect 502026 705562 502262 705798
rect 502346 705562 502582 705798
rect 502026 705242 502262 705478
rect 502346 705242 502582 705478
rect 533186 710362 533422 710598
rect 533506 710362 533742 710598
rect 533186 710042 533422 710278
rect 533506 710042 533742 710278
rect 529466 708442 529702 708678
rect 529786 708442 530022 708678
rect 529466 708122 529702 708358
rect 529786 708122 530022 708358
rect 525746 706522 525982 706758
rect 526066 706522 526302 706758
rect 525746 706202 525982 706438
rect 526066 706202 526302 706438
rect 522026 704602 522262 704838
rect 522346 704602 522582 704838
rect 522026 704282 522262 704518
rect 522346 704282 522582 704518
rect 553186 711322 553422 711558
rect 553506 711322 553742 711558
rect 553186 711002 553422 711238
rect 553506 711002 553742 711238
rect 549466 709402 549702 709638
rect 549786 709402 550022 709638
rect 549466 709082 549702 709318
rect 549786 709082 550022 709318
rect 545746 707482 545982 707718
rect 546066 707482 546302 707718
rect 545746 707162 545982 707398
rect 546066 707162 546302 707398
rect 542026 705562 542262 705798
rect 542346 705562 542582 705798
rect 542026 705242 542262 705478
rect 542346 705242 542582 705478
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 573186 710362 573422 710598
rect 573506 710362 573742 710598
rect 573186 710042 573422 710278
rect 573506 710042 573742 710278
rect 569466 708442 569702 708678
rect 569786 708442 570022 708678
rect 569466 708122 569702 708358
rect 569786 708122 570022 708358
rect 565746 706522 565982 706758
rect 566066 706522 566302 706758
rect 565746 706202 565982 706438
rect 566066 706202 566302 706438
rect 562026 704602 562262 704838
rect 562346 704602 562582 704838
rect 562026 704282 562262 704518
rect 562346 704282 562582 704518
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect -1974 683418 -1738 683654
rect -1654 683418 -1418 683654
rect -1974 683098 -1738 683334
rect -1654 683098 -1418 683334
rect 9116 683418 9352 683654
rect 9436 683418 9672 683654
rect 9116 683098 9352 683334
rect 9436 683098 9672 683334
rect 56652 683418 56888 683654
rect 56972 683418 57208 683654
rect 56652 683098 56888 683334
rect 56972 683098 57208 683334
rect 92652 683418 92888 683654
rect 92972 683418 93208 683654
rect 92652 683098 92888 683334
rect 92972 683098 93208 683334
rect 128652 683418 128888 683654
rect 128972 683418 129208 683654
rect 128652 683098 128888 683334
rect 128972 683098 129208 683334
rect 164652 683418 164888 683654
rect 164972 683418 165208 683654
rect 164652 683098 164888 683334
rect 164972 683098 165208 683334
rect 200652 683418 200888 683654
rect 200972 683418 201208 683654
rect 200652 683098 200888 683334
rect 200972 683098 201208 683334
rect 236652 683418 236888 683654
rect 236972 683418 237208 683654
rect 236652 683098 236888 683334
rect 236972 683098 237208 683334
rect 272652 683418 272888 683654
rect 272972 683418 273208 683654
rect 272652 683098 272888 683334
rect 272972 683098 273208 683334
rect 308652 683418 308888 683654
rect 308972 683418 309208 683654
rect 308652 683098 308888 683334
rect 308972 683098 309208 683334
rect 344652 683418 344888 683654
rect 344972 683418 345208 683654
rect 344652 683098 344888 683334
rect 344972 683098 345208 683334
rect 380652 683418 380888 683654
rect 380972 683418 381208 683654
rect 380652 683098 380888 683334
rect 380972 683098 381208 683334
rect 416652 683418 416888 683654
rect 416972 683418 417208 683654
rect 416652 683098 416888 683334
rect 416972 683098 417208 683334
rect 452652 683418 452888 683654
rect 452972 683418 453208 683654
rect 452652 683098 452888 683334
rect 452972 683098 453208 683334
rect 488652 683418 488888 683654
rect 488972 683418 489208 683654
rect 488652 683098 488888 683334
rect 488972 683098 489208 683334
rect 524652 683418 524888 683654
rect 524972 683418 525208 683654
rect 524652 683098 524888 683334
rect 524972 683098 525208 683334
rect 560652 683418 560888 683654
rect 560972 683418 561208 683654
rect 560652 683098 560888 683334
rect 560972 683098 561208 683334
rect 570292 683418 570528 683654
rect 570612 683418 570848 683654
rect 570292 683098 570528 683334
rect 570612 683098 570848 683334
rect 585342 683418 585578 683654
rect 585662 683418 585898 683654
rect 585342 683098 585578 683334
rect 585662 683098 585898 683334
rect 7876 663418 8112 663654
rect 8196 663418 8432 663654
rect 7876 663098 8112 663334
rect 8196 663098 8432 663334
rect 38032 663418 38268 663654
rect 38352 663418 38588 663654
rect 38032 663098 38268 663334
rect 38352 663098 38588 663334
rect 74032 663418 74268 663654
rect 74352 663418 74588 663654
rect 74032 663098 74268 663334
rect 74352 663098 74588 663334
rect 110032 663418 110268 663654
rect 110352 663418 110588 663654
rect 110032 663098 110268 663334
rect 110352 663098 110588 663334
rect 146032 663418 146268 663654
rect 146352 663418 146588 663654
rect 146032 663098 146268 663334
rect 146352 663098 146588 663334
rect 182032 663418 182268 663654
rect 182352 663418 182588 663654
rect 182032 663098 182268 663334
rect 182352 663098 182588 663334
rect 218032 663418 218268 663654
rect 218352 663418 218588 663654
rect 218032 663098 218268 663334
rect 218352 663098 218588 663334
rect 254032 663418 254268 663654
rect 254352 663418 254588 663654
rect 254032 663098 254268 663334
rect 254352 663098 254588 663334
rect 290032 663418 290268 663654
rect 290352 663418 290588 663654
rect 290032 663098 290268 663334
rect 290352 663098 290588 663334
rect 326032 663418 326268 663654
rect 326352 663418 326588 663654
rect 326032 663098 326268 663334
rect 326352 663098 326588 663334
rect 362032 663418 362268 663654
rect 362352 663418 362588 663654
rect 362032 663098 362268 663334
rect 362352 663098 362588 663334
rect 398032 663418 398268 663654
rect 398352 663418 398588 663654
rect 398032 663098 398268 663334
rect 398352 663098 398588 663334
rect 434032 663418 434268 663654
rect 434352 663418 434588 663654
rect 434032 663098 434268 663334
rect 434352 663098 434588 663334
rect 470032 663418 470268 663654
rect 470352 663418 470588 663654
rect 470032 663098 470268 663334
rect 470352 663098 470588 663334
rect 506032 663418 506268 663654
rect 506352 663418 506588 663654
rect 506032 663098 506268 663334
rect 506352 663098 506588 663334
rect 542032 663418 542268 663654
rect 542352 663418 542588 663654
rect 542032 663098 542268 663334
rect 542352 663098 542588 663334
rect 571532 663418 571768 663654
rect 571852 663418 572088 663654
rect 571532 663098 571768 663334
rect 571852 663098 572088 663334
rect -1974 643418 -1738 643654
rect -1654 643418 -1418 643654
rect -1974 643098 -1738 643334
rect -1654 643098 -1418 643334
rect 9116 643418 9352 643654
rect 9436 643418 9672 643654
rect 9116 643098 9352 643334
rect 9436 643098 9672 643334
rect 56652 643418 56888 643654
rect 56972 643418 57208 643654
rect 56652 643098 56888 643334
rect 56972 643098 57208 643334
rect 92652 643418 92888 643654
rect 92972 643418 93208 643654
rect 92652 643098 92888 643334
rect 92972 643098 93208 643334
rect 128652 643418 128888 643654
rect 128972 643418 129208 643654
rect 128652 643098 128888 643334
rect 128972 643098 129208 643334
rect 164652 643418 164888 643654
rect 164972 643418 165208 643654
rect 164652 643098 164888 643334
rect 164972 643098 165208 643334
rect 200652 643418 200888 643654
rect 200972 643418 201208 643654
rect 200652 643098 200888 643334
rect 200972 643098 201208 643334
rect 236652 643418 236888 643654
rect 236972 643418 237208 643654
rect 236652 643098 236888 643334
rect 236972 643098 237208 643334
rect 272652 643418 272888 643654
rect 272972 643418 273208 643654
rect 272652 643098 272888 643334
rect 272972 643098 273208 643334
rect 308652 643418 308888 643654
rect 308972 643418 309208 643654
rect 308652 643098 308888 643334
rect 308972 643098 309208 643334
rect 344652 643418 344888 643654
rect 344972 643418 345208 643654
rect 344652 643098 344888 643334
rect 344972 643098 345208 643334
rect 380652 643418 380888 643654
rect 380972 643418 381208 643654
rect 380652 643098 380888 643334
rect 380972 643098 381208 643334
rect 416652 643418 416888 643654
rect 416972 643418 417208 643654
rect 416652 643098 416888 643334
rect 416972 643098 417208 643334
rect 452652 643418 452888 643654
rect 452972 643418 453208 643654
rect 452652 643098 452888 643334
rect 452972 643098 453208 643334
rect 488652 643418 488888 643654
rect 488972 643418 489208 643654
rect 488652 643098 488888 643334
rect 488972 643098 489208 643334
rect 524652 643418 524888 643654
rect 524972 643418 525208 643654
rect 524652 643098 524888 643334
rect 524972 643098 525208 643334
rect 560652 643418 560888 643654
rect 560972 643418 561208 643654
rect 560652 643098 560888 643334
rect 560972 643098 561208 643334
rect 570292 643418 570528 643654
rect 570612 643418 570848 643654
rect 570292 643098 570528 643334
rect 570612 643098 570848 643334
rect 585342 643418 585578 643654
rect 585662 643418 585898 643654
rect 585342 643098 585578 643334
rect 585662 643098 585898 643334
rect 7876 623418 8112 623654
rect 8196 623418 8432 623654
rect 7876 623098 8112 623334
rect 8196 623098 8432 623334
rect 38032 623418 38268 623654
rect 38352 623418 38588 623654
rect 38032 623098 38268 623334
rect 38352 623098 38588 623334
rect 74032 623418 74268 623654
rect 74352 623418 74588 623654
rect 74032 623098 74268 623334
rect 74352 623098 74588 623334
rect 110032 623418 110268 623654
rect 110352 623418 110588 623654
rect 110032 623098 110268 623334
rect 110352 623098 110588 623334
rect 146032 623418 146268 623654
rect 146352 623418 146588 623654
rect 146032 623098 146268 623334
rect 146352 623098 146588 623334
rect 182032 623418 182268 623654
rect 182352 623418 182588 623654
rect 182032 623098 182268 623334
rect 182352 623098 182588 623334
rect 218032 623418 218268 623654
rect 218352 623418 218588 623654
rect 218032 623098 218268 623334
rect 218352 623098 218588 623334
rect 254032 623418 254268 623654
rect 254352 623418 254588 623654
rect 254032 623098 254268 623334
rect 254352 623098 254588 623334
rect 290032 623418 290268 623654
rect 290352 623418 290588 623654
rect 290032 623098 290268 623334
rect 290352 623098 290588 623334
rect 326032 623418 326268 623654
rect 326352 623418 326588 623654
rect 326032 623098 326268 623334
rect 326352 623098 326588 623334
rect 362032 623418 362268 623654
rect 362352 623418 362588 623654
rect 362032 623098 362268 623334
rect 362352 623098 362588 623334
rect 398032 623418 398268 623654
rect 398352 623418 398588 623654
rect 398032 623098 398268 623334
rect 398352 623098 398588 623334
rect 434032 623418 434268 623654
rect 434352 623418 434588 623654
rect 434032 623098 434268 623334
rect 434352 623098 434588 623334
rect 470032 623418 470268 623654
rect 470352 623418 470588 623654
rect 470032 623098 470268 623334
rect 470352 623098 470588 623334
rect 506032 623418 506268 623654
rect 506352 623418 506588 623654
rect 506032 623098 506268 623334
rect 506352 623098 506588 623334
rect 542032 623418 542268 623654
rect 542352 623418 542588 623654
rect 542032 623098 542268 623334
rect 542352 623098 542588 623334
rect 571532 623418 571768 623654
rect 571852 623418 572088 623654
rect 571532 623098 571768 623334
rect 571852 623098 572088 623334
rect -1974 603418 -1738 603654
rect -1654 603418 -1418 603654
rect -1974 603098 -1738 603334
rect -1654 603098 -1418 603334
rect 9116 603418 9352 603654
rect 9436 603418 9672 603654
rect 9116 603098 9352 603334
rect 9436 603098 9672 603334
rect 56652 603418 56888 603654
rect 56972 603418 57208 603654
rect 56652 603098 56888 603334
rect 56972 603098 57208 603334
rect 92652 603418 92888 603654
rect 92972 603418 93208 603654
rect 92652 603098 92888 603334
rect 92972 603098 93208 603334
rect 128652 603418 128888 603654
rect 128972 603418 129208 603654
rect 128652 603098 128888 603334
rect 128972 603098 129208 603334
rect 164652 603418 164888 603654
rect 164972 603418 165208 603654
rect 164652 603098 164888 603334
rect 164972 603098 165208 603334
rect 200652 603418 200888 603654
rect 200972 603418 201208 603654
rect 200652 603098 200888 603334
rect 200972 603098 201208 603334
rect 236652 603418 236888 603654
rect 236972 603418 237208 603654
rect 236652 603098 236888 603334
rect 236972 603098 237208 603334
rect 272652 603418 272888 603654
rect 272972 603418 273208 603654
rect 272652 603098 272888 603334
rect 272972 603098 273208 603334
rect 308652 603418 308888 603654
rect 308972 603418 309208 603654
rect 308652 603098 308888 603334
rect 308972 603098 309208 603334
rect 344652 603418 344888 603654
rect 344972 603418 345208 603654
rect 344652 603098 344888 603334
rect 344972 603098 345208 603334
rect 380652 603418 380888 603654
rect 380972 603418 381208 603654
rect 380652 603098 380888 603334
rect 380972 603098 381208 603334
rect 416652 603418 416888 603654
rect 416972 603418 417208 603654
rect 416652 603098 416888 603334
rect 416972 603098 417208 603334
rect 452652 603418 452888 603654
rect 452972 603418 453208 603654
rect 452652 603098 452888 603334
rect 452972 603098 453208 603334
rect 488652 603418 488888 603654
rect 488972 603418 489208 603654
rect 488652 603098 488888 603334
rect 488972 603098 489208 603334
rect 524652 603418 524888 603654
rect 524972 603418 525208 603654
rect 524652 603098 524888 603334
rect 524972 603098 525208 603334
rect 560652 603418 560888 603654
rect 560972 603418 561208 603654
rect 560652 603098 560888 603334
rect 560972 603098 561208 603334
rect 570292 603418 570528 603654
rect 570612 603418 570848 603654
rect 570292 603098 570528 603334
rect 570612 603098 570848 603334
rect 585342 603418 585578 603654
rect 585662 603418 585898 603654
rect 585342 603098 585578 603334
rect 585662 603098 585898 603334
rect 7876 583418 8112 583654
rect 8196 583418 8432 583654
rect 7876 583098 8112 583334
rect 8196 583098 8432 583334
rect 38032 583418 38268 583654
rect 38352 583418 38588 583654
rect 38032 583098 38268 583334
rect 38352 583098 38588 583334
rect 74032 583418 74268 583654
rect 74352 583418 74588 583654
rect 74032 583098 74268 583334
rect 74352 583098 74588 583334
rect 110032 583418 110268 583654
rect 110352 583418 110588 583654
rect 110032 583098 110268 583334
rect 110352 583098 110588 583334
rect 146032 583418 146268 583654
rect 146352 583418 146588 583654
rect 146032 583098 146268 583334
rect 146352 583098 146588 583334
rect 182032 583418 182268 583654
rect 182352 583418 182588 583654
rect 182032 583098 182268 583334
rect 182352 583098 182588 583334
rect 218032 583418 218268 583654
rect 218352 583418 218588 583654
rect 218032 583098 218268 583334
rect 218352 583098 218588 583334
rect 254032 583418 254268 583654
rect 254352 583418 254588 583654
rect 254032 583098 254268 583334
rect 254352 583098 254588 583334
rect 290032 583418 290268 583654
rect 290352 583418 290588 583654
rect 290032 583098 290268 583334
rect 290352 583098 290588 583334
rect 326032 583418 326268 583654
rect 326352 583418 326588 583654
rect 326032 583098 326268 583334
rect 326352 583098 326588 583334
rect 362032 583418 362268 583654
rect 362352 583418 362588 583654
rect 362032 583098 362268 583334
rect 362352 583098 362588 583334
rect 398032 583418 398268 583654
rect 398352 583418 398588 583654
rect 398032 583098 398268 583334
rect 398352 583098 398588 583334
rect 434032 583418 434268 583654
rect 434352 583418 434588 583654
rect 434032 583098 434268 583334
rect 434352 583098 434588 583334
rect 470032 583418 470268 583654
rect 470352 583418 470588 583654
rect 470032 583098 470268 583334
rect 470352 583098 470588 583334
rect 506032 583418 506268 583654
rect 506352 583418 506588 583654
rect 506032 583098 506268 583334
rect 506352 583098 506588 583334
rect 542032 583418 542268 583654
rect 542352 583418 542588 583654
rect 542032 583098 542268 583334
rect 542352 583098 542588 583334
rect 571532 583418 571768 583654
rect 571852 583418 572088 583654
rect 571532 583098 571768 583334
rect 571852 583098 572088 583334
rect -1974 563418 -1738 563654
rect -1654 563418 -1418 563654
rect -1974 563098 -1738 563334
rect -1654 563098 -1418 563334
rect 9116 563418 9352 563654
rect 9436 563418 9672 563654
rect 9116 563098 9352 563334
rect 9436 563098 9672 563334
rect 56652 563418 56888 563654
rect 56972 563418 57208 563654
rect 56652 563098 56888 563334
rect 56972 563098 57208 563334
rect 92652 563418 92888 563654
rect 92972 563418 93208 563654
rect 92652 563098 92888 563334
rect 92972 563098 93208 563334
rect 128652 563418 128888 563654
rect 128972 563418 129208 563654
rect 128652 563098 128888 563334
rect 128972 563098 129208 563334
rect 164652 563418 164888 563654
rect 164972 563418 165208 563654
rect 164652 563098 164888 563334
rect 164972 563098 165208 563334
rect 200652 563418 200888 563654
rect 200972 563418 201208 563654
rect 200652 563098 200888 563334
rect 200972 563098 201208 563334
rect 236652 563418 236888 563654
rect 236972 563418 237208 563654
rect 236652 563098 236888 563334
rect 236972 563098 237208 563334
rect 272652 563418 272888 563654
rect 272972 563418 273208 563654
rect 272652 563098 272888 563334
rect 272972 563098 273208 563334
rect 308652 563418 308888 563654
rect 308972 563418 309208 563654
rect 308652 563098 308888 563334
rect 308972 563098 309208 563334
rect 344652 563418 344888 563654
rect 344972 563418 345208 563654
rect 344652 563098 344888 563334
rect 344972 563098 345208 563334
rect 380652 563418 380888 563654
rect 380972 563418 381208 563654
rect 380652 563098 380888 563334
rect 380972 563098 381208 563334
rect 416652 563418 416888 563654
rect 416972 563418 417208 563654
rect 416652 563098 416888 563334
rect 416972 563098 417208 563334
rect 452652 563418 452888 563654
rect 452972 563418 453208 563654
rect 452652 563098 452888 563334
rect 452972 563098 453208 563334
rect 488652 563418 488888 563654
rect 488972 563418 489208 563654
rect 488652 563098 488888 563334
rect 488972 563098 489208 563334
rect 524652 563418 524888 563654
rect 524972 563418 525208 563654
rect 524652 563098 524888 563334
rect 524972 563098 525208 563334
rect 560652 563418 560888 563654
rect 560972 563418 561208 563654
rect 560652 563098 560888 563334
rect 560972 563098 561208 563334
rect 570292 563418 570528 563654
rect 570612 563418 570848 563654
rect 570292 563098 570528 563334
rect 570612 563098 570848 563334
rect 585342 563418 585578 563654
rect 585662 563418 585898 563654
rect 585342 563098 585578 563334
rect 585662 563098 585898 563334
rect 7876 543418 8112 543654
rect 8196 543418 8432 543654
rect 7876 543098 8112 543334
rect 8196 543098 8432 543334
rect 38032 543418 38268 543654
rect 38352 543418 38588 543654
rect 38032 543098 38268 543334
rect 38352 543098 38588 543334
rect 74032 543418 74268 543654
rect 74352 543418 74588 543654
rect 74032 543098 74268 543334
rect 74352 543098 74588 543334
rect 110032 543418 110268 543654
rect 110352 543418 110588 543654
rect 110032 543098 110268 543334
rect 110352 543098 110588 543334
rect 146032 543418 146268 543654
rect 146352 543418 146588 543654
rect 146032 543098 146268 543334
rect 146352 543098 146588 543334
rect 182032 543418 182268 543654
rect 182352 543418 182588 543654
rect 182032 543098 182268 543334
rect 182352 543098 182588 543334
rect 218032 543418 218268 543654
rect 218352 543418 218588 543654
rect 218032 543098 218268 543334
rect 218352 543098 218588 543334
rect 254032 543418 254268 543654
rect 254352 543418 254588 543654
rect 254032 543098 254268 543334
rect 254352 543098 254588 543334
rect 290032 543418 290268 543654
rect 290352 543418 290588 543654
rect 290032 543098 290268 543334
rect 290352 543098 290588 543334
rect 326032 543418 326268 543654
rect 326352 543418 326588 543654
rect 326032 543098 326268 543334
rect 326352 543098 326588 543334
rect 362032 543418 362268 543654
rect 362352 543418 362588 543654
rect 362032 543098 362268 543334
rect 362352 543098 362588 543334
rect 398032 543418 398268 543654
rect 398352 543418 398588 543654
rect 398032 543098 398268 543334
rect 398352 543098 398588 543334
rect 434032 543418 434268 543654
rect 434352 543418 434588 543654
rect 434032 543098 434268 543334
rect 434352 543098 434588 543334
rect 470032 543418 470268 543654
rect 470352 543418 470588 543654
rect 470032 543098 470268 543334
rect 470352 543098 470588 543334
rect 506032 543418 506268 543654
rect 506352 543418 506588 543654
rect 506032 543098 506268 543334
rect 506352 543098 506588 543334
rect 542032 543418 542268 543654
rect 542352 543418 542588 543654
rect 542032 543098 542268 543334
rect 542352 543098 542588 543334
rect 571532 543418 571768 543654
rect 571852 543418 572088 543654
rect 571532 543098 571768 543334
rect 571852 543098 572088 543334
rect -1974 523418 -1738 523654
rect -1654 523418 -1418 523654
rect -1974 523098 -1738 523334
rect -1654 523098 -1418 523334
rect 9116 523418 9352 523654
rect 9436 523418 9672 523654
rect 9116 523098 9352 523334
rect 9436 523098 9672 523334
rect 56652 523418 56888 523654
rect 56972 523418 57208 523654
rect 56652 523098 56888 523334
rect 56972 523098 57208 523334
rect 92652 523418 92888 523654
rect 92972 523418 93208 523654
rect 92652 523098 92888 523334
rect 92972 523098 93208 523334
rect 128652 523418 128888 523654
rect 128972 523418 129208 523654
rect 128652 523098 128888 523334
rect 128972 523098 129208 523334
rect 164652 523418 164888 523654
rect 164972 523418 165208 523654
rect 164652 523098 164888 523334
rect 164972 523098 165208 523334
rect 200652 523418 200888 523654
rect 200972 523418 201208 523654
rect 200652 523098 200888 523334
rect 200972 523098 201208 523334
rect 236652 523418 236888 523654
rect 236972 523418 237208 523654
rect 236652 523098 236888 523334
rect 236972 523098 237208 523334
rect 272652 523418 272888 523654
rect 272972 523418 273208 523654
rect 272652 523098 272888 523334
rect 272972 523098 273208 523334
rect 308652 523418 308888 523654
rect 308972 523418 309208 523654
rect 308652 523098 308888 523334
rect 308972 523098 309208 523334
rect 344652 523418 344888 523654
rect 344972 523418 345208 523654
rect 344652 523098 344888 523334
rect 344972 523098 345208 523334
rect 380652 523418 380888 523654
rect 380972 523418 381208 523654
rect 380652 523098 380888 523334
rect 380972 523098 381208 523334
rect 416652 523418 416888 523654
rect 416972 523418 417208 523654
rect 416652 523098 416888 523334
rect 416972 523098 417208 523334
rect 452652 523418 452888 523654
rect 452972 523418 453208 523654
rect 452652 523098 452888 523334
rect 452972 523098 453208 523334
rect 488652 523418 488888 523654
rect 488972 523418 489208 523654
rect 488652 523098 488888 523334
rect 488972 523098 489208 523334
rect 524652 523418 524888 523654
rect 524972 523418 525208 523654
rect 524652 523098 524888 523334
rect 524972 523098 525208 523334
rect 560652 523418 560888 523654
rect 560972 523418 561208 523654
rect 560652 523098 560888 523334
rect 560972 523098 561208 523334
rect 570292 523418 570528 523654
rect 570612 523418 570848 523654
rect 570292 523098 570528 523334
rect 570612 523098 570848 523334
rect 585342 523418 585578 523654
rect 585662 523418 585898 523654
rect 585342 523098 585578 523334
rect 585662 523098 585898 523334
rect 7876 503418 8112 503654
rect 8196 503418 8432 503654
rect 7876 503098 8112 503334
rect 8196 503098 8432 503334
rect 38032 503418 38268 503654
rect 38352 503418 38588 503654
rect 38032 503098 38268 503334
rect 38352 503098 38588 503334
rect 60622 503418 60858 503654
rect 60622 503098 60858 503334
rect 159098 503418 159334 503654
rect 159098 503098 159334 503334
rect 182032 503418 182268 503654
rect 182352 503418 182588 503654
rect 182032 503098 182268 503334
rect 182352 503098 182588 503334
rect 185622 503418 185858 503654
rect 185622 503098 185858 503334
rect 284098 503418 284334 503654
rect 284098 503098 284334 503334
rect 290032 503418 290268 503654
rect 290352 503418 290588 503654
rect 290032 503098 290268 503334
rect 290352 503098 290588 503334
rect 310622 503418 310858 503654
rect 310622 503098 310858 503334
rect 409098 503418 409334 503654
rect 409098 503098 409334 503334
rect 434032 503418 434268 503654
rect 434352 503418 434588 503654
rect 434032 503098 434268 503334
rect 434352 503098 434588 503334
rect 436622 503418 436858 503654
rect 436622 503098 436858 503334
rect 535098 503418 535334 503654
rect 535098 503098 535334 503334
rect 542032 503418 542268 503654
rect 542352 503418 542588 503654
rect 542032 503098 542268 503334
rect 542352 503098 542588 503334
rect 571532 503418 571768 503654
rect 571852 503418 572088 503654
rect 571532 503098 571768 503334
rect 571852 503098 572088 503334
rect -1974 483418 -1738 483654
rect -1654 483418 -1418 483654
rect -1974 483098 -1738 483334
rect -1654 483098 -1418 483334
rect 9116 483418 9352 483654
rect 9436 483418 9672 483654
rect 9116 483098 9352 483334
rect 9436 483098 9672 483334
rect 56652 483418 56888 483654
rect 56972 483418 57208 483654
rect 56652 483098 56888 483334
rect 56972 483098 57208 483334
rect 61342 483418 61578 483654
rect 61342 483098 61578 483334
rect 158378 483418 158614 483654
rect 158378 483098 158614 483334
rect 164652 483418 164888 483654
rect 164972 483418 165208 483654
rect 164652 483098 164888 483334
rect 164972 483098 165208 483334
rect 186342 483418 186578 483654
rect 186342 483098 186578 483334
rect 283378 483418 283614 483654
rect 283378 483098 283614 483334
rect 308652 483418 308888 483654
rect 308972 483418 309208 483654
rect 308652 483098 308888 483334
rect 308972 483098 309208 483334
rect 311342 483418 311578 483654
rect 311342 483098 311578 483334
rect 408378 483418 408614 483654
rect 408378 483098 408614 483334
rect 416652 483418 416888 483654
rect 416972 483418 417208 483654
rect 416652 483098 416888 483334
rect 416972 483098 417208 483334
rect 437342 483418 437578 483654
rect 437342 483098 437578 483334
rect 534378 483418 534614 483654
rect 534378 483098 534614 483334
rect 560652 483418 560888 483654
rect 560972 483418 561208 483654
rect 560652 483098 560888 483334
rect 560972 483098 561208 483334
rect 570292 483418 570528 483654
rect 570612 483418 570848 483654
rect 570292 483098 570528 483334
rect 570612 483098 570848 483334
rect 585342 483418 585578 483654
rect 585662 483418 585898 483654
rect 585342 483098 585578 483334
rect 585662 483098 585898 483334
rect 7876 463418 8112 463654
rect 8196 463418 8432 463654
rect 7876 463098 8112 463334
rect 8196 463098 8432 463334
rect 38032 463418 38268 463654
rect 38352 463418 38588 463654
rect 38032 463098 38268 463334
rect 38352 463098 38588 463334
rect 60622 463418 60858 463654
rect 60622 463098 60858 463334
rect 159098 463418 159334 463654
rect 159098 463098 159334 463334
rect 182032 463418 182268 463654
rect 182352 463418 182588 463654
rect 182032 463098 182268 463334
rect 182352 463098 182588 463334
rect 185622 463418 185858 463654
rect 185622 463098 185858 463334
rect 284098 463418 284334 463654
rect 284098 463098 284334 463334
rect 290032 463418 290268 463654
rect 290352 463418 290588 463654
rect 290032 463098 290268 463334
rect 290352 463098 290588 463334
rect 310622 463418 310858 463654
rect 310622 463098 310858 463334
rect 409098 463418 409334 463654
rect 409098 463098 409334 463334
rect 434032 463418 434268 463654
rect 434352 463418 434588 463654
rect 434032 463098 434268 463334
rect 434352 463098 434588 463334
rect 436622 463418 436858 463654
rect 436622 463098 436858 463334
rect 535098 463418 535334 463654
rect 535098 463098 535334 463334
rect 542032 463418 542268 463654
rect 542352 463418 542588 463654
rect 542032 463098 542268 463334
rect 542352 463098 542588 463334
rect 571532 463418 571768 463654
rect 571852 463418 572088 463654
rect 571532 463098 571768 463334
rect 571852 463098 572088 463334
rect -1974 443418 -1738 443654
rect -1654 443418 -1418 443654
rect -1974 443098 -1738 443334
rect -1654 443098 -1418 443334
rect 9116 443418 9352 443654
rect 9436 443418 9672 443654
rect 9116 443098 9352 443334
rect 9436 443098 9672 443334
rect 56652 443418 56888 443654
rect 56972 443418 57208 443654
rect 56652 443098 56888 443334
rect 56972 443098 57208 443334
rect 61342 443418 61578 443654
rect 61342 443098 61578 443334
rect 158378 443418 158614 443654
rect 158378 443098 158614 443334
rect 164652 443418 164888 443654
rect 164972 443418 165208 443654
rect 164652 443098 164888 443334
rect 164972 443098 165208 443334
rect 186342 443418 186578 443654
rect 186342 443098 186578 443334
rect 283378 443418 283614 443654
rect 283378 443098 283614 443334
rect 308652 443418 308888 443654
rect 308972 443418 309208 443654
rect 308652 443098 308888 443334
rect 308972 443098 309208 443334
rect 311342 443418 311578 443654
rect 311342 443098 311578 443334
rect 408378 443418 408614 443654
rect 408378 443098 408614 443334
rect 416652 443418 416888 443654
rect 416972 443418 417208 443654
rect 416652 443098 416888 443334
rect 416972 443098 417208 443334
rect 437342 443418 437578 443654
rect 437342 443098 437578 443334
rect 534378 443418 534614 443654
rect 534378 443098 534614 443334
rect 560652 443418 560888 443654
rect 560972 443418 561208 443654
rect 560652 443098 560888 443334
rect 560972 443098 561208 443334
rect 570292 443418 570528 443654
rect 570612 443418 570848 443654
rect 570292 443098 570528 443334
rect 570612 443098 570848 443334
rect 585342 443418 585578 443654
rect 585662 443418 585898 443654
rect 585342 443098 585578 443334
rect 585662 443098 585898 443334
rect 7876 423418 8112 423654
rect 8196 423418 8432 423654
rect 7876 423098 8112 423334
rect 8196 423098 8432 423334
rect 38032 423418 38268 423654
rect 38352 423418 38588 423654
rect 38032 423098 38268 423334
rect 38352 423098 38588 423334
rect 74032 423418 74268 423654
rect 74352 423418 74588 423654
rect 74032 423098 74268 423334
rect 74352 423098 74588 423334
rect 110032 423418 110268 423654
rect 110352 423418 110588 423654
rect 110032 423098 110268 423334
rect 110352 423098 110588 423334
rect 146032 423418 146268 423654
rect 146352 423418 146588 423654
rect 146032 423098 146268 423334
rect 146352 423098 146588 423334
rect 182032 423418 182268 423654
rect 182352 423418 182588 423654
rect 182032 423098 182268 423334
rect 182352 423098 182588 423334
rect 218032 423418 218268 423654
rect 218352 423418 218588 423654
rect 218032 423098 218268 423334
rect 218352 423098 218588 423334
rect 254032 423418 254268 423654
rect 254352 423418 254588 423654
rect 254032 423098 254268 423334
rect 254352 423098 254588 423334
rect 290032 423418 290268 423654
rect 290352 423418 290588 423654
rect 290032 423098 290268 423334
rect 290352 423098 290588 423334
rect 326032 423418 326268 423654
rect 326352 423418 326588 423654
rect 326032 423098 326268 423334
rect 326352 423098 326588 423334
rect 362032 423418 362268 423654
rect 362352 423418 362588 423654
rect 362032 423098 362268 423334
rect 362352 423098 362588 423334
rect 398032 423418 398268 423654
rect 398352 423418 398588 423654
rect 398032 423098 398268 423334
rect 398352 423098 398588 423334
rect 434032 423418 434268 423654
rect 434352 423418 434588 423654
rect 434032 423098 434268 423334
rect 434352 423098 434588 423334
rect 470032 423418 470268 423654
rect 470352 423418 470588 423654
rect 470032 423098 470268 423334
rect 470352 423098 470588 423334
rect 506032 423418 506268 423654
rect 506352 423418 506588 423654
rect 506032 423098 506268 423334
rect 506352 423098 506588 423334
rect 542032 423418 542268 423654
rect 542352 423418 542588 423654
rect 542032 423098 542268 423334
rect 542352 423098 542588 423334
rect 571532 423418 571768 423654
rect 571852 423418 572088 423654
rect 571532 423098 571768 423334
rect 571852 423098 572088 423334
rect -1974 403418 -1738 403654
rect -1654 403418 -1418 403654
rect -1974 403098 -1738 403334
rect -1654 403098 -1418 403334
rect 9116 403418 9352 403654
rect 9436 403418 9672 403654
rect 9116 403098 9352 403334
rect 9436 403098 9672 403334
rect 56652 403418 56888 403654
rect 56972 403418 57208 403654
rect 56652 403098 56888 403334
rect 56972 403098 57208 403334
rect 92652 403418 92888 403654
rect 92972 403418 93208 403654
rect 92652 403098 92888 403334
rect 92972 403098 93208 403334
rect 128652 403418 128888 403654
rect 128972 403418 129208 403654
rect 128652 403098 128888 403334
rect 128972 403098 129208 403334
rect 164652 403418 164888 403654
rect 164972 403418 165208 403654
rect 164652 403098 164888 403334
rect 164972 403098 165208 403334
rect 200652 403418 200888 403654
rect 200972 403418 201208 403654
rect 200652 403098 200888 403334
rect 200972 403098 201208 403334
rect 236652 403418 236888 403654
rect 236972 403418 237208 403654
rect 236652 403098 236888 403334
rect 236972 403098 237208 403334
rect 272652 403418 272888 403654
rect 272972 403418 273208 403654
rect 272652 403098 272888 403334
rect 272972 403098 273208 403334
rect 308652 403418 308888 403654
rect 308972 403418 309208 403654
rect 308652 403098 308888 403334
rect 308972 403098 309208 403334
rect 344652 403418 344888 403654
rect 344972 403418 345208 403654
rect 344652 403098 344888 403334
rect 344972 403098 345208 403334
rect 380652 403418 380888 403654
rect 380972 403418 381208 403654
rect 380652 403098 380888 403334
rect 380972 403098 381208 403334
rect 416652 403418 416888 403654
rect 416972 403418 417208 403654
rect 416652 403098 416888 403334
rect 416972 403098 417208 403334
rect 452652 403418 452888 403654
rect 452972 403418 453208 403654
rect 452652 403098 452888 403334
rect 452972 403098 453208 403334
rect 488652 403418 488888 403654
rect 488972 403418 489208 403654
rect 488652 403098 488888 403334
rect 488972 403098 489208 403334
rect 524652 403418 524888 403654
rect 524972 403418 525208 403654
rect 524652 403098 524888 403334
rect 524972 403098 525208 403334
rect 560652 403418 560888 403654
rect 560972 403418 561208 403654
rect 560652 403098 560888 403334
rect 560972 403098 561208 403334
rect 570292 403418 570528 403654
rect 570612 403418 570848 403654
rect 570292 403098 570528 403334
rect 570612 403098 570848 403334
rect 585342 403418 585578 403654
rect 585662 403418 585898 403654
rect 585342 403098 585578 403334
rect 585662 403098 585898 403334
rect 7876 383418 8112 383654
rect 8196 383418 8432 383654
rect 7876 383098 8112 383334
rect 8196 383098 8432 383334
rect 38032 383418 38268 383654
rect 38352 383418 38588 383654
rect 38032 383098 38268 383334
rect 38352 383098 38588 383334
rect 74032 383418 74268 383654
rect 74352 383418 74588 383654
rect 74032 383098 74268 383334
rect 74352 383098 74588 383334
rect 110032 383418 110268 383654
rect 110352 383418 110588 383654
rect 110032 383098 110268 383334
rect 110352 383098 110588 383334
rect 146032 383418 146268 383654
rect 146352 383418 146588 383654
rect 146032 383098 146268 383334
rect 146352 383098 146588 383334
rect 182032 383418 182268 383654
rect 182352 383418 182588 383654
rect 182032 383098 182268 383334
rect 182352 383098 182588 383334
rect 218032 383418 218268 383654
rect 218352 383418 218588 383654
rect 218032 383098 218268 383334
rect 218352 383098 218588 383334
rect 254032 383418 254268 383654
rect 254352 383418 254588 383654
rect 254032 383098 254268 383334
rect 254352 383098 254588 383334
rect 290032 383418 290268 383654
rect 290352 383418 290588 383654
rect 290032 383098 290268 383334
rect 290352 383098 290588 383334
rect 326032 383418 326268 383654
rect 326352 383418 326588 383654
rect 326032 383098 326268 383334
rect 326352 383098 326588 383334
rect 362032 383418 362268 383654
rect 362352 383418 362588 383654
rect 362032 383098 362268 383334
rect 362352 383098 362588 383334
rect 398032 383418 398268 383654
rect 398352 383418 398588 383654
rect 398032 383098 398268 383334
rect 398352 383098 398588 383334
rect 434032 383418 434268 383654
rect 434352 383418 434588 383654
rect 434032 383098 434268 383334
rect 434352 383098 434588 383334
rect 470032 383418 470268 383654
rect 470352 383418 470588 383654
rect 470032 383098 470268 383334
rect 470352 383098 470588 383334
rect 506032 383418 506268 383654
rect 506352 383418 506588 383654
rect 506032 383098 506268 383334
rect 506352 383098 506588 383334
rect 542032 383418 542268 383654
rect 542352 383418 542588 383654
rect 542032 383098 542268 383334
rect 542352 383098 542588 383334
rect 571532 383418 571768 383654
rect 571852 383418 572088 383654
rect 571532 383098 571768 383334
rect 571852 383098 572088 383334
rect -1974 363418 -1738 363654
rect -1654 363418 -1418 363654
rect -1974 363098 -1738 363334
rect -1654 363098 -1418 363334
rect 9116 363418 9352 363654
rect 9436 363418 9672 363654
rect 9116 363098 9352 363334
rect 9436 363098 9672 363334
rect 56652 363418 56888 363654
rect 56972 363418 57208 363654
rect 56652 363098 56888 363334
rect 56972 363098 57208 363334
rect 92652 363418 92888 363654
rect 92972 363418 93208 363654
rect 92652 363098 92888 363334
rect 92972 363098 93208 363334
rect 128652 363418 128888 363654
rect 128972 363418 129208 363654
rect 128652 363098 128888 363334
rect 128972 363098 129208 363334
rect 164652 363418 164888 363654
rect 164972 363418 165208 363654
rect 164652 363098 164888 363334
rect 164972 363098 165208 363334
rect 200652 363418 200888 363654
rect 200972 363418 201208 363654
rect 200652 363098 200888 363334
rect 200972 363098 201208 363334
rect 236652 363418 236888 363654
rect 236972 363418 237208 363654
rect 236652 363098 236888 363334
rect 236972 363098 237208 363334
rect 272652 363418 272888 363654
rect 272972 363418 273208 363654
rect 272652 363098 272888 363334
rect 272972 363098 273208 363334
rect 308652 363418 308888 363654
rect 308972 363418 309208 363654
rect 308652 363098 308888 363334
rect 308972 363098 309208 363334
rect 344652 363418 344888 363654
rect 344972 363418 345208 363654
rect 344652 363098 344888 363334
rect 344972 363098 345208 363334
rect 380652 363418 380888 363654
rect 380972 363418 381208 363654
rect 380652 363098 380888 363334
rect 380972 363098 381208 363334
rect 416652 363418 416888 363654
rect 416972 363418 417208 363654
rect 416652 363098 416888 363334
rect 416972 363098 417208 363334
rect 452652 363418 452888 363654
rect 452972 363418 453208 363654
rect 452652 363098 452888 363334
rect 452972 363098 453208 363334
rect 488652 363418 488888 363654
rect 488972 363418 489208 363654
rect 488652 363098 488888 363334
rect 488972 363098 489208 363334
rect 524652 363418 524888 363654
rect 524972 363418 525208 363654
rect 524652 363098 524888 363334
rect 524972 363098 525208 363334
rect 560652 363418 560888 363654
rect 560972 363418 561208 363654
rect 560652 363098 560888 363334
rect 560972 363098 561208 363334
rect 570292 363418 570528 363654
rect 570612 363418 570848 363654
rect 570292 363098 570528 363334
rect 570612 363098 570848 363334
rect 585342 363418 585578 363654
rect 585662 363418 585898 363654
rect 585342 363098 585578 363334
rect 585662 363098 585898 363334
rect 7876 343418 8112 343654
rect 8196 343418 8432 343654
rect 7876 343098 8112 343334
rect 8196 343098 8432 343334
rect 38032 343418 38268 343654
rect 38352 343418 38588 343654
rect 38032 343098 38268 343334
rect 38352 343098 38588 343334
rect 74032 343418 74268 343654
rect 74352 343418 74588 343654
rect 74032 343098 74268 343334
rect 74352 343098 74588 343334
rect 110032 343418 110268 343654
rect 110352 343418 110588 343654
rect 110032 343098 110268 343334
rect 110352 343098 110588 343334
rect 146032 343418 146268 343654
rect 146352 343418 146588 343654
rect 146032 343098 146268 343334
rect 146352 343098 146588 343334
rect 182032 343418 182268 343654
rect 182352 343418 182588 343654
rect 182032 343098 182268 343334
rect 182352 343098 182588 343334
rect 218032 343418 218268 343654
rect 218352 343418 218588 343654
rect 218032 343098 218268 343334
rect 218352 343098 218588 343334
rect 254032 343418 254268 343654
rect 254352 343418 254588 343654
rect 254032 343098 254268 343334
rect 254352 343098 254588 343334
rect 290032 343418 290268 343654
rect 290352 343418 290588 343654
rect 290032 343098 290268 343334
rect 290352 343098 290588 343334
rect 326032 343418 326268 343654
rect 326352 343418 326588 343654
rect 326032 343098 326268 343334
rect 326352 343098 326588 343334
rect 362032 343418 362268 343654
rect 362352 343418 362588 343654
rect 362032 343098 362268 343334
rect 362352 343098 362588 343334
rect 398032 343418 398268 343654
rect 398352 343418 398588 343654
rect 398032 343098 398268 343334
rect 398352 343098 398588 343334
rect 434032 343418 434268 343654
rect 434352 343418 434588 343654
rect 434032 343098 434268 343334
rect 434352 343098 434588 343334
rect 470032 343418 470268 343654
rect 470352 343418 470588 343654
rect 470032 343098 470268 343334
rect 470352 343098 470588 343334
rect 506032 343418 506268 343654
rect 506352 343418 506588 343654
rect 506032 343098 506268 343334
rect 506352 343098 506588 343334
rect 542032 343418 542268 343654
rect 542352 343418 542588 343654
rect 542032 343098 542268 343334
rect 542352 343098 542588 343334
rect 571532 343418 571768 343654
rect 571852 343418 572088 343654
rect 571532 343098 571768 343334
rect 571852 343098 572088 343334
rect -1974 323418 -1738 323654
rect -1654 323418 -1418 323654
rect -1974 323098 -1738 323334
rect -1654 323098 -1418 323334
rect 9116 323418 9352 323654
rect 9436 323418 9672 323654
rect 9116 323098 9352 323334
rect 9436 323098 9672 323334
rect 56652 323418 56888 323654
rect 56972 323418 57208 323654
rect 56652 323098 56888 323334
rect 56972 323098 57208 323334
rect 92652 323418 92888 323654
rect 92972 323418 93208 323654
rect 92652 323098 92888 323334
rect 92972 323098 93208 323334
rect 128652 323418 128888 323654
rect 128972 323418 129208 323654
rect 128652 323098 128888 323334
rect 128972 323098 129208 323334
rect 164652 323418 164888 323654
rect 164972 323418 165208 323654
rect 164652 323098 164888 323334
rect 164972 323098 165208 323334
rect 200652 323418 200888 323654
rect 200972 323418 201208 323654
rect 200652 323098 200888 323334
rect 200972 323098 201208 323334
rect 236652 323418 236888 323654
rect 236972 323418 237208 323654
rect 236652 323098 236888 323334
rect 236972 323098 237208 323334
rect 272652 323418 272888 323654
rect 272972 323418 273208 323654
rect 272652 323098 272888 323334
rect 272972 323098 273208 323334
rect 308652 323418 308888 323654
rect 308972 323418 309208 323654
rect 308652 323098 308888 323334
rect 308972 323098 309208 323334
rect 344652 323418 344888 323654
rect 344972 323418 345208 323654
rect 344652 323098 344888 323334
rect 344972 323098 345208 323334
rect 380652 323418 380888 323654
rect 380972 323418 381208 323654
rect 380652 323098 380888 323334
rect 380972 323098 381208 323334
rect 416652 323418 416888 323654
rect 416972 323418 417208 323654
rect 416652 323098 416888 323334
rect 416972 323098 417208 323334
rect 452652 323418 452888 323654
rect 452972 323418 453208 323654
rect 452652 323098 452888 323334
rect 452972 323098 453208 323334
rect 488652 323418 488888 323654
rect 488972 323418 489208 323654
rect 488652 323098 488888 323334
rect 488972 323098 489208 323334
rect 524652 323418 524888 323654
rect 524972 323418 525208 323654
rect 524652 323098 524888 323334
rect 524972 323098 525208 323334
rect 560652 323418 560888 323654
rect 560972 323418 561208 323654
rect 560652 323098 560888 323334
rect 560972 323098 561208 323334
rect 570292 323418 570528 323654
rect 570612 323418 570848 323654
rect 570292 323098 570528 323334
rect 570612 323098 570848 323334
rect 585342 323418 585578 323654
rect 585662 323418 585898 323654
rect 585342 323098 585578 323334
rect 585662 323098 585898 323334
rect 7876 303418 8112 303654
rect 8196 303418 8432 303654
rect 7876 303098 8112 303334
rect 8196 303098 8432 303334
rect 38032 303418 38268 303654
rect 38352 303418 38588 303654
rect 38032 303098 38268 303334
rect 38352 303098 38588 303334
rect 74032 303418 74268 303654
rect 74352 303418 74588 303654
rect 74032 303098 74268 303334
rect 74352 303098 74588 303334
rect 110032 303418 110268 303654
rect 110352 303418 110588 303654
rect 110032 303098 110268 303334
rect 110352 303098 110588 303334
rect 146032 303418 146268 303654
rect 146352 303418 146588 303654
rect 146032 303098 146268 303334
rect 146352 303098 146588 303334
rect 182032 303418 182268 303654
rect 182352 303418 182588 303654
rect 182032 303098 182268 303334
rect 182352 303098 182588 303334
rect 218032 303418 218268 303654
rect 218352 303418 218588 303654
rect 218032 303098 218268 303334
rect 218352 303098 218588 303334
rect 254032 303418 254268 303654
rect 254352 303418 254588 303654
rect 254032 303098 254268 303334
rect 254352 303098 254588 303334
rect 290032 303418 290268 303654
rect 290352 303418 290588 303654
rect 290032 303098 290268 303334
rect 290352 303098 290588 303334
rect 326032 303418 326268 303654
rect 326352 303418 326588 303654
rect 326032 303098 326268 303334
rect 326352 303098 326588 303334
rect 362032 303418 362268 303654
rect 362352 303418 362588 303654
rect 362032 303098 362268 303334
rect 362352 303098 362588 303334
rect 398032 303418 398268 303654
rect 398352 303418 398588 303654
rect 398032 303098 398268 303334
rect 398352 303098 398588 303334
rect 434032 303418 434268 303654
rect 434352 303418 434588 303654
rect 434032 303098 434268 303334
rect 434352 303098 434588 303334
rect 470032 303418 470268 303654
rect 470352 303418 470588 303654
rect 470032 303098 470268 303334
rect 470352 303098 470588 303334
rect 506032 303418 506268 303654
rect 506352 303418 506588 303654
rect 506032 303098 506268 303334
rect 506352 303098 506588 303334
rect 542032 303418 542268 303654
rect 542352 303418 542588 303654
rect 542032 303098 542268 303334
rect 542352 303098 542588 303334
rect 571532 303418 571768 303654
rect 571852 303418 572088 303654
rect 571532 303098 571768 303334
rect 571852 303098 572088 303334
rect -1974 283418 -1738 283654
rect -1654 283418 -1418 283654
rect -1974 283098 -1738 283334
rect -1654 283098 -1418 283334
rect 9116 283418 9352 283654
rect 9436 283418 9672 283654
rect 9116 283098 9352 283334
rect 9436 283098 9672 283334
rect 56652 283418 56888 283654
rect 56972 283418 57208 283654
rect 56652 283098 56888 283334
rect 56972 283098 57208 283334
rect 92652 283418 92888 283654
rect 92972 283418 93208 283654
rect 92652 283098 92888 283334
rect 92972 283098 93208 283334
rect 128652 283418 128888 283654
rect 128972 283418 129208 283654
rect 128652 283098 128888 283334
rect 128972 283098 129208 283334
rect 164652 283418 164888 283654
rect 164972 283418 165208 283654
rect 164652 283098 164888 283334
rect 164972 283098 165208 283334
rect 200652 283418 200888 283654
rect 200972 283418 201208 283654
rect 200652 283098 200888 283334
rect 200972 283098 201208 283334
rect 236652 283418 236888 283654
rect 236972 283418 237208 283654
rect 236652 283098 236888 283334
rect 236972 283098 237208 283334
rect 272652 283418 272888 283654
rect 272972 283418 273208 283654
rect 272652 283098 272888 283334
rect 272972 283098 273208 283334
rect 308652 283418 308888 283654
rect 308972 283418 309208 283654
rect 308652 283098 308888 283334
rect 308972 283098 309208 283334
rect 344652 283418 344888 283654
rect 344972 283418 345208 283654
rect 344652 283098 344888 283334
rect 344972 283098 345208 283334
rect 380652 283418 380888 283654
rect 380972 283418 381208 283654
rect 380652 283098 380888 283334
rect 380972 283098 381208 283334
rect 416652 283418 416888 283654
rect 416972 283418 417208 283654
rect 416652 283098 416888 283334
rect 416972 283098 417208 283334
rect 452652 283418 452888 283654
rect 452972 283418 453208 283654
rect 452652 283098 452888 283334
rect 452972 283098 453208 283334
rect 488652 283418 488888 283654
rect 488972 283418 489208 283654
rect 488652 283098 488888 283334
rect 488972 283098 489208 283334
rect 524652 283418 524888 283654
rect 524972 283418 525208 283654
rect 524652 283098 524888 283334
rect 524972 283098 525208 283334
rect 560652 283418 560888 283654
rect 560972 283418 561208 283654
rect 560652 283098 560888 283334
rect 560972 283098 561208 283334
rect 570292 283418 570528 283654
rect 570612 283418 570848 283654
rect 570292 283098 570528 283334
rect 570612 283098 570848 283334
rect 585342 283418 585578 283654
rect 585662 283418 585898 283654
rect 585342 283098 585578 283334
rect 585662 283098 585898 283334
rect 7876 263418 8112 263654
rect 8196 263418 8432 263654
rect 7876 263098 8112 263334
rect 8196 263098 8432 263334
rect 38032 263418 38268 263654
rect 38352 263418 38588 263654
rect 38032 263098 38268 263334
rect 38352 263098 38588 263334
rect 74032 263418 74268 263654
rect 74352 263418 74588 263654
rect 74032 263098 74268 263334
rect 74352 263098 74588 263334
rect 110032 263418 110268 263654
rect 110352 263418 110588 263654
rect 110032 263098 110268 263334
rect 110352 263098 110588 263334
rect 146032 263418 146268 263654
rect 146352 263418 146588 263654
rect 146032 263098 146268 263334
rect 146352 263098 146588 263334
rect 182032 263418 182268 263654
rect 182352 263418 182588 263654
rect 182032 263098 182268 263334
rect 182352 263098 182588 263334
rect 218032 263418 218268 263654
rect 218352 263418 218588 263654
rect 218032 263098 218268 263334
rect 218352 263098 218588 263334
rect 254032 263418 254268 263654
rect 254352 263418 254588 263654
rect 254032 263098 254268 263334
rect 254352 263098 254588 263334
rect 290032 263418 290268 263654
rect 290352 263418 290588 263654
rect 290032 263098 290268 263334
rect 290352 263098 290588 263334
rect 326032 263418 326268 263654
rect 326352 263418 326588 263654
rect 326032 263098 326268 263334
rect 326352 263098 326588 263334
rect 362032 263418 362268 263654
rect 362352 263418 362588 263654
rect 362032 263098 362268 263334
rect 362352 263098 362588 263334
rect 398032 263418 398268 263654
rect 398352 263418 398588 263654
rect 398032 263098 398268 263334
rect 398352 263098 398588 263334
rect 434032 263418 434268 263654
rect 434352 263418 434588 263654
rect 434032 263098 434268 263334
rect 434352 263098 434588 263334
rect 470032 263418 470268 263654
rect 470352 263418 470588 263654
rect 470032 263098 470268 263334
rect 470352 263098 470588 263334
rect 506032 263418 506268 263654
rect 506352 263418 506588 263654
rect 506032 263098 506268 263334
rect 506352 263098 506588 263334
rect 542032 263418 542268 263654
rect 542352 263418 542588 263654
rect 542032 263098 542268 263334
rect 542352 263098 542588 263334
rect 571532 263418 571768 263654
rect 571852 263418 572088 263654
rect 571532 263098 571768 263334
rect 571852 263098 572088 263334
rect -1974 243418 -1738 243654
rect -1654 243418 -1418 243654
rect -1974 243098 -1738 243334
rect -1654 243098 -1418 243334
rect 9116 243418 9352 243654
rect 9436 243418 9672 243654
rect 9116 243098 9352 243334
rect 9436 243098 9672 243334
rect 56652 243418 56888 243654
rect 56972 243418 57208 243654
rect 56652 243098 56888 243334
rect 56972 243098 57208 243334
rect 92652 243418 92888 243654
rect 92972 243418 93208 243654
rect 92652 243098 92888 243334
rect 92972 243098 93208 243334
rect 128652 243418 128888 243654
rect 128972 243418 129208 243654
rect 128652 243098 128888 243334
rect 128972 243098 129208 243334
rect 164652 243418 164888 243654
rect 164972 243418 165208 243654
rect 164652 243098 164888 243334
rect 164972 243098 165208 243334
rect 200652 243418 200888 243654
rect 200972 243418 201208 243654
rect 200652 243098 200888 243334
rect 200972 243098 201208 243334
rect 236652 243418 236888 243654
rect 236972 243418 237208 243654
rect 236652 243098 236888 243334
rect 236972 243098 237208 243334
rect 272652 243418 272888 243654
rect 272972 243418 273208 243654
rect 272652 243098 272888 243334
rect 272972 243098 273208 243334
rect 308652 243418 308888 243654
rect 308972 243418 309208 243654
rect 308652 243098 308888 243334
rect 308972 243098 309208 243334
rect 344652 243418 344888 243654
rect 344972 243418 345208 243654
rect 344652 243098 344888 243334
rect 344972 243098 345208 243334
rect 380652 243418 380888 243654
rect 380972 243418 381208 243654
rect 380652 243098 380888 243334
rect 380972 243098 381208 243334
rect 416652 243418 416888 243654
rect 416972 243418 417208 243654
rect 416652 243098 416888 243334
rect 416972 243098 417208 243334
rect 452652 243418 452888 243654
rect 452972 243418 453208 243654
rect 452652 243098 452888 243334
rect 452972 243098 453208 243334
rect 488652 243418 488888 243654
rect 488972 243418 489208 243654
rect 488652 243098 488888 243334
rect 488972 243098 489208 243334
rect 524652 243418 524888 243654
rect 524972 243418 525208 243654
rect 524652 243098 524888 243334
rect 524972 243098 525208 243334
rect 560652 243418 560888 243654
rect 560972 243418 561208 243654
rect 560652 243098 560888 243334
rect 560972 243098 561208 243334
rect 570292 243418 570528 243654
rect 570612 243418 570848 243654
rect 570292 243098 570528 243334
rect 570612 243098 570848 243334
rect 585342 243418 585578 243654
rect 585662 243418 585898 243654
rect 585342 243098 585578 243334
rect 585662 243098 585898 243334
rect 7876 223418 8112 223654
rect 8196 223418 8432 223654
rect 7876 223098 8112 223334
rect 8196 223098 8432 223334
rect 38032 223418 38268 223654
rect 38352 223418 38588 223654
rect 38032 223098 38268 223334
rect 38352 223098 38588 223334
rect 74032 223418 74268 223654
rect 74352 223418 74588 223654
rect 74032 223098 74268 223334
rect 74352 223098 74588 223334
rect 110032 223418 110268 223654
rect 110352 223418 110588 223654
rect 110032 223098 110268 223334
rect 110352 223098 110588 223334
rect 146032 223418 146268 223654
rect 146352 223418 146588 223654
rect 146032 223098 146268 223334
rect 146352 223098 146588 223334
rect 182032 223418 182268 223654
rect 182352 223418 182588 223654
rect 182032 223098 182268 223334
rect 182352 223098 182588 223334
rect 218032 223418 218268 223654
rect 218352 223418 218588 223654
rect 218032 223098 218268 223334
rect 218352 223098 218588 223334
rect 254032 223418 254268 223654
rect 254352 223418 254588 223654
rect 254032 223098 254268 223334
rect 254352 223098 254588 223334
rect 290032 223418 290268 223654
rect 290352 223418 290588 223654
rect 290032 223098 290268 223334
rect 290352 223098 290588 223334
rect 326032 223418 326268 223654
rect 326352 223418 326588 223654
rect 326032 223098 326268 223334
rect 326352 223098 326588 223334
rect 362032 223418 362268 223654
rect 362352 223418 362588 223654
rect 362032 223098 362268 223334
rect 362352 223098 362588 223334
rect 398032 223418 398268 223654
rect 398352 223418 398588 223654
rect 398032 223098 398268 223334
rect 398352 223098 398588 223334
rect 434032 223418 434268 223654
rect 434352 223418 434588 223654
rect 434032 223098 434268 223334
rect 434352 223098 434588 223334
rect 470032 223418 470268 223654
rect 470352 223418 470588 223654
rect 470032 223098 470268 223334
rect 470352 223098 470588 223334
rect 506032 223418 506268 223654
rect 506352 223418 506588 223654
rect 506032 223098 506268 223334
rect 506352 223098 506588 223334
rect 542032 223418 542268 223654
rect 542352 223418 542588 223654
rect 542032 223098 542268 223334
rect 542352 223098 542588 223334
rect 571532 223418 571768 223654
rect 571852 223418 572088 223654
rect 571532 223098 571768 223334
rect 571852 223098 572088 223334
rect -1974 203418 -1738 203654
rect -1654 203418 -1418 203654
rect -1974 203098 -1738 203334
rect -1654 203098 -1418 203334
rect 9116 203418 9352 203654
rect 9436 203418 9672 203654
rect 9116 203098 9352 203334
rect 9436 203098 9672 203334
rect 56652 203418 56888 203654
rect 56972 203418 57208 203654
rect 56652 203098 56888 203334
rect 56972 203098 57208 203334
rect 92652 203418 92888 203654
rect 92972 203418 93208 203654
rect 92652 203098 92888 203334
rect 92972 203098 93208 203334
rect 128652 203418 128888 203654
rect 128972 203418 129208 203654
rect 128652 203098 128888 203334
rect 128972 203098 129208 203334
rect 164652 203418 164888 203654
rect 164972 203418 165208 203654
rect 164652 203098 164888 203334
rect 164972 203098 165208 203334
rect 200652 203418 200888 203654
rect 200972 203418 201208 203654
rect 200652 203098 200888 203334
rect 200972 203098 201208 203334
rect 236652 203418 236888 203654
rect 236972 203418 237208 203654
rect 236652 203098 236888 203334
rect 236972 203098 237208 203334
rect 272652 203418 272888 203654
rect 272972 203418 273208 203654
rect 272652 203098 272888 203334
rect 272972 203098 273208 203334
rect 308652 203418 308888 203654
rect 308972 203418 309208 203654
rect 308652 203098 308888 203334
rect 308972 203098 309208 203334
rect 344652 203418 344888 203654
rect 344972 203418 345208 203654
rect 344652 203098 344888 203334
rect 344972 203098 345208 203334
rect 380652 203418 380888 203654
rect 380972 203418 381208 203654
rect 380652 203098 380888 203334
rect 380972 203098 381208 203334
rect 416652 203418 416888 203654
rect 416972 203418 417208 203654
rect 416652 203098 416888 203334
rect 416972 203098 417208 203334
rect 452652 203418 452888 203654
rect 452972 203418 453208 203654
rect 452652 203098 452888 203334
rect 452972 203098 453208 203334
rect 488652 203418 488888 203654
rect 488972 203418 489208 203654
rect 488652 203098 488888 203334
rect 488972 203098 489208 203334
rect 524652 203418 524888 203654
rect 524972 203418 525208 203654
rect 524652 203098 524888 203334
rect 524972 203098 525208 203334
rect 560652 203418 560888 203654
rect 560972 203418 561208 203654
rect 560652 203098 560888 203334
rect 560972 203098 561208 203334
rect 570292 203418 570528 203654
rect 570612 203418 570848 203654
rect 570292 203098 570528 203334
rect 570612 203098 570848 203334
rect 585342 203418 585578 203654
rect 585662 203418 585898 203654
rect 585342 203098 585578 203334
rect 585662 203098 585898 203334
rect 7876 183418 8112 183654
rect 8196 183418 8432 183654
rect 7876 183098 8112 183334
rect 8196 183098 8432 183334
rect 38032 183418 38268 183654
rect 38352 183418 38588 183654
rect 38032 183098 38268 183334
rect 38352 183098 38588 183334
rect 60622 183418 60858 183654
rect 60622 183098 60858 183334
rect 159098 183418 159334 183654
rect 159098 183098 159334 183334
rect 182032 183418 182268 183654
rect 182352 183418 182588 183654
rect 182032 183098 182268 183334
rect 182352 183098 182588 183334
rect 185622 183418 185858 183654
rect 185622 183098 185858 183334
rect 284098 183418 284334 183654
rect 284098 183098 284334 183334
rect 290032 183418 290268 183654
rect 290352 183418 290588 183654
rect 290032 183098 290268 183334
rect 290352 183098 290588 183334
rect 310622 183418 310858 183654
rect 310622 183098 310858 183334
rect 409098 183418 409334 183654
rect 409098 183098 409334 183334
rect 434032 183418 434268 183654
rect 434352 183418 434588 183654
rect 434032 183098 434268 183334
rect 434352 183098 434588 183334
rect 436622 183418 436858 183654
rect 436622 183098 436858 183334
rect 535098 183418 535334 183654
rect 535098 183098 535334 183334
rect 542032 183418 542268 183654
rect 542352 183418 542588 183654
rect 542032 183098 542268 183334
rect 542352 183098 542588 183334
rect 571532 183418 571768 183654
rect 571852 183418 572088 183654
rect 571532 183098 571768 183334
rect 571852 183098 572088 183334
rect -1974 163418 -1738 163654
rect -1654 163418 -1418 163654
rect -1974 163098 -1738 163334
rect -1654 163098 -1418 163334
rect 9116 163418 9352 163654
rect 9436 163418 9672 163654
rect 9116 163098 9352 163334
rect 9436 163098 9672 163334
rect 56652 163418 56888 163654
rect 56972 163418 57208 163654
rect 56652 163098 56888 163334
rect 56972 163098 57208 163334
rect 61342 163418 61578 163654
rect 61342 163098 61578 163334
rect 158378 163418 158614 163654
rect 158378 163098 158614 163334
rect 164652 163418 164888 163654
rect 164972 163418 165208 163654
rect 164652 163098 164888 163334
rect 164972 163098 165208 163334
rect 186342 163418 186578 163654
rect 186342 163098 186578 163334
rect 283378 163418 283614 163654
rect 283378 163098 283614 163334
rect 308652 163418 308888 163654
rect 308972 163418 309208 163654
rect 308652 163098 308888 163334
rect 308972 163098 309208 163334
rect 311342 163418 311578 163654
rect 311342 163098 311578 163334
rect 408378 163418 408614 163654
rect 408378 163098 408614 163334
rect 416652 163418 416888 163654
rect 416972 163418 417208 163654
rect 416652 163098 416888 163334
rect 416972 163098 417208 163334
rect 437342 163418 437578 163654
rect 437342 163098 437578 163334
rect 534378 163418 534614 163654
rect 534378 163098 534614 163334
rect 560652 163418 560888 163654
rect 560972 163418 561208 163654
rect 560652 163098 560888 163334
rect 560972 163098 561208 163334
rect 570292 163418 570528 163654
rect 570612 163418 570848 163654
rect 570292 163098 570528 163334
rect 570612 163098 570848 163334
rect 585342 163418 585578 163654
rect 585662 163418 585898 163654
rect 585342 163098 585578 163334
rect 585662 163098 585898 163334
rect 7876 143418 8112 143654
rect 8196 143418 8432 143654
rect 7876 143098 8112 143334
rect 8196 143098 8432 143334
rect 38032 143418 38268 143654
rect 38352 143418 38588 143654
rect 38032 143098 38268 143334
rect 38352 143098 38588 143334
rect 60622 143418 60858 143654
rect 60622 143098 60858 143334
rect 159098 143418 159334 143654
rect 159098 143098 159334 143334
rect 182032 143418 182268 143654
rect 182352 143418 182588 143654
rect 182032 143098 182268 143334
rect 182352 143098 182588 143334
rect 185622 143418 185858 143654
rect 185622 143098 185858 143334
rect 284098 143418 284334 143654
rect 284098 143098 284334 143334
rect 290032 143418 290268 143654
rect 290352 143418 290588 143654
rect 290032 143098 290268 143334
rect 290352 143098 290588 143334
rect 310622 143418 310858 143654
rect 310622 143098 310858 143334
rect 409098 143418 409334 143654
rect 409098 143098 409334 143334
rect 434032 143418 434268 143654
rect 434352 143418 434588 143654
rect 434032 143098 434268 143334
rect 434352 143098 434588 143334
rect 436622 143418 436858 143654
rect 436622 143098 436858 143334
rect 535098 143418 535334 143654
rect 535098 143098 535334 143334
rect 542032 143418 542268 143654
rect 542352 143418 542588 143654
rect 542032 143098 542268 143334
rect 542352 143098 542588 143334
rect 571532 143418 571768 143654
rect 571852 143418 572088 143654
rect 571532 143098 571768 143334
rect 571852 143098 572088 143334
rect -1974 123418 -1738 123654
rect -1654 123418 -1418 123654
rect -1974 123098 -1738 123334
rect -1654 123098 -1418 123334
rect 9116 123418 9352 123654
rect 9436 123418 9672 123654
rect 9116 123098 9352 123334
rect 9436 123098 9672 123334
rect 56652 123418 56888 123654
rect 56972 123418 57208 123654
rect 56652 123098 56888 123334
rect 56972 123098 57208 123334
rect 61342 123418 61578 123654
rect 61342 123098 61578 123334
rect 158378 123418 158614 123654
rect 158378 123098 158614 123334
rect 164652 123418 164888 123654
rect 164972 123418 165208 123654
rect 164652 123098 164888 123334
rect 164972 123098 165208 123334
rect 186342 123418 186578 123654
rect 186342 123098 186578 123334
rect 283378 123418 283614 123654
rect 283378 123098 283614 123334
rect 308652 123418 308888 123654
rect 308972 123418 309208 123654
rect 308652 123098 308888 123334
rect 308972 123098 309208 123334
rect 311342 123418 311578 123654
rect 311342 123098 311578 123334
rect 408378 123418 408614 123654
rect 408378 123098 408614 123334
rect 416652 123418 416888 123654
rect 416972 123418 417208 123654
rect 416652 123098 416888 123334
rect 416972 123098 417208 123334
rect 437342 123418 437578 123654
rect 437342 123098 437578 123334
rect 534378 123418 534614 123654
rect 534378 123098 534614 123334
rect 560652 123418 560888 123654
rect 560972 123418 561208 123654
rect 560652 123098 560888 123334
rect 560972 123098 561208 123334
rect 570292 123418 570528 123654
rect 570612 123418 570848 123654
rect 570292 123098 570528 123334
rect 570612 123098 570848 123334
rect 585342 123418 585578 123654
rect 585662 123418 585898 123654
rect 585342 123098 585578 123334
rect 585662 123098 585898 123334
rect 7876 103418 8112 103654
rect 8196 103418 8432 103654
rect 7876 103098 8112 103334
rect 8196 103098 8432 103334
rect 38032 103418 38268 103654
rect 38352 103418 38588 103654
rect 38032 103098 38268 103334
rect 38352 103098 38588 103334
rect 74032 103418 74268 103654
rect 74352 103418 74588 103654
rect 74032 103098 74268 103334
rect 74352 103098 74588 103334
rect 110032 103418 110268 103654
rect 110352 103418 110588 103654
rect 110032 103098 110268 103334
rect 110352 103098 110588 103334
rect 146032 103418 146268 103654
rect 146352 103418 146588 103654
rect 146032 103098 146268 103334
rect 146352 103098 146588 103334
rect 182032 103418 182268 103654
rect 182352 103418 182588 103654
rect 182032 103098 182268 103334
rect 182352 103098 182588 103334
rect 218032 103418 218268 103654
rect 218352 103418 218588 103654
rect 218032 103098 218268 103334
rect 218352 103098 218588 103334
rect 254032 103418 254268 103654
rect 254352 103418 254588 103654
rect 254032 103098 254268 103334
rect 254352 103098 254588 103334
rect 290032 103418 290268 103654
rect 290352 103418 290588 103654
rect 290032 103098 290268 103334
rect 290352 103098 290588 103334
rect 326032 103418 326268 103654
rect 326352 103418 326588 103654
rect 326032 103098 326268 103334
rect 326352 103098 326588 103334
rect 362032 103418 362268 103654
rect 362352 103418 362588 103654
rect 362032 103098 362268 103334
rect 362352 103098 362588 103334
rect 398032 103418 398268 103654
rect 398352 103418 398588 103654
rect 398032 103098 398268 103334
rect 398352 103098 398588 103334
rect 434032 103418 434268 103654
rect 434352 103418 434588 103654
rect 434032 103098 434268 103334
rect 434352 103098 434588 103334
rect 470032 103418 470268 103654
rect 470352 103418 470588 103654
rect 470032 103098 470268 103334
rect 470352 103098 470588 103334
rect 506032 103418 506268 103654
rect 506352 103418 506588 103654
rect 506032 103098 506268 103334
rect 506352 103098 506588 103334
rect 542032 103418 542268 103654
rect 542352 103418 542588 103654
rect 542032 103098 542268 103334
rect 542352 103098 542588 103334
rect 571532 103418 571768 103654
rect 571852 103418 572088 103654
rect 571532 103098 571768 103334
rect 571852 103098 572088 103334
rect -1974 83418 -1738 83654
rect -1654 83418 -1418 83654
rect -1974 83098 -1738 83334
rect -1654 83098 -1418 83334
rect 9116 83418 9352 83654
rect 9436 83418 9672 83654
rect 9116 83098 9352 83334
rect 9436 83098 9672 83334
rect 56652 83418 56888 83654
rect 56972 83418 57208 83654
rect 56652 83098 56888 83334
rect 56972 83098 57208 83334
rect 61342 83418 61578 83654
rect 61342 83098 61578 83334
rect 158378 83418 158614 83654
rect 158378 83098 158614 83334
rect 164652 83418 164888 83654
rect 164972 83418 165208 83654
rect 164652 83098 164888 83334
rect 164972 83098 165208 83334
rect 186342 83418 186578 83654
rect 186342 83098 186578 83334
rect 283378 83418 283614 83654
rect 283378 83098 283614 83334
rect 308652 83418 308888 83654
rect 308972 83418 309208 83654
rect 308652 83098 308888 83334
rect 308972 83098 309208 83334
rect 311342 83418 311578 83654
rect 311342 83098 311578 83334
rect 408378 83418 408614 83654
rect 408378 83098 408614 83334
rect 416652 83418 416888 83654
rect 416972 83418 417208 83654
rect 416652 83098 416888 83334
rect 416972 83098 417208 83334
rect 437342 83418 437578 83654
rect 437342 83098 437578 83334
rect 534378 83418 534614 83654
rect 534378 83098 534614 83334
rect 560652 83418 560888 83654
rect 560972 83418 561208 83654
rect 560652 83098 560888 83334
rect 560972 83098 561208 83334
rect 570292 83418 570528 83654
rect 570612 83418 570848 83654
rect 570292 83098 570528 83334
rect 570612 83098 570848 83334
rect 585342 83418 585578 83654
rect 585662 83418 585898 83654
rect 585342 83098 585578 83334
rect 585662 83098 585898 83334
rect 7876 63418 8112 63654
rect 8196 63418 8432 63654
rect 7876 63098 8112 63334
rect 8196 63098 8432 63334
rect 38032 63418 38268 63654
rect 38352 63418 38588 63654
rect 38032 63098 38268 63334
rect 38352 63098 38588 63334
rect 60622 63418 60858 63654
rect 60622 63098 60858 63334
rect 159098 63418 159334 63654
rect 159098 63098 159334 63334
rect 182032 63418 182268 63654
rect 182352 63418 182588 63654
rect 182032 63098 182268 63334
rect 182352 63098 182588 63334
rect 185622 63418 185858 63654
rect 185622 63098 185858 63334
rect 284098 63418 284334 63654
rect 284098 63098 284334 63334
rect 290032 63418 290268 63654
rect 290352 63418 290588 63654
rect 290032 63098 290268 63334
rect 290352 63098 290588 63334
rect 310622 63418 310858 63654
rect 310622 63098 310858 63334
rect 409098 63418 409334 63654
rect 409098 63098 409334 63334
rect 434032 63418 434268 63654
rect 434352 63418 434588 63654
rect 434032 63098 434268 63334
rect 434352 63098 434588 63334
rect 436622 63418 436858 63654
rect 436622 63098 436858 63334
rect 535098 63418 535334 63654
rect 535098 63098 535334 63334
rect 542032 63418 542268 63654
rect 542352 63418 542588 63654
rect 542032 63098 542268 63334
rect 542352 63098 542588 63334
rect 571532 63418 571768 63654
rect 571852 63418 572088 63654
rect 571532 63098 571768 63334
rect 571852 63098 572088 63334
rect -1974 43418 -1738 43654
rect -1654 43418 -1418 43654
rect -1974 43098 -1738 43334
rect -1654 43098 -1418 43334
rect 9116 43418 9352 43654
rect 9436 43418 9672 43654
rect 9116 43098 9352 43334
rect 9436 43098 9672 43334
rect 56652 43418 56888 43654
rect 56972 43418 57208 43654
rect 56652 43098 56888 43334
rect 56972 43098 57208 43334
rect 61342 43418 61578 43654
rect 61342 43098 61578 43334
rect 158378 43418 158614 43654
rect 158378 43098 158614 43334
rect 164652 43418 164888 43654
rect 164972 43418 165208 43654
rect 164652 43098 164888 43334
rect 164972 43098 165208 43334
rect 186342 43418 186578 43654
rect 186342 43098 186578 43334
rect 283378 43418 283614 43654
rect 283378 43098 283614 43334
rect 308652 43418 308888 43654
rect 308972 43418 309208 43654
rect 308652 43098 308888 43334
rect 308972 43098 309208 43334
rect 311342 43418 311578 43654
rect 311342 43098 311578 43334
rect 408378 43418 408614 43654
rect 408378 43098 408614 43334
rect 416652 43418 416888 43654
rect 416972 43418 417208 43654
rect 416652 43098 416888 43334
rect 416972 43098 417208 43334
rect 437342 43418 437578 43654
rect 437342 43098 437578 43334
rect 534378 43418 534614 43654
rect 534378 43098 534614 43334
rect 560652 43418 560888 43654
rect 560972 43418 561208 43654
rect 560652 43098 560888 43334
rect 560972 43098 561208 43334
rect 570292 43418 570528 43654
rect 570612 43418 570848 43654
rect 570292 43098 570528 43334
rect 570612 43098 570848 43334
rect 585342 43418 585578 43654
rect 585662 43418 585898 43654
rect 585342 43098 585578 43334
rect 585662 43098 585898 43334
rect 7876 23418 8112 23654
rect 8196 23418 8432 23654
rect 7876 23098 8112 23334
rect 8196 23098 8432 23334
rect 38032 23418 38268 23654
rect 38352 23418 38588 23654
rect 38032 23098 38268 23334
rect 38352 23098 38588 23334
rect 60622 23418 60858 23654
rect 60622 23098 60858 23334
rect 159098 23418 159334 23654
rect 159098 23098 159334 23334
rect 182032 23418 182268 23654
rect 182352 23418 182588 23654
rect 182032 23098 182268 23334
rect 182352 23098 182588 23334
rect 185622 23418 185858 23654
rect 185622 23098 185858 23334
rect 284098 23418 284334 23654
rect 284098 23098 284334 23334
rect 290032 23418 290268 23654
rect 290352 23418 290588 23654
rect 290032 23098 290268 23334
rect 290352 23098 290588 23334
rect 310622 23418 310858 23654
rect 310622 23098 310858 23334
rect 409098 23418 409334 23654
rect 409098 23098 409334 23334
rect 434032 23418 434268 23654
rect 434352 23418 434588 23654
rect 434032 23098 434268 23334
rect 434352 23098 434588 23334
rect 436622 23418 436858 23654
rect 436622 23098 436858 23334
rect 535098 23418 535334 23654
rect 535098 23098 535334 23334
rect 542032 23418 542268 23654
rect 542352 23418 542588 23654
rect 542032 23098 542268 23334
rect 542352 23098 542588 23334
rect 571532 23418 571768 23654
rect 571852 23418 572088 23654
rect 571532 23098 571768 23334
rect 571852 23098 572088 23334
rect -1974 3418 -1738 3654
rect -1654 3418 -1418 3654
rect -1974 3098 -1738 3334
rect -1654 3098 -1418 3334
rect 585342 3418 585578 3654
rect 585662 3418 585898 3654
rect 585342 3098 585578 3334
rect 585662 3098 585898 3334
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 2026 -582 2262 -346
rect 2346 -582 2582 -346
rect 2026 -902 2262 -666
rect 2346 -902 2582 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5746 -2502 5982 -2266
rect 6066 -2502 6302 -2266
rect 5746 -2822 5982 -2586
rect 6066 -2822 6302 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9466 -4422 9702 -4186
rect 9786 -4422 10022 -4186
rect 9466 -4742 9702 -4506
rect 9786 -4742 10022 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 22026 -1542 22262 -1306
rect 22346 -1542 22582 -1306
rect 22026 -1862 22262 -1626
rect 22346 -1862 22582 -1626
rect 25746 -3462 25982 -3226
rect 26066 -3462 26302 -3226
rect 25746 -3782 25982 -3546
rect 26066 -3782 26302 -3546
rect 29466 -5382 29702 -5146
rect 29786 -5382 30022 -5146
rect 29466 -5702 29702 -5466
rect 29786 -5702 30022 -5466
rect 13186 -6342 13422 -6106
rect 13506 -6342 13742 -6106
rect 13186 -6662 13422 -6426
rect 13506 -6662 13742 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 42026 -582 42262 -346
rect 42346 -582 42582 -346
rect 42026 -902 42262 -666
rect 42346 -902 42582 -666
rect 45746 -2502 45982 -2266
rect 46066 -2502 46302 -2266
rect 45746 -2822 45982 -2586
rect 46066 -2822 46302 -2586
rect 49466 -4422 49702 -4186
rect 49786 -4422 50022 -4186
rect 49466 -4742 49702 -4506
rect 49786 -4742 50022 -4506
rect 33186 -7302 33422 -7066
rect 33506 -7302 33742 -7066
rect 33186 -7622 33422 -7386
rect 33506 -7622 33742 -7386
rect 62026 -1542 62262 -1306
rect 62346 -1542 62582 -1306
rect 62026 -1862 62262 -1626
rect 62346 -1862 62582 -1626
rect 65746 -3462 65982 -3226
rect 66066 -3462 66302 -3226
rect 65746 -3782 65982 -3546
rect 66066 -3782 66302 -3546
rect 69466 -5382 69702 -5146
rect 69786 -5382 70022 -5146
rect 69466 -5702 69702 -5466
rect 69786 -5702 70022 -5466
rect 53186 -6342 53422 -6106
rect 53506 -6342 53742 -6106
rect 53186 -6662 53422 -6426
rect 53506 -6662 53742 -6426
rect 82026 -582 82262 -346
rect 82346 -582 82582 -346
rect 82026 -902 82262 -666
rect 82346 -902 82582 -666
rect 85746 -2502 85982 -2266
rect 86066 -2502 86302 -2266
rect 85746 -2822 85982 -2586
rect 86066 -2822 86302 -2586
rect 89466 -4422 89702 -4186
rect 89786 -4422 90022 -4186
rect 89466 -4742 89702 -4506
rect 89786 -4742 90022 -4506
rect 73186 -7302 73422 -7066
rect 73506 -7302 73742 -7066
rect 73186 -7622 73422 -7386
rect 73506 -7622 73742 -7386
rect 102026 -1542 102262 -1306
rect 102346 -1542 102582 -1306
rect 102026 -1862 102262 -1626
rect 102346 -1862 102582 -1626
rect 105746 -3462 105982 -3226
rect 106066 -3462 106302 -3226
rect 105746 -3782 105982 -3546
rect 106066 -3782 106302 -3546
rect 109466 -5382 109702 -5146
rect 109786 -5382 110022 -5146
rect 109466 -5702 109702 -5466
rect 109786 -5702 110022 -5466
rect 93186 -6342 93422 -6106
rect 93506 -6342 93742 -6106
rect 93186 -6662 93422 -6426
rect 93506 -6662 93742 -6426
rect 122026 -582 122262 -346
rect 122346 -582 122582 -346
rect 122026 -902 122262 -666
rect 122346 -902 122582 -666
rect 125746 -2502 125982 -2266
rect 126066 -2502 126302 -2266
rect 125746 -2822 125982 -2586
rect 126066 -2822 126302 -2586
rect 129466 -4422 129702 -4186
rect 129786 -4422 130022 -4186
rect 129466 -4742 129702 -4506
rect 129786 -4742 130022 -4506
rect 113186 -7302 113422 -7066
rect 113506 -7302 113742 -7066
rect 113186 -7622 113422 -7386
rect 113506 -7622 113742 -7386
rect 142026 -1542 142262 -1306
rect 142346 -1542 142582 -1306
rect 142026 -1862 142262 -1626
rect 142346 -1862 142582 -1626
rect 145746 -3462 145982 -3226
rect 146066 -3462 146302 -3226
rect 145746 -3782 145982 -3546
rect 146066 -3782 146302 -3546
rect 149466 -5382 149702 -5146
rect 149786 -5382 150022 -5146
rect 149466 -5702 149702 -5466
rect 149786 -5702 150022 -5466
rect 133186 -6342 133422 -6106
rect 133506 -6342 133742 -6106
rect 133186 -6662 133422 -6426
rect 133506 -6662 133742 -6426
rect 162026 -582 162262 -346
rect 162346 -582 162582 -346
rect 162026 -902 162262 -666
rect 162346 -902 162582 -666
rect 165746 -2502 165982 -2266
rect 166066 -2502 166302 -2266
rect 165746 -2822 165982 -2586
rect 166066 -2822 166302 -2586
rect 169466 -4422 169702 -4186
rect 169786 -4422 170022 -4186
rect 169466 -4742 169702 -4506
rect 169786 -4742 170022 -4506
rect 153186 -7302 153422 -7066
rect 153506 -7302 153742 -7066
rect 153186 -7622 153422 -7386
rect 153506 -7622 153742 -7386
rect 182026 -1542 182262 -1306
rect 182346 -1542 182582 -1306
rect 182026 -1862 182262 -1626
rect 182346 -1862 182582 -1626
rect 185746 -3462 185982 -3226
rect 186066 -3462 186302 -3226
rect 185746 -3782 185982 -3546
rect 186066 -3782 186302 -3546
rect 189466 -5382 189702 -5146
rect 189786 -5382 190022 -5146
rect 189466 -5702 189702 -5466
rect 189786 -5702 190022 -5466
rect 173186 -6342 173422 -6106
rect 173506 -6342 173742 -6106
rect 173186 -6662 173422 -6426
rect 173506 -6662 173742 -6426
rect 202026 -582 202262 -346
rect 202346 -582 202582 -346
rect 202026 -902 202262 -666
rect 202346 -902 202582 -666
rect 205746 -2502 205982 -2266
rect 206066 -2502 206302 -2266
rect 205746 -2822 205982 -2586
rect 206066 -2822 206302 -2586
rect 209466 -4422 209702 -4186
rect 209786 -4422 210022 -4186
rect 209466 -4742 209702 -4506
rect 209786 -4742 210022 -4506
rect 193186 -7302 193422 -7066
rect 193506 -7302 193742 -7066
rect 193186 -7622 193422 -7386
rect 193506 -7622 193742 -7386
rect 222026 -1542 222262 -1306
rect 222346 -1542 222582 -1306
rect 222026 -1862 222262 -1626
rect 222346 -1862 222582 -1626
rect 225746 -3462 225982 -3226
rect 226066 -3462 226302 -3226
rect 225746 -3782 225982 -3546
rect 226066 -3782 226302 -3546
rect 229466 -5382 229702 -5146
rect 229786 -5382 230022 -5146
rect 229466 -5702 229702 -5466
rect 229786 -5702 230022 -5466
rect 213186 -6342 213422 -6106
rect 213506 -6342 213742 -6106
rect 213186 -6662 213422 -6426
rect 213506 -6662 213742 -6426
rect 242026 -582 242262 -346
rect 242346 -582 242582 -346
rect 242026 -902 242262 -666
rect 242346 -902 242582 -666
rect 245746 -2502 245982 -2266
rect 246066 -2502 246302 -2266
rect 245746 -2822 245982 -2586
rect 246066 -2822 246302 -2586
rect 249466 -4422 249702 -4186
rect 249786 -4422 250022 -4186
rect 249466 -4742 249702 -4506
rect 249786 -4742 250022 -4506
rect 233186 -7302 233422 -7066
rect 233506 -7302 233742 -7066
rect 233186 -7622 233422 -7386
rect 233506 -7622 233742 -7386
rect 262026 -1542 262262 -1306
rect 262346 -1542 262582 -1306
rect 262026 -1862 262262 -1626
rect 262346 -1862 262582 -1626
rect 265746 -3462 265982 -3226
rect 266066 -3462 266302 -3226
rect 265746 -3782 265982 -3546
rect 266066 -3782 266302 -3546
rect 269466 -5382 269702 -5146
rect 269786 -5382 270022 -5146
rect 269466 -5702 269702 -5466
rect 269786 -5702 270022 -5466
rect 253186 -6342 253422 -6106
rect 253506 -6342 253742 -6106
rect 253186 -6662 253422 -6426
rect 253506 -6662 253742 -6426
rect 282026 -582 282262 -346
rect 282346 -582 282582 -346
rect 282026 -902 282262 -666
rect 282346 -902 282582 -666
rect 285746 -2502 285982 -2266
rect 286066 -2502 286302 -2266
rect 285746 -2822 285982 -2586
rect 286066 -2822 286302 -2586
rect 289466 -4422 289702 -4186
rect 289786 -4422 290022 -4186
rect 289466 -4742 289702 -4506
rect 289786 -4742 290022 -4506
rect 273186 -7302 273422 -7066
rect 273506 -7302 273742 -7066
rect 273186 -7622 273422 -7386
rect 273506 -7622 273742 -7386
rect 302026 -1542 302262 -1306
rect 302346 -1542 302582 -1306
rect 302026 -1862 302262 -1626
rect 302346 -1862 302582 -1626
rect 305746 -3462 305982 -3226
rect 306066 -3462 306302 -3226
rect 305746 -3782 305982 -3546
rect 306066 -3782 306302 -3546
rect 309466 -5382 309702 -5146
rect 309786 -5382 310022 -5146
rect 309466 -5702 309702 -5466
rect 309786 -5702 310022 -5466
rect 293186 -6342 293422 -6106
rect 293506 -6342 293742 -6106
rect 293186 -6662 293422 -6426
rect 293506 -6662 293742 -6426
rect 322026 -582 322262 -346
rect 322346 -582 322582 -346
rect 322026 -902 322262 -666
rect 322346 -902 322582 -666
rect 325746 -2502 325982 -2266
rect 326066 -2502 326302 -2266
rect 325746 -2822 325982 -2586
rect 326066 -2822 326302 -2586
rect 329466 -4422 329702 -4186
rect 329786 -4422 330022 -4186
rect 329466 -4742 329702 -4506
rect 329786 -4742 330022 -4506
rect 313186 -7302 313422 -7066
rect 313506 -7302 313742 -7066
rect 313186 -7622 313422 -7386
rect 313506 -7622 313742 -7386
rect 342026 -1542 342262 -1306
rect 342346 -1542 342582 -1306
rect 342026 -1862 342262 -1626
rect 342346 -1862 342582 -1626
rect 345746 -3462 345982 -3226
rect 346066 -3462 346302 -3226
rect 345746 -3782 345982 -3546
rect 346066 -3782 346302 -3546
rect 349466 -5382 349702 -5146
rect 349786 -5382 350022 -5146
rect 349466 -5702 349702 -5466
rect 349786 -5702 350022 -5466
rect 333186 -6342 333422 -6106
rect 333506 -6342 333742 -6106
rect 333186 -6662 333422 -6426
rect 333506 -6662 333742 -6426
rect 362026 -582 362262 -346
rect 362346 -582 362582 -346
rect 362026 -902 362262 -666
rect 362346 -902 362582 -666
rect 365746 -2502 365982 -2266
rect 366066 -2502 366302 -2266
rect 365746 -2822 365982 -2586
rect 366066 -2822 366302 -2586
rect 369466 -4422 369702 -4186
rect 369786 -4422 370022 -4186
rect 369466 -4742 369702 -4506
rect 369786 -4742 370022 -4506
rect 353186 -7302 353422 -7066
rect 353506 -7302 353742 -7066
rect 353186 -7622 353422 -7386
rect 353506 -7622 353742 -7386
rect 382026 -1542 382262 -1306
rect 382346 -1542 382582 -1306
rect 382026 -1862 382262 -1626
rect 382346 -1862 382582 -1626
rect 385746 -3462 385982 -3226
rect 386066 -3462 386302 -3226
rect 385746 -3782 385982 -3546
rect 386066 -3782 386302 -3546
rect 389466 -5382 389702 -5146
rect 389786 -5382 390022 -5146
rect 389466 -5702 389702 -5466
rect 389786 -5702 390022 -5466
rect 373186 -6342 373422 -6106
rect 373506 -6342 373742 -6106
rect 373186 -6662 373422 -6426
rect 373506 -6662 373742 -6426
rect 402026 -582 402262 -346
rect 402346 -582 402582 -346
rect 402026 -902 402262 -666
rect 402346 -902 402582 -666
rect 405746 -2502 405982 -2266
rect 406066 -2502 406302 -2266
rect 405746 -2822 405982 -2586
rect 406066 -2822 406302 -2586
rect 409466 -4422 409702 -4186
rect 409786 -4422 410022 -4186
rect 409466 -4742 409702 -4506
rect 409786 -4742 410022 -4506
rect 393186 -7302 393422 -7066
rect 393506 -7302 393742 -7066
rect 393186 -7622 393422 -7386
rect 393506 -7622 393742 -7386
rect 422026 -1542 422262 -1306
rect 422346 -1542 422582 -1306
rect 422026 -1862 422262 -1626
rect 422346 -1862 422582 -1626
rect 425746 -3462 425982 -3226
rect 426066 -3462 426302 -3226
rect 425746 -3782 425982 -3546
rect 426066 -3782 426302 -3546
rect 429466 -5382 429702 -5146
rect 429786 -5382 430022 -5146
rect 429466 -5702 429702 -5466
rect 429786 -5702 430022 -5466
rect 413186 -6342 413422 -6106
rect 413506 -6342 413742 -6106
rect 413186 -6662 413422 -6426
rect 413506 -6662 413742 -6426
rect 442026 -582 442262 -346
rect 442346 -582 442582 -346
rect 442026 -902 442262 -666
rect 442346 -902 442582 -666
rect 445746 -2502 445982 -2266
rect 446066 -2502 446302 -2266
rect 445746 -2822 445982 -2586
rect 446066 -2822 446302 -2586
rect 449466 -4422 449702 -4186
rect 449786 -4422 450022 -4186
rect 449466 -4742 449702 -4506
rect 449786 -4742 450022 -4506
rect 433186 -7302 433422 -7066
rect 433506 -7302 433742 -7066
rect 433186 -7622 433422 -7386
rect 433506 -7622 433742 -7386
rect 462026 -1542 462262 -1306
rect 462346 -1542 462582 -1306
rect 462026 -1862 462262 -1626
rect 462346 -1862 462582 -1626
rect 465746 -3462 465982 -3226
rect 466066 -3462 466302 -3226
rect 465746 -3782 465982 -3546
rect 466066 -3782 466302 -3546
rect 469466 -5382 469702 -5146
rect 469786 -5382 470022 -5146
rect 469466 -5702 469702 -5466
rect 469786 -5702 470022 -5466
rect 453186 -6342 453422 -6106
rect 453506 -6342 453742 -6106
rect 453186 -6662 453422 -6426
rect 453506 -6662 453742 -6426
rect 482026 -582 482262 -346
rect 482346 -582 482582 -346
rect 482026 -902 482262 -666
rect 482346 -902 482582 -666
rect 485746 -2502 485982 -2266
rect 486066 -2502 486302 -2266
rect 485746 -2822 485982 -2586
rect 486066 -2822 486302 -2586
rect 489466 -4422 489702 -4186
rect 489786 -4422 490022 -4186
rect 489466 -4742 489702 -4506
rect 489786 -4742 490022 -4506
rect 473186 -7302 473422 -7066
rect 473506 -7302 473742 -7066
rect 473186 -7622 473422 -7386
rect 473506 -7622 473742 -7386
rect 502026 -1542 502262 -1306
rect 502346 -1542 502582 -1306
rect 502026 -1862 502262 -1626
rect 502346 -1862 502582 -1626
rect 505746 -3462 505982 -3226
rect 506066 -3462 506302 -3226
rect 505746 -3782 505982 -3546
rect 506066 -3782 506302 -3546
rect 509466 -5382 509702 -5146
rect 509786 -5382 510022 -5146
rect 509466 -5702 509702 -5466
rect 509786 -5702 510022 -5466
rect 493186 -6342 493422 -6106
rect 493506 -6342 493742 -6106
rect 493186 -6662 493422 -6426
rect 493506 -6662 493742 -6426
rect 522026 -582 522262 -346
rect 522346 -582 522582 -346
rect 522026 -902 522262 -666
rect 522346 -902 522582 -666
rect 525746 -2502 525982 -2266
rect 526066 -2502 526302 -2266
rect 525746 -2822 525982 -2586
rect 526066 -2822 526302 -2586
rect 529466 -4422 529702 -4186
rect 529786 -4422 530022 -4186
rect 529466 -4742 529702 -4506
rect 529786 -4742 530022 -4506
rect 513186 -7302 513422 -7066
rect 513506 -7302 513742 -7066
rect 513186 -7622 513422 -7386
rect 513506 -7622 513742 -7386
rect 542026 -1542 542262 -1306
rect 542346 -1542 542582 -1306
rect 542026 -1862 542262 -1626
rect 542346 -1862 542582 -1626
rect 545746 -3462 545982 -3226
rect 546066 -3462 546302 -3226
rect 545746 -3782 545982 -3546
rect 546066 -3782 546302 -3546
rect 549466 -5382 549702 -5146
rect 549786 -5382 550022 -5146
rect 549466 -5702 549702 -5466
rect 549786 -5702 550022 -5466
rect 533186 -6342 533422 -6106
rect 533506 -6342 533742 -6106
rect 533186 -6662 533422 -6426
rect 533506 -6662 533742 -6426
rect 562026 -582 562262 -346
rect 562346 -582 562582 -346
rect 562026 -902 562262 -666
rect 562346 -902 562582 -666
rect 565746 -2502 565982 -2266
rect 566066 -2502 566302 -2266
rect 565746 -2822 565982 -2586
rect 566066 -2822 566302 -2586
rect 569466 -4422 569702 -4186
rect 569786 -4422 570022 -4186
rect 569466 -4742 569702 -4506
rect 569786 -4742 570022 -4506
rect 553186 -7302 553422 -7066
rect 553506 -7302 553742 -7066
rect 553186 -7622 553422 -7386
rect 553506 -7622 553742 -7386
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 663418 586538 663654
rect 586622 663418 586858 663654
rect 586302 663098 586538 663334
rect 586622 663098 586858 663334
rect 586302 623418 586538 623654
rect 586622 623418 586858 623654
rect 586302 623098 586538 623334
rect 586622 623098 586858 623334
rect 586302 583418 586538 583654
rect 586622 583418 586858 583654
rect 586302 583098 586538 583334
rect 586622 583098 586858 583334
rect 586302 543418 586538 543654
rect 586622 543418 586858 543654
rect 586302 543098 586538 543334
rect 586622 543098 586858 543334
rect 586302 503418 586538 503654
rect 586622 503418 586858 503654
rect 586302 503098 586538 503334
rect 586622 503098 586858 503334
rect 586302 463418 586538 463654
rect 586622 463418 586858 463654
rect 586302 463098 586538 463334
rect 586622 463098 586858 463334
rect 586302 423418 586538 423654
rect 586622 423418 586858 423654
rect 586302 423098 586538 423334
rect 586622 423098 586858 423334
rect 586302 383418 586538 383654
rect 586622 383418 586858 383654
rect 586302 383098 586538 383334
rect 586622 383098 586858 383334
rect 586302 343418 586538 343654
rect 586622 343418 586858 343654
rect 586302 343098 586538 343334
rect 586622 343098 586858 343334
rect 586302 303418 586538 303654
rect 586622 303418 586858 303654
rect 586302 303098 586538 303334
rect 586622 303098 586858 303334
rect 586302 263418 586538 263654
rect 586622 263418 586858 263654
rect 586302 263098 586538 263334
rect 586622 263098 586858 263334
rect 586302 223418 586538 223654
rect 586622 223418 586858 223654
rect 586302 223098 586538 223334
rect 586622 223098 586858 223334
rect 586302 183418 586538 183654
rect 586622 183418 586858 183654
rect 586302 183098 586538 183334
rect 586622 183098 586858 183334
rect 586302 143418 586538 143654
rect 586622 143418 586858 143654
rect 586302 143098 586538 143334
rect 586622 143098 586858 143334
rect 586302 103418 586538 103654
rect 586622 103418 586858 103654
rect 586302 103098 586538 103334
rect 586622 103098 586858 103334
rect 586302 63418 586538 63654
rect 586622 63418 586858 63654
rect 586302 63098 586538 63334
rect 586622 63098 586858 63334
rect 586302 23418 586538 23654
rect 586622 23418 586858 23654
rect 586302 23098 586538 23334
rect 586622 23098 586858 23334
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 687138 587498 687374
rect 587582 687138 587818 687374
rect 587262 686818 587498 687054
rect 587582 686818 587818 687054
rect 587262 647138 587498 647374
rect 587582 647138 587818 647374
rect 587262 646818 587498 647054
rect 587582 646818 587818 647054
rect 587262 607138 587498 607374
rect 587582 607138 587818 607374
rect 587262 606818 587498 607054
rect 587582 606818 587818 607054
rect 587262 567138 587498 567374
rect 587582 567138 587818 567374
rect 587262 566818 587498 567054
rect 587582 566818 587818 567054
rect 587262 527138 587498 527374
rect 587582 527138 587818 527374
rect 587262 526818 587498 527054
rect 587582 526818 587818 527054
rect 587262 487138 587498 487374
rect 587582 487138 587818 487374
rect 587262 486818 587498 487054
rect 587582 486818 587818 487054
rect 587262 447138 587498 447374
rect 587582 447138 587818 447374
rect 587262 446818 587498 447054
rect 587582 446818 587818 447054
rect 587262 407138 587498 407374
rect 587582 407138 587818 407374
rect 587262 406818 587498 407054
rect 587582 406818 587818 407054
rect 587262 367138 587498 367374
rect 587582 367138 587818 367374
rect 587262 366818 587498 367054
rect 587582 366818 587818 367054
rect 587262 327138 587498 327374
rect 587582 327138 587818 327374
rect 587262 326818 587498 327054
rect 587582 326818 587818 327054
rect 587262 287138 587498 287374
rect 587582 287138 587818 287374
rect 587262 286818 587498 287054
rect 587582 286818 587818 287054
rect 587262 247138 587498 247374
rect 587582 247138 587818 247374
rect 587262 246818 587498 247054
rect 587582 246818 587818 247054
rect 587262 207138 587498 207374
rect 587582 207138 587818 207374
rect 587262 206818 587498 207054
rect 587582 206818 587818 207054
rect 587262 167138 587498 167374
rect 587582 167138 587818 167374
rect 587262 166818 587498 167054
rect 587582 166818 587818 167054
rect 587262 127138 587498 127374
rect 587582 127138 587818 127374
rect 587262 126818 587498 127054
rect 587582 126818 587818 127054
rect 587262 87138 587498 87374
rect 587582 87138 587818 87374
rect 587262 86818 587498 87054
rect 587582 86818 587818 87054
rect 587262 47138 587498 47374
rect 587582 47138 587818 47374
rect 587262 46818 587498 47054
rect 587582 46818 587818 47054
rect 587262 7138 587498 7374
rect 587582 7138 587818 7374
rect 587262 6818 587498 7054
rect 587582 6818 587818 7054
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 667138 588458 667374
rect 588542 667138 588778 667374
rect 588222 666818 588458 667054
rect 588542 666818 588778 667054
rect 588222 627138 588458 627374
rect 588542 627138 588778 627374
rect 588222 626818 588458 627054
rect 588542 626818 588778 627054
rect 588222 587138 588458 587374
rect 588542 587138 588778 587374
rect 588222 586818 588458 587054
rect 588542 586818 588778 587054
rect 588222 547138 588458 547374
rect 588542 547138 588778 547374
rect 588222 546818 588458 547054
rect 588542 546818 588778 547054
rect 588222 507138 588458 507374
rect 588542 507138 588778 507374
rect 588222 506818 588458 507054
rect 588542 506818 588778 507054
rect 588222 467138 588458 467374
rect 588542 467138 588778 467374
rect 588222 466818 588458 467054
rect 588542 466818 588778 467054
rect 588222 427138 588458 427374
rect 588542 427138 588778 427374
rect 588222 426818 588458 427054
rect 588542 426818 588778 427054
rect 588222 387138 588458 387374
rect 588542 387138 588778 387374
rect 588222 386818 588458 387054
rect 588542 386818 588778 387054
rect 588222 347138 588458 347374
rect 588542 347138 588778 347374
rect 588222 346818 588458 347054
rect 588542 346818 588778 347054
rect 588222 307138 588458 307374
rect 588542 307138 588778 307374
rect 588222 306818 588458 307054
rect 588542 306818 588778 307054
rect 588222 267138 588458 267374
rect 588542 267138 588778 267374
rect 588222 266818 588458 267054
rect 588542 266818 588778 267054
rect 588222 227138 588458 227374
rect 588542 227138 588778 227374
rect 588222 226818 588458 227054
rect 588542 226818 588778 227054
rect 588222 187138 588458 187374
rect 588542 187138 588778 187374
rect 588222 186818 588458 187054
rect 588542 186818 588778 187054
rect 588222 147138 588458 147374
rect 588542 147138 588778 147374
rect 588222 146818 588458 147054
rect 588542 146818 588778 147054
rect 588222 107138 588458 107374
rect 588542 107138 588778 107374
rect 588222 106818 588458 107054
rect 588542 106818 588778 107054
rect 588222 67138 588458 67374
rect 588542 67138 588778 67374
rect 588222 66818 588458 67054
rect 588542 66818 588778 67054
rect 588222 27138 588458 27374
rect 588542 27138 588778 27374
rect 588222 26818 588458 27054
rect 588542 26818 588778 27054
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 690858 589418 691094
rect 589502 690858 589738 691094
rect 589182 690538 589418 690774
rect 589502 690538 589738 690774
rect 589182 650858 589418 651094
rect 589502 650858 589738 651094
rect 589182 650538 589418 650774
rect 589502 650538 589738 650774
rect 589182 610858 589418 611094
rect 589502 610858 589738 611094
rect 589182 610538 589418 610774
rect 589502 610538 589738 610774
rect 589182 570858 589418 571094
rect 589502 570858 589738 571094
rect 589182 570538 589418 570774
rect 589502 570538 589738 570774
rect 589182 530858 589418 531094
rect 589502 530858 589738 531094
rect 589182 530538 589418 530774
rect 589502 530538 589738 530774
rect 589182 490858 589418 491094
rect 589502 490858 589738 491094
rect 589182 490538 589418 490774
rect 589502 490538 589738 490774
rect 589182 450858 589418 451094
rect 589502 450858 589738 451094
rect 589182 450538 589418 450774
rect 589502 450538 589738 450774
rect 589182 410858 589418 411094
rect 589502 410858 589738 411094
rect 589182 410538 589418 410774
rect 589502 410538 589738 410774
rect 589182 370858 589418 371094
rect 589502 370858 589738 371094
rect 589182 370538 589418 370774
rect 589502 370538 589738 370774
rect 589182 330858 589418 331094
rect 589502 330858 589738 331094
rect 589182 330538 589418 330774
rect 589502 330538 589738 330774
rect 589182 290858 589418 291094
rect 589502 290858 589738 291094
rect 589182 290538 589418 290774
rect 589502 290538 589738 290774
rect 589182 250858 589418 251094
rect 589502 250858 589738 251094
rect 589182 250538 589418 250774
rect 589502 250538 589738 250774
rect 589182 210858 589418 211094
rect 589502 210858 589738 211094
rect 589182 210538 589418 210774
rect 589502 210538 589738 210774
rect 589182 170858 589418 171094
rect 589502 170858 589738 171094
rect 589182 170538 589418 170774
rect 589502 170538 589738 170774
rect 589182 130858 589418 131094
rect 589502 130858 589738 131094
rect 589182 130538 589418 130774
rect 589502 130538 589738 130774
rect 589182 90858 589418 91094
rect 589502 90858 589738 91094
rect 589182 90538 589418 90774
rect 589502 90538 589738 90774
rect 589182 50858 589418 51094
rect 589502 50858 589738 51094
rect 589182 50538 589418 50774
rect 589502 50538 589738 50774
rect 589182 10858 589418 11094
rect 589502 10858 589738 11094
rect 589182 10538 589418 10774
rect 589502 10538 589738 10774
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 670858 590378 671094
rect 590462 670858 590698 671094
rect 590142 670538 590378 670774
rect 590462 670538 590698 670774
rect 590142 630858 590378 631094
rect 590462 630858 590698 631094
rect 590142 630538 590378 630774
rect 590462 630538 590698 630774
rect 590142 590858 590378 591094
rect 590462 590858 590698 591094
rect 590142 590538 590378 590774
rect 590462 590538 590698 590774
rect 590142 550858 590378 551094
rect 590462 550858 590698 551094
rect 590142 550538 590378 550774
rect 590462 550538 590698 550774
rect 590142 510858 590378 511094
rect 590462 510858 590698 511094
rect 590142 510538 590378 510774
rect 590462 510538 590698 510774
rect 590142 470858 590378 471094
rect 590462 470858 590698 471094
rect 590142 470538 590378 470774
rect 590462 470538 590698 470774
rect 590142 430858 590378 431094
rect 590462 430858 590698 431094
rect 590142 430538 590378 430774
rect 590462 430538 590698 430774
rect 590142 390858 590378 391094
rect 590462 390858 590698 391094
rect 590142 390538 590378 390774
rect 590462 390538 590698 390774
rect 590142 350858 590378 351094
rect 590462 350858 590698 351094
rect 590142 350538 590378 350774
rect 590462 350538 590698 350774
rect 590142 310858 590378 311094
rect 590462 310858 590698 311094
rect 590142 310538 590378 310774
rect 590462 310538 590698 310774
rect 590142 270858 590378 271094
rect 590462 270858 590698 271094
rect 590142 270538 590378 270774
rect 590462 270538 590698 270774
rect 590142 230858 590378 231094
rect 590462 230858 590698 231094
rect 590142 230538 590378 230774
rect 590462 230538 590698 230774
rect 590142 190858 590378 191094
rect 590462 190858 590698 191094
rect 590142 190538 590378 190774
rect 590462 190538 590698 190774
rect 590142 150858 590378 151094
rect 590462 150858 590698 151094
rect 590142 150538 590378 150774
rect 590462 150538 590698 150774
rect 590142 110858 590378 111094
rect 590462 110858 590698 111094
rect 590142 110538 590378 110774
rect 590462 110538 590698 110774
rect 590142 70858 590378 71094
rect 590462 70858 590698 71094
rect 590142 70538 590378 70774
rect 590462 70538 590698 70774
rect 590142 30858 590378 31094
rect 590462 30858 590698 31094
rect 590142 30538 590378 30774
rect 590462 30538 590698 30774
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 694578 591338 694814
rect 591422 694578 591658 694814
rect 591102 694258 591338 694494
rect 591422 694258 591658 694494
rect 591102 654578 591338 654814
rect 591422 654578 591658 654814
rect 591102 654258 591338 654494
rect 591422 654258 591658 654494
rect 591102 614578 591338 614814
rect 591422 614578 591658 614814
rect 591102 614258 591338 614494
rect 591422 614258 591658 614494
rect 591102 574578 591338 574814
rect 591422 574578 591658 574814
rect 591102 574258 591338 574494
rect 591422 574258 591658 574494
rect 591102 534578 591338 534814
rect 591422 534578 591658 534814
rect 591102 534258 591338 534494
rect 591422 534258 591658 534494
rect 591102 494578 591338 494814
rect 591422 494578 591658 494814
rect 591102 494258 591338 494494
rect 591422 494258 591658 494494
rect 591102 454578 591338 454814
rect 591422 454578 591658 454814
rect 591102 454258 591338 454494
rect 591422 454258 591658 454494
rect 591102 414578 591338 414814
rect 591422 414578 591658 414814
rect 591102 414258 591338 414494
rect 591422 414258 591658 414494
rect 591102 374578 591338 374814
rect 591422 374578 591658 374814
rect 591102 374258 591338 374494
rect 591422 374258 591658 374494
rect 591102 334578 591338 334814
rect 591422 334578 591658 334814
rect 591102 334258 591338 334494
rect 591422 334258 591658 334494
rect 591102 294578 591338 294814
rect 591422 294578 591658 294814
rect 591102 294258 591338 294494
rect 591422 294258 591658 294494
rect 591102 254578 591338 254814
rect 591422 254578 591658 254814
rect 591102 254258 591338 254494
rect 591422 254258 591658 254494
rect 591102 214578 591338 214814
rect 591422 214578 591658 214814
rect 591102 214258 591338 214494
rect 591422 214258 591658 214494
rect 591102 174578 591338 174814
rect 591422 174578 591658 174814
rect 591102 174258 591338 174494
rect 591422 174258 591658 174494
rect 591102 134578 591338 134814
rect 591422 134578 591658 134814
rect 591102 134258 591338 134494
rect 591422 134258 591658 134494
rect 591102 94578 591338 94814
rect 591422 94578 591658 94814
rect 591102 94258 591338 94494
rect 591422 94258 591658 94494
rect 591102 54578 591338 54814
rect 591422 54578 591658 54814
rect 591102 54258 591338 54494
rect 591422 54258 591658 54494
rect 591102 14578 591338 14814
rect 591422 14578 591658 14814
rect 591102 14258 591338 14494
rect 591422 14258 591658 14494
rect 573186 -6342 573422 -6106
rect 573506 -6342 573742 -6106
rect 573186 -6662 573422 -6426
rect 573506 -6662 573742 -6426
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 674578 592298 674814
rect 592382 674578 592618 674814
rect 592062 674258 592298 674494
rect 592382 674258 592618 674494
rect 592062 634578 592298 634814
rect 592382 634578 592618 634814
rect 592062 634258 592298 634494
rect 592382 634258 592618 634494
rect 592062 594578 592298 594814
rect 592382 594578 592618 594814
rect 592062 594258 592298 594494
rect 592382 594258 592618 594494
rect 592062 554578 592298 554814
rect 592382 554578 592618 554814
rect 592062 554258 592298 554494
rect 592382 554258 592618 554494
rect 592062 514578 592298 514814
rect 592382 514578 592618 514814
rect 592062 514258 592298 514494
rect 592382 514258 592618 514494
rect 592062 474578 592298 474814
rect 592382 474578 592618 474814
rect 592062 474258 592298 474494
rect 592382 474258 592618 474494
rect 592062 434578 592298 434814
rect 592382 434578 592618 434814
rect 592062 434258 592298 434494
rect 592382 434258 592618 434494
rect 592062 394578 592298 394814
rect 592382 394578 592618 394814
rect 592062 394258 592298 394494
rect 592382 394258 592618 394494
rect 592062 354578 592298 354814
rect 592382 354578 592618 354814
rect 592062 354258 592298 354494
rect 592382 354258 592618 354494
rect 592062 314578 592298 314814
rect 592382 314578 592618 314814
rect 592062 314258 592298 314494
rect 592382 314258 592618 314494
rect 592062 274578 592298 274814
rect 592382 274578 592618 274814
rect 592062 274258 592298 274494
rect 592382 274258 592618 274494
rect 592062 234578 592298 234814
rect 592382 234578 592618 234814
rect 592062 234258 592298 234494
rect 592382 234258 592618 234494
rect 592062 194578 592298 194814
rect 592382 194578 592618 194814
rect 592062 194258 592298 194494
rect 592382 194258 592618 194494
rect 592062 154578 592298 154814
rect 592382 154578 592618 154814
rect 592062 154258 592298 154494
rect 592382 154258 592618 154494
rect 592062 114578 592298 114814
rect 592382 114578 592618 114814
rect 592062 114258 592298 114494
rect 592382 114258 592618 114494
rect 592062 74578 592298 74814
rect 592382 74578 592618 74814
rect 592062 74258 592298 74494
rect 592382 74258 592618 74494
rect 592062 34578 592298 34814
rect 592382 34578 592618 34814
rect 592062 34258 592298 34494
rect 592382 34258 592618 34494
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33186 711558
rect 33422 711322 33506 711558
rect 33742 711322 73186 711558
rect 73422 711322 73506 711558
rect 73742 711322 113186 711558
rect 113422 711322 113506 711558
rect 113742 711322 153186 711558
rect 153422 711322 153506 711558
rect 153742 711322 193186 711558
rect 193422 711322 193506 711558
rect 193742 711322 233186 711558
rect 233422 711322 233506 711558
rect 233742 711322 273186 711558
rect 273422 711322 273506 711558
rect 273742 711322 313186 711558
rect 313422 711322 313506 711558
rect 313742 711322 353186 711558
rect 353422 711322 353506 711558
rect 353742 711322 393186 711558
rect 393422 711322 393506 711558
rect 393742 711322 433186 711558
rect 433422 711322 433506 711558
rect 433742 711322 473186 711558
rect 473422 711322 473506 711558
rect 473742 711322 513186 711558
rect 513422 711322 513506 711558
rect 513742 711322 553186 711558
rect 553422 711322 553506 711558
rect 553742 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33186 711238
rect 33422 711002 33506 711238
rect 33742 711002 73186 711238
rect 73422 711002 73506 711238
rect 73742 711002 113186 711238
rect 113422 711002 113506 711238
rect 113742 711002 153186 711238
rect 153422 711002 153506 711238
rect 153742 711002 193186 711238
rect 193422 711002 193506 711238
rect 193742 711002 233186 711238
rect 233422 711002 233506 711238
rect 233742 711002 273186 711238
rect 273422 711002 273506 711238
rect 273742 711002 313186 711238
rect 313422 711002 313506 711238
rect 313742 711002 353186 711238
rect 353422 711002 353506 711238
rect 353742 711002 393186 711238
rect 393422 711002 393506 711238
rect 393742 711002 433186 711238
rect 433422 711002 433506 711238
rect 433742 711002 473186 711238
rect 473422 711002 473506 711238
rect 473742 711002 513186 711238
rect 513422 711002 513506 711238
rect 513742 711002 553186 711238
rect 553422 711002 553506 711238
rect 553742 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 13186 710598
rect 13422 710362 13506 710598
rect 13742 710362 53186 710598
rect 53422 710362 53506 710598
rect 53742 710362 93186 710598
rect 93422 710362 93506 710598
rect 93742 710362 133186 710598
rect 133422 710362 133506 710598
rect 133742 710362 173186 710598
rect 173422 710362 173506 710598
rect 173742 710362 213186 710598
rect 213422 710362 213506 710598
rect 213742 710362 253186 710598
rect 253422 710362 253506 710598
rect 253742 710362 293186 710598
rect 293422 710362 293506 710598
rect 293742 710362 333186 710598
rect 333422 710362 333506 710598
rect 333742 710362 373186 710598
rect 373422 710362 373506 710598
rect 373742 710362 413186 710598
rect 413422 710362 413506 710598
rect 413742 710362 453186 710598
rect 453422 710362 453506 710598
rect 453742 710362 493186 710598
rect 493422 710362 493506 710598
rect 493742 710362 533186 710598
rect 533422 710362 533506 710598
rect 533742 710362 573186 710598
rect 573422 710362 573506 710598
rect 573742 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 13186 710278
rect 13422 710042 13506 710278
rect 13742 710042 53186 710278
rect 53422 710042 53506 710278
rect 53742 710042 93186 710278
rect 93422 710042 93506 710278
rect 93742 710042 133186 710278
rect 133422 710042 133506 710278
rect 133742 710042 173186 710278
rect 173422 710042 173506 710278
rect 173742 710042 213186 710278
rect 213422 710042 213506 710278
rect 213742 710042 253186 710278
rect 253422 710042 253506 710278
rect 253742 710042 293186 710278
rect 293422 710042 293506 710278
rect 293742 710042 333186 710278
rect 333422 710042 333506 710278
rect 333742 710042 373186 710278
rect 373422 710042 373506 710278
rect 373742 710042 413186 710278
rect 413422 710042 413506 710278
rect 413742 710042 453186 710278
rect 453422 710042 453506 710278
rect 453742 710042 493186 710278
rect 493422 710042 493506 710278
rect 493742 710042 533186 710278
rect 533422 710042 533506 710278
rect 533742 710042 573186 710278
rect 573422 710042 573506 710278
rect 573742 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 29466 709638
rect 29702 709402 29786 709638
rect 30022 709402 69466 709638
rect 69702 709402 69786 709638
rect 70022 709402 109466 709638
rect 109702 709402 109786 709638
rect 110022 709402 149466 709638
rect 149702 709402 149786 709638
rect 150022 709402 189466 709638
rect 189702 709402 189786 709638
rect 190022 709402 229466 709638
rect 229702 709402 229786 709638
rect 230022 709402 269466 709638
rect 269702 709402 269786 709638
rect 270022 709402 309466 709638
rect 309702 709402 309786 709638
rect 310022 709402 349466 709638
rect 349702 709402 349786 709638
rect 350022 709402 389466 709638
rect 389702 709402 389786 709638
rect 390022 709402 429466 709638
rect 429702 709402 429786 709638
rect 430022 709402 469466 709638
rect 469702 709402 469786 709638
rect 470022 709402 509466 709638
rect 509702 709402 509786 709638
rect 510022 709402 549466 709638
rect 549702 709402 549786 709638
rect 550022 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 29466 709318
rect 29702 709082 29786 709318
rect 30022 709082 69466 709318
rect 69702 709082 69786 709318
rect 70022 709082 109466 709318
rect 109702 709082 109786 709318
rect 110022 709082 149466 709318
rect 149702 709082 149786 709318
rect 150022 709082 189466 709318
rect 189702 709082 189786 709318
rect 190022 709082 229466 709318
rect 229702 709082 229786 709318
rect 230022 709082 269466 709318
rect 269702 709082 269786 709318
rect 270022 709082 309466 709318
rect 309702 709082 309786 709318
rect 310022 709082 349466 709318
rect 349702 709082 349786 709318
rect 350022 709082 389466 709318
rect 389702 709082 389786 709318
rect 390022 709082 429466 709318
rect 429702 709082 429786 709318
rect 430022 709082 469466 709318
rect 469702 709082 469786 709318
rect 470022 709082 509466 709318
rect 509702 709082 509786 709318
rect 510022 709082 549466 709318
rect 549702 709082 549786 709318
rect 550022 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9466 708678
rect 9702 708442 9786 708678
rect 10022 708442 49466 708678
rect 49702 708442 49786 708678
rect 50022 708442 89466 708678
rect 89702 708442 89786 708678
rect 90022 708442 129466 708678
rect 129702 708442 129786 708678
rect 130022 708442 169466 708678
rect 169702 708442 169786 708678
rect 170022 708442 209466 708678
rect 209702 708442 209786 708678
rect 210022 708442 249466 708678
rect 249702 708442 249786 708678
rect 250022 708442 289466 708678
rect 289702 708442 289786 708678
rect 290022 708442 329466 708678
rect 329702 708442 329786 708678
rect 330022 708442 369466 708678
rect 369702 708442 369786 708678
rect 370022 708442 409466 708678
rect 409702 708442 409786 708678
rect 410022 708442 449466 708678
rect 449702 708442 449786 708678
rect 450022 708442 489466 708678
rect 489702 708442 489786 708678
rect 490022 708442 529466 708678
rect 529702 708442 529786 708678
rect 530022 708442 569466 708678
rect 569702 708442 569786 708678
rect 570022 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9466 708358
rect 9702 708122 9786 708358
rect 10022 708122 49466 708358
rect 49702 708122 49786 708358
rect 50022 708122 89466 708358
rect 89702 708122 89786 708358
rect 90022 708122 129466 708358
rect 129702 708122 129786 708358
rect 130022 708122 169466 708358
rect 169702 708122 169786 708358
rect 170022 708122 209466 708358
rect 209702 708122 209786 708358
rect 210022 708122 249466 708358
rect 249702 708122 249786 708358
rect 250022 708122 289466 708358
rect 289702 708122 289786 708358
rect 290022 708122 329466 708358
rect 329702 708122 329786 708358
rect 330022 708122 369466 708358
rect 369702 708122 369786 708358
rect 370022 708122 409466 708358
rect 409702 708122 409786 708358
rect 410022 708122 449466 708358
rect 449702 708122 449786 708358
rect 450022 708122 489466 708358
rect 489702 708122 489786 708358
rect 490022 708122 529466 708358
rect 529702 708122 529786 708358
rect 530022 708122 569466 708358
rect 569702 708122 569786 708358
rect 570022 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 25746 707718
rect 25982 707482 26066 707718
rect 26302 707482 65746 707718
rect 65982 707482 66066 707718
rect 66302 707482 105746 707718
rect 105982 707482 106066 707718
rect 106302 707482 145746 707718
rect 145982 707482 146066 707718
rect 146302 707482 185746 707718
rect 185982 707482 186066 707718
rect 186302 707482 225746 707718
rect 225982 707482 226066 707718
rect 226302 707482 265746 707718
rect 265982 707482 266066 707718
rect 266302 707482 305746 707718
rect 305982 707482 306066 707718
rect 306302 707482 345746 707718
rect 345982 707482 346066 707718
rect 346302 707482 385746 707718
rect 385982 707482 386066 707718
rect 386302 707482 425746 707718
rect 425982 707482 426066 707718
rect 426302 707482 465746 707718
rect 465982 707482 466066 707718
rect 466302 707482 505746 707718
rect 505982 707482 506066 707718
rect 506302 707482 545746 707718
rect 545982 707482 546066 707718
rect 546302 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 25746 707398
rect 25982 707162 26066 707398
rect 26302 707162 65746 707398
rect 65982 707162 66066 707398
rect 66302 707162 105746 707398
rect 105982 707162 106066 707398
rect 106302 707162 145746 707398
rect 145982 707162 146066 707398
rect 146302 707162 185746 707398
rect 185982 707162 186066 707398
rect 186302 707162 225746 707398
rect 225982 707162 226066 707398
rect 226302 707162 265746 707398
rect 265982 707162 266066 707398
rect 266302 707162 305746 707398
rect 305982 707162 306066 707398
rect 306302 707162 345746 707398
rect 345982 707162 346066 707398
rect 346302 707162 385746 707398
rect 385982 707162 386066 707398
rect 386302 707162 425746 707398
rect 425982 707162 426066 707398
rect 426302 707162 465746 707398
rect 465982 707162 466066 707398
rect 466302 707162 505746 707398
rect 505982 707162 506066 707398
rect 506302 707162 545746 707398
rect 545982 707162 546066 707398
rect 546302 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5746 706758
rect 5982 706522 6066 706758
rect 6302 706522 45746 706758
rect 45982 706522 46066 706758
rect 46302 706522 85746 706758
rect 85982 706522 86066 706758
rect 86302 706522 125746 706758
rect 125982 706522 126066 706758
rect 126302 706522 165746 706758
rect 165982 706522 166066 706758
rect 166302 706522 205746 706758
rect 205982 706522 206066 706758
rect 206302 706522 245746 706758
rect 245982 706522 246066 706758
rect 246302 706522 285746 706758
rect 285982 706522 286066 706758
rect 286302 706522 325746 706758
rect 325982 706522 326066 706758
rect 326302 706522 365746 706758
rect 365982 706522 366066 706758
rect 366302 706522 405746 706758
rect 405982 706522 406066 706758
rect 406302 706522 445746 706758
rect 445982 706522 446066 706758
rect 446302 706522 485746 706758
rect 485982 706522 486066 706758
rect 486302 706522 525746 706758
rect 525982 706522 526066 706758
rect 526302 706522 565746 706758
rect 565982 706522 566066 706758
rect 566302 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5746 706438
rect 5982 706202 6066 706438
rect 6302 706202 45746 706438
rect 45982 706202 46066 706438
rect 46302 706202 85746 706438
rect 85982 706202 86066 706438
rect 86302 706202 125746 706438
rect 125982 706202 126066 706438
rect 126302 706202 165746 706438
rect 165982 706202 166066 706438
rect 166302 706202 205746 706438
rect 205982 706202 206066 706438
rect 206302 706202 245746 706438
rect 245982 706202 246066 706438
rect 246302 706202 285746 706438
rect 285982 706202 286066 706438
rect 286302 706202 325746 706438
rect 325982 706202 326066 706438
rect 326302 706202 365746 706438
rect 365982 706202 366066 706438
rect 366302 706202 405746 706438
rect 405982 706202 406066 706438
rect 406302 706202 445746 706438
rect 445982 706202 446066 706438
rect 446302 706202 485746 706438
rect 485982 706202 486066 706438
rect 486302 706202 525746 706438
rect 525982 706202 526066 706438
rect 526302 706202 565746 706438
rect 565982 706202 566066 706438
rect 566302 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 22026 705798
rect 22262 705562 22346 705798
rect 22582 705562 62026 705798
rect 62262 705562 62346 705798
rect 62582 705562 102026 705798
rect 102262 705562 102346 705798
rect 102582 705562 142026 705798
rect 142262 705562 142346 705798
rect 142582 705562 182026 705798
rect 182262 705562 182346 705798
rect 182582 705562 222026 705798
rect 222262 705562 222346 705798
rect 222582 705562 262026 705798
rect 262262 705562 262346 705798
rect 262582 705562 302026 705798
rect 302262 705562 302346 705798
rect 302582 705562 342026 705798
rect 342262 705562 342346 705798
rect 342582 705562 382026 705798
rect 382262 705562 382346 705798
rect 382582 705562 422026 705798
rect 422262 705562 422346 705798
rect 422582 705562 462026 705798
rect 462262 705562 462346 705798
rect 462582 705562 502026 705798
rect 502262 705562 502346 705798
rect 502582 705562 542026 705798
rect 542262 705562 542346 705798
rect 542582 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 22026 705478
rect 22262 705242 22346 705478
rect 22582 705242 62026 705478
rect 62262 705242 62346 705478
rect 62582 705242 102026 705478
rect 102262 705242 102346 705478
rect 102582 705242 142026 705478
rect 142262 705242 142346 705478
rect 142582 705242 182026 705478
rect 182262 705242 182346 705478
rect 182582 705242 222026 705478
rect 222262 705242 222346 705478
rect 222582 705242 262026 705478
rect 262262 705242 262346 705478
rect 262582 705242 302026 705478
rect 302262 705242 302346 705478
rect 302582 705242 342026 705478
rect 342262 705242 342346 705478
rect 342582 705242 382026 705478
rect 382262 705242 382346 705478
rect 382582 705242 422026 705478
rect 422262 705242 422346 705478
rect 422582 705242 462026 705478
rect 462262 705242 462346 705478
rect 462582 705242 502026 705478
rect 502262 705242 502346 705478
rect 502582 705242 542026 705478
rect 542262 705242 542346 705478
rect 542582 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 2026 704838
rect 2262 704602 2346 704838
rect 2582 704602 42026 704838
rect 42262 704602 42346 704838
rect 42582 704602 82026 704838
rect 82262 704602 82346 704838
rect 82582 704602 122026 704838
rect 122262 704602 122346 704838
rect 122582 704602 162026 704838
rect 162262 704602 162346 704838
rect 162582 704602 202026 704838
rect 202262 704602 202346 704838
rect 202582 704602 242026 704838
rect 242262 704602 242346 704838
rect 242582 704602 282026 704838
rect 282262 704602 282346 704838
rect 282582 704602 322026 704838
rect 322262 704602 322346 704838
rect 322582 704602 362026 704838
rect 362262 704602 362346 704838
rect 362582 704602 402026 704838
rect 402262 704602 402346 704838
rect 402582 704602 442026 704838
rect 442262 704602 442346 704838
rect 442582 704602 482026 704838
rect 482262 704602 482346 704838
rect 482582 704602 522026 704838
rect 522262 704602 522346 704838
rect 522582 704602 562026 704838
rect 562262 704602 562346 704838
rect 562582 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 2026 704518
rect 2262 704282 2346 704518
rect 2582 704282 42026 704518
rect 42262 704282 42346 704518
rect 42582 704282 82026 704518
rect 82262 704282 82346 704518
rect 82582 704282 122026 704518
rect 122262 704282 122346 704518
rect 122582 704282 162026 704518
rect 162262 704282 162346 704518
rect 162582 704282 202026 704518
rect 202262 704282 202346 704518
rect 202582 704282 242026 704518
rect 242262 704282 242346 704518
rect 242582 704282 282026 704518
rect 282262 704282 282346 704518
rect 282582 704282 322026 704518
rect 322262 704282 322346 704518
rect 322582 704282 362026 704518
rect 362262 704282 362346 704518
rect 362582 704282 402026 704518
rect 402262 704282 402346 704518
rect 402582 704282 442026 704518
rect 442262 704282 442346 704518
rect 442582 704282 482026 704518
rect 482262 704282 482346 704518
rect 482582 704282 522026 704518
rect 522262 704282 522346 704518
rect 522582 704282 562026 704518
rect 562262 704282 562346 704518
rect 562582 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 694814 592650 694846
rect -8726 694578 -7734 694814
rect -7498 694578 -7414 694814
rect -7178 694578 591102 694814
rect 591338 694578 591422 694814
rect 591658 694578 592650 694814
rect -8726 694494 592650 694578
rect -8726 694258 -7734 694494
rect -7498 694258 -7414 694494
rect -7178 694258 591102 694494
rect 591338 694258 591422 694494
rect 591658 694258 592650 694494
rect -8726 694226 592650 694258
rect -6806 691094 590730 691126
rect -6806 690858 -5814 691094
rect -5578 690858 -5494 691094
rect -5258 690858 589182 691094
rect 589418 690858 589502 691094
rect 589738 690858 590730 691094
rect -6806 690774 590730 690858
rect -6806 690538 -5814 690774
rect -5578 690538 -5494 690774
rect -5258 690538 589182 690774
rect 589418 690538 589502 690774
rect 589738 690538 590730 690774
rect -6806 690506 590730 690538
rect -4886 687374 588810 687406
rect -4886 687138 -3894 687374
rect -3658 687138 -3574 687374
rect -3338 687138 587262 687374
rect 587498 687138 587582 687374
rect 587818 687138 588810 687374
rect -4886 687054 588810 687138
rect -4886 686818 -3894 687054
rect -3658 686818 -3574 687054
rect -3338 686818 587262 687054
rect 587498 686818 587582 687054
rect 587818 686818 588810 687054
rect -4886 686786 588810 686818
rect -2966 683654 586890 683686
rect -2966 683418 -1974 683654
rect -1738 683418 -1654 683654
rect -1418 683418 9116 683654
rect 9352 683418 9436 683654
rect 9672 683418 56652 683654
rect 56888 683418 56972 683654
rect 57208 683418 92652 683654
rect 92888 683418 92972 683654
rect 93208 683418 128652 683654
rect 128888 683418 128972 683654
rect 129208 683418 164652 683654
rect 164888 683418 164972 683654
rect 165208 683418 200652 683654
rect 200888 683418 200972 683654
rect 201208 683418 236652 683654
rect 236888 683418 236972 683654
rect 237208 683418 272652 683654
rect 272888 683418 272972 683654
rect 273208 683418 308652 683654
rect 308888 683418 308972 683654
rect 309208 683418 344652 683654
rect 344888 683418 344972 683654
rect 345208 683418 380652 683654
rect 380888 683418 380972 683654
rect 381208 683418 416652 683654
rect 416888 683418 416972 683654
rect 417208 683418 452652 683654
rect 452888 683418 452972 683654
rect 453208 683418 488652 683654
rect 488888 683418 488972 683654
rect 489208 683418 524652 683654
rect 524888 683418 524972 683654
rect 525208 683418 560652 683654
rect 560888 683418 560972 683654
rect 561208 683418 570292 683654
rect 570528 683418 570612 683654
rect 570848 683418 585342 683654
rect 585578 683418 585662 683654
rect 585898 683418 586890 683654
rect -2966 683334 586890 683418
rect -2966 683098 -1974 683334
rect -1738 683098 -1654 683334
rect -1418 683098 9116 683334
rect 9352 683098 9436 683334
rect 9672 683098 56652 683334
rect 56888 683098 56972 683334
rect 57208 683098 92652 683334
rect 92888 683098 92972 683334
rect 93208 683098 128652 683334
rect 128888 683098 128972 683334
rect 129208 683098 164652 683334
rect 164888 683098 164972 683334
rect 165208 683098 200652 683334
rect 200888 683098 200972 683334
rect 201208 683098 236652 683334
rect 236888 683098 236972 683334
rect 237208 683098 272652 683334
rect 272888 683098 272972 683334
rect 273208 683098 308652 683334
rect 308888 683098 308972 683334
rect 309208 683098 344652 683334
rect 344888 683098 344972 683334
rect 345208 683098 380652 683334
rect 380888 683098 380972 683334
rect 381208 683098 416652 683334
rect 416888 683098 416972 683334
rect 417208 683098 452652 683334
rect 452888 683098 452972 683334
rect 453208 683098 488652 683334
rect 488888 683098 488972 683334
rect 489208 683098 524652 683334
rect 524888 683098 524972 683334
rect 525208 683098 560652 683334
rect 560888 683098 560972 683334
rect 561208 683098 570292 683334
rect 570528 683098 570612 683334
rect 570848 683098 585342 683334
rect 585578 683098 585662 683334
rect 585898 683098 586890 683334
rect -2966 683066 586890 683098
rect -8726 674814 592650 674846
rect -8726 674578 -8694 674814
rect -8458 674578 -8374 674814
rect -8138 674578 592062 674814
rect 592298 674578 592382 674814
rect 592618 674578 592650 674814
rect -8726 674494 592650 674578
rect -8726 674258 -8694 674494
rect -8458 674258 -8374 674494
rect -8138 674258 592062 674494
rect 592298 674258 592382 674494
rect 592618 674258 592650 674494
rect -8726 674226 592650 674258
rect -6806 671094 590730 671126
rect -6806 670858 -6774 671094
rect -6538 670858 -6454 671094
rect -6218 670858 590142 671094
rect 590378 670858 590462 671094
rect 590698 670858 590730 671094
rect -6806 670774 590730 670858
rect -6806 670538 -6774 670774
rect -6538 670538 -6454 670774
rect -6218 670538 590142 670774
rect 590378 670538 590462 670774
rect 590698 670538 590730 670774
rect -6806 670506 590730 670538
rect -4886 667374 588810 667406
rect -4886 667138 -4854 667374
rect -4618 667138 -4534 667374
rect -4298 667138 588222 667374
rect 588458 667138 588542 667374
rect 588778 667138 588810 667374
rect -4886 667054 588810 667138
rect -4886 666818 -4854 667054
rect -4618 666818 -4534 667054
rect -4298 666818 588222 667054
rect 588458 666818 588542 667054
rect 588778 666818 588810 667054
rect -4886 666786 588810 666818
rect -2966 663654 586890 663686
rect -2966 663418 -2934 663654
rect -2698 663418 -2614 663654
rect -2378 663418 7876 663654
rect 8112 663418 8196 663654
rect 8432 663418 38032 663654
rect 38268 663418 38352 663654
rect 38588 663418 74032 663654
rect 74268 663418 74352 663654
rect 74588 663418 110032 663654
rect 110268 663418 110352 663654
rect 110588 663418 146032 663654
rect 146268 663418 146352 663654
rect 146588 663418 182032 663654
rect 182268 663418 182352 663654
rect 182588 663418 218032 663654
rect 218268 663418 218352 663654
rect 218588 663418 254032 663654
rect 254268 663418 254352 663654
rect 254588 663418 290032 663654
rect 290268 663418 290352 663654
rect 290588 663418 326032 663654
rect 326268 663418 326352 663654
rect 326588 663418 362032 663654
rect 362268 663418 362352 663654
rect 362588 663418 398032 663654
rect 398268 663418 398352 663654
rect 398588 663418 434032 663654
rect 434268 663418 434352 663654
rect 434588 663418 470032 663654
rect 470268 663418 470352 663654
rect 470588 663418 506032 663654
rect 506268 663418 506352 663654
rect 506588 663418 542032 663654
rect 542268 663418 542352 663654
rect 542588 663418 571532 663654
rect 571768 663418 571852 663654
rect 572088 663418 586302 663654
rect 586538 663418 586622 663654
rect 586858 663418 586890 663654
rect -2966 663334 586890 663418
rect -2966 663098 -2934 663334
rect -2698 663098 -2614 663334
rect -2378 663098 7876 663334
rect 8112 663098 8196 663334
rect 8432 663098 38032 663334
rect 38268 663098 38352 663334
rect 38588 663098 74032 663334
rect 74268 663098 74352 663334
rect 74588 663098 110032 663334
rect 110268 663098 110352 663334
rect 110588 663098 146032 663334
rect 146268 663098 146352 663334
rect 146588 663098 182032 663334
rect 182268 663098 182352 663334
rect 182588 663098 218032 663334
rect 218268 663098 218352 663334
rect 218588 663098 254032 663334
rect 254268 663098 254352 663334
rect 254588 663098 290032 663334
rect 290268 663098 290352 663334
rect 290588 663098 326032 663334
rect 326268 663098 326352 663334
rect 326588 663098 362032 663334
rect 362268 663098 362352 663334
rect 362588 663098 398032 663334
rect 398268 663098 398352 663334
rect 398588 663098 434032 663334
rect 434268 663098 434352 663334
rect 434588 663098 470032 663334
rect 470268 663098 470352 663334
rect 470588 663098 506032 663334
rect 506268 663098 506352 663334
rect 506588 663098 542032 663334
rect 542268 663098 542352 663334
rect 542588 663098 571532 663334
rect 571768 663098 571852 663334
rect 572088 663098 586302 663334
rect 586538 663098 586622 663334
rect 586858 663098 586890 663334
rect -2966 663066 586890 663098
rect -8726 654814 592650 654846
rect -8726 654578 -7734 654814
rect -7498 654578 -7414 654814
rect -7178 654578 591102 654814
rect 591338 654578 591422 654814
rect 591658 654578 592650 654814
rect -8726 654494 592650 654578
rect -8726 654258 -7734 654494
rect -7498 654258 -7414 654494
rect -7178 654258 591102 654494
rect 591338 654258 591422 654494
rect 591658 654258 592650 654494
rect -8726 654226 592650 654258
rect -6806 651094 590730 651126
rect -6806 650858 -5814 651094
rect -5578 650858 -5494 651094
rect -5258 650858 589182 651094
rect 589418 650858 589502 651094
rect 589738 650858 590730 651094
rect -6806 650774 590730 650858
rect -6806 650538 -5814 650774
rect -5578 650538 -5494 650774
rect -5258 650538 589182 650774
rect 589418 650538 589502 650774
rect 589738 650538 590730 650774
rect -6806 650506 590730 650538
rect -4886 647374 588810 647406
rect -4886 647138 -3894 647374
rect -3658 647138 -3574 647374
rect -3338 647138 587262 647374
rect 587498 647138 587582 647374
rect 587818 647138 588810 647374
rect -4886 647054 588810 647138
rect -4886 646818 -3894 647054
rect -3658 646818 -3574 647054
rect -3338 646818 587262 647054
rect 587498 646818 587582 647054
rect 587818 646818 588810 647054
rect -4886 646786 588810 646818
rect -2966 643654 586890 643686
rect -2966 643418 -1974 643654
rect -1738 643418 -1654 643654
rect -1418 643418 9116 643654
rect 9352 643418 9436 643654
rect 9672 643418 56652 643654
rect 56888 643418 56972 643654
rect 57208 643418 92652 643654
rect 92888 643418 92972 643654
rect 93208 643418 128652 643654
rect 128888 643418 128972 643654
rect 129208 643418 164652 643654
rect 164888 643418 164972 643654
rect 165208 643418 200652 643654
rect 200888 643418 200972 643654
rect 201208 643418 236652 643654
rect 236888 643418 236972 643654
rect 237208 643418 272652 643654
rect 272888 643418 272972 643654
rect 273208 643418 308652 643654
rect 308888 643418 308972 643654
rect 309208 643418 344652 643654
rect 344888 643418 344972 643654
rect 345208 643418 380652 643654
rect 380888 643418 380972 643654
rect 381208 643418 416652 643654
rect 416888 643418 416972 643654
rect 417208 643418 452652 643654
rect 452888 643418 452972 643654
rect 453208 643418 488652 643654
rect 488888 643418 488972 643654
rect 489208 643418 524652 643654
rect 524888 643418 524972 643654
rect 525208 643418 560652 643654
rect 560888 643418 560972 643654
rect 561208 643418 570292 643654
rect 570528 643418 570612 643654
rect 570848 643418 585342 643654
rect 585578 643418 585662 643654
rect 585898 643418 586890 643654
rect -2966 643334 586890 643418
rect -2966 643098 -1974 643334
rect -1738 643098 -1654 643334
rect -1418 643098 9116 643334
rect 9352 643098 9436 643334
rect 9672 643098 56652 643334
rect 56888 643098 56972 643334
rect 57208 643098 92652 643334
rect 92888 643098 92972 643334
rect 93208 643098 128652 643334
rect 128888 643098 128972 643334
rect 129208 643098 164652 643334
rect 164888 643098 164972 643334
rect 165208 643098 200652 643334
rect 200888 643098 200972 643334
rect 201208 643098 236652 643334
rect 236888 643098 236972 643334
rect 237208 643098 272652 643334
rect 272888 643098 272972 643334
rect 273208 643098 308652 643334
rect 308888 643098 308972 643334
rect 309208 643098 344652 643334
rect 344888 643098 344972 643334
rect 345208 643098 380652 643334
rect 380888 643098 380972 643334
rect 381208 643098 416652 643334
rect 416888 643098 416972 643334
rect 417208 643098 452652 643334
rect 452888 643098 452972 643334
rect 453208 643098 488652 643334
rect 488888 643098 488972 643334
rect 489208 643098 524652 643334
rect 524888 643098 524972 643334
rect 525208 643098 560652 643334
rect 560888 643098 560972 643334
rect 561208 643098 570292 643334
rect 570528 643098 570612 643334
rect 570848 643098 585342 643334
rect 585578 643098 585662 643334
rect 585898 643098 586890 643334
rect -2966 643066 586890 643098
rect -8726 634814 592650 634846
rect -8726 634578 -8694 634814
rect -8458 634578 -8374 634814
rect -8138 634578 592062 634814
rect 592298 634578 592382 634814
rect 592618 634578 592650 634814
rect -8726 634494 592650 634578
rect -8726 634258 -8694 634494
rect -8458 634258 -8374 634494
rect -8138 634258 592062 634494
rect 592298 634258 592382 634494
rect 592618 634258 592650 634494
rect -8726 634226 592650 634258
rect -6806 631094 590730 631126
rect -6806 630858 -6774 631094
rect -6538 630858 -6454 631094
rect -6218 630858 590142 631094
rect 590378 630858 590462 631094
rect 590698 630858 590730 631094
rect -6806 630774 590730 630858
rect -6806 630538 -6774 630774
rect -6538 630538 -6454 630774
rect -6218 630538 590142 630774
rect 590378 630538 590462 630774
rect 590698 630538 590730 630774
rect -6806 630506 590730 630538
rect -4886 627374 588810 627406
rect -4886 627138 -4854 627374
rect -4618 627138 -4534 627374
rect -4298 627138 588222 627374
rect 588458 627138 588542 627374
rect 588778 627138 588810 627374
rect -4886 627054 588810 627138
rect -4886 626818 -4854 627054
rect -4618 626818 -4534 627054
rect -4298 626818 588222 627054
rect 588458 626818 588542 627054
rect 588778 626818 588810 627054
rect -4886 626786 588810 626818
rect -2966 623654 586890 623686
rect -2966 623418 -2934 623654
rect -2698 623418 -2614 623654
rect -2378 623418 7876 623654
rect 8112 623418 8196 623654
rect 8432 623418 38032 623654
rect 38268 623418 38352 623654
rect 38588 623418 74032 623654
rect 74268 623418 74352 623654
rect 74588 623418 110032 623654
rect 110268 623418 110352 623654
rect 110588 623418 146032 623654
rect 146268 623418 146352 623654
rect 146588 623418 182032 623654
rect 182268 623418 182352 623654
rect 182588 623418 218032 623654
rect 218268 623418 218352 623654
rect 218588 623418 254032 623654
rect 254268 623418 254352 623654
rect 254588 623418 290032 623654
rect 290268 623418 290352 623654
rect 290588 623418 326032 623654
rect 326268 623418 326352 623654
rect 326588 623418 362032 623654
rect 362268 623418 362352 623654
rect 362588 623418 398032 623654
rect 398268 623418 398352 623654
rect 398588 623418 434032 623654
rect 434268 623418 434352 623654
rect 434588 623418 470032 623654
rect 470268 623418 470352 623654
rect 470588 623418 506032 623654
rect 506268 623418 506352 623654
rect 506588 623418 542032 623654
rect 542268 623418 542352 623654
rect 542588 623418 571532 623654
rect 571768 623418 571852 623654
rect 572088 623418 586302 623654
rect 586538 623418 586622 623654
rect 586858 623418 586890 623654
rect -2966 623334 586890 623418
rect -2966 623098 -2934 623334
rect -2698 623098 -2614 623334
rect -2378 623098 7876 623334
rect 8112 623098 8196 623334
rect 8432 623098 38032 623334
rect 38268 623098 38352 623334
rect 38588 623098 74032 623334
rect 74268 623098 74352 623334
rect 74588 623098 110032 623334
rect 110268 623098 110352 623334
rect 110588 623098 146032 623334
rect 146268 623098 146352 623334
rect 146588 623098 182032 623334
rect 182268 623098 182352 623334
rect 182588 623098 218032 623334
rect 218268 623098 218352 623334
rect 218588 623098 254032 623334
rect 254268 623098 254352 623334
rect 254588 623098 290032 623334
rect 290268 623098 290352 623334
rect 290588 623098 326032 623334
rect 326268 623098 326352 623334
rect 326588 623098 362032 623334
rect 362268 623098 362352 623334
rect 362588 623098 398032 623334
rect 398268 623098 398352 623334
rect 398588 623098 434032 623334
rect 434268 623098 434352 623334
rect 434588 623098 470032 623334
rect 470268 623098 470352 623334
rect 470588 623098 506032 623334
rect 506268 623098 506352 623334
rect 506588 623098 542032 623334
rect 542268 623098 542352 623334
rect 542588 623098 571532 623334
rect 571768 623098 571852 623334
rect 572088 623098 586302 623334
rect 586538 623098 586622 623334
rect 586858 623098 586890 623334
rect -2966 623066 586890 623098
rect -8726 614814 592650 614846
rect -8726 614578 -7734 614814
rect -7498 614578 -7414 614814
rect -7178 614578 591102 614814
rect 591338 614578 591422 614814
rect 591658 614578 592650 614814
rect -8726 614494 592650 614578
rect -8726 614258 -7734 614494
rect -7498 614258 -7414 614494
rect -7178 614258 591102 614494
rect 591338 614258 591422 614494
rect 591658 614258 592650 614494
rect -8726 614226 592650 614258
rect -6806 611094 590730 611126
rect -6806 610858 -5814 611094
rect -5578 610858 -5494 611094
rect -5258 610858 589182 611094
rect 589418 610858 589502 611094
rect 589738 610858 590730 611094
rect -6806 610774 590730 610858
rect -6806 610538 -5814 610774
rect -5578 610538 -5494 610774
rect -5258 610538 589182 610774
rect 589418 610538 589502 610774
rect 589738 610538 590730 610774
rect -6806 610506 590730 610538
rect -4886 607374 588810 607406
rect -4886 607138 -3894 607374
rect -3658 607138 -3574 607374
rect -3338 607138 587262 607374
rect 587498 607138 587582 607374
rect 587818 607138 588810 607374
rect -4886 607054 588810 607138
rect -4886 606818 -3894 607054
rect -3658 606818 -3574 607054
rect -3338 606818 587262 607054
rect 587498 606818 587582 607054
rect 587818 606818 588810 607054
rect -4886 606786 588810 606818
rect -2966 603654 586890 603686
rect -2966 603418 -1974 603654
rect -1738 603418 -1654 603654
rect -1418 603418 9116 603654
rect 9352 603418 9436 603654
rect 9672 603418 56652 603654
rect 56888 603418 56972 603654
rect 57208 603418 92652 603654
rect 92888 603418 92972 603654
rect 93208 603418 128652 603654
rect 128888 603418 128972 603654
rect 129208 603418 164652 603654
rect 164888 603418 164972 603654
rect 165208 603418 200652 603654
rect 200888 603418 200972 603654
rect 201208 603418 236652 603654
rect 236888 603418 236972 603654
rect 237208 603418 272652 603654
rect 272888 603418 272972 603654
rect 273208 603418 308652 603654
rect 308888 603418 308972 603654
rect 309208 603418 344652 603654
rect 344888 603418 344972 603654
rect 345208 603418 380652 603654
rect 380888 603418 380972 603654
rect 381208 603418 416652 603654
rect 416888 603418 416972 603654
rect 417208 603418 452652 603654
rect 452888 603418 452972 603654
rect 453208 603418 488652 603654
rect 488888 603418 488972 603654
rect 489208 603418 524652 603654
rect 524888 603418 524972 603654
rect 525208 603418 560652 603654
rect 560888 603418 560972 603654
rect 561208 603418 570292 603654
rect 570528 603418 570612 603654
rect 570848 603418 585342 603654
rect 585578 603418 585662 603654
rect 585898 603418 586890 603654
rect -2966 603334 586890 603418
rect -2966 603098 -1974 603334
rect -1738 603098 -1654 603334
rect -1418 603098 9116 603334
rect 9352 603098 9436 603334
rect 9672 603098 56652 603334
rect 56888 603098 56972 603334
rect 57208 603098 92652 603334
rect 92888 603098 92972 603334
rect 93208 603098 128652 603334
rect 128888 603098 128972 603334
rect 129208 603098 164652 603334
rect 164888 603098 164972 603334
rect 165208 603098 200652 603334
rect 200888 603098 200972 603334
rect 201208 603098 236652 603334
rect 236888 603098 236972 603334
rect 237208 603098 272652 603334
rect 272888 603098 272972 603334
rect 273208 603098 308652 603334
rect 308888 603098 308972 603334
rect 309208 603098 344652 603334
rect 344888 603098 344972 603334
rect 345208 603098 380652 603334
rect 380888 603098 380972 603334
rect 381208 603098 416652 603334
rect 416888 603098 416972 603334
rect 417208 603098 452652 603334
rect 452888 603098 452972 603334
rect 453208 603098 488652 603334
rect 488888 603098 488972 603334
rect 489208 603098 524652 603334
rect 524888 603098 524972 603334
rect 525208 603098 560652 603334
rect 560888 603098 560972 603334
rect 561208 603098 570292 603334
rect 570528 603098 570612 603334
rect 570848 603098 585342 603334
rect 585578 603098 585662 603334
rect 585898 603098 586890 603334
rect -2966 603066 586890 603098
rect -8726 594814 592650 594846
rect -8726 594578 -8694 594814
rect -8458 594578 -8374 594814
rect -8138 594578 592062 594814
rect 592298 594578 592382 594814
rect 592618 594578 592650 594814
rect -8726 594494 592650 594578
rect -8726 594258 -8694 594494
rect -8458 594258 -8374 594494
rect -8138 594258 592062 594494
rect 592298 594258 592382 594494
rect 592618 594258 592650 594494
rect -8726 594226 592650 594258
rect -6806 591094 590730 591126
rect -6806 590858 -6774 591094
rect -6538 590858 -6454 591094
rect -6218 590858 590142 591094
rect 590378 590858 590462 591094
rect 590698 590858 590730 591094
rect -6806 590774 590730 590858
rect -6806 590538 -6774 590774
rect -6538 590538 -6454 590774
rect -6218 590538 590142 590774
rect 590378 590538 590462 590774
rect 590698 590538 590730 590774
rect -6806 590506 590730 590538
rect -4886 587374 588810 587406
rect -4886 587138 -4854 587374
rect -4618 587138 -4534 587374
rect -4298 587138 588222 587374
rect 588458 587138 588542 587374
rect 588778 587138 588810 587374
rect -4886 587054 588810 587138
rect -4886 586818 -4854 587054
rect -4618 586818 -4534 587054
rect -4298 586818 588222 587054
rect 588458 586818 588542 587054
rect 588778 586818 588810 587054
rect -4886 586786 588810 586818
rect -2966 583654 586890 583686
rect -2966 583418 -2934 583654
rect -2698 583418 -2614 583654
rect -2378 583418 7876 583654
rect 8112 583418 8196 583654
rect 8432 583418 38032 583654
rect 38268 583418 38352 583654
rect 38588 583418 74032 583654
rect 74268 583418 74352 583654
rect 74588 583418 110032 583654
rect 110268 583418 110352 583654
rect 110588 583418 146032 583654
rect 146268 583418 146352 583654
rect 146588 583418 182032 583654
rect 182268 583418 182352 583654
rect 182588 583418 218032 583654
rect 218268 583418 218352 583654
rect 218588 583418 254032 583654
rect 254268 583418 254352 583654
rect 254588 583418 290032 583654
rect 290268 583418 290352 583654
rect 290588 583418 326032 583654
rect 326268 583418 326352 583654
rect 326588 583418 362032 583654
rect 362268 583418 362352 583654
rect 362588 583418 398032 583654
rect 398268 583418 398352 583654
rect 398588 583418 434032 583654
rect 434268 583418 434352 583654
rect 434588 583418 470032 583654
rect 470268 583418 470352 583654
rect 470588 583418 506032 583654
rect 506268 583418 506352 583654
rect 506588 583418 542032 583654
rect 542268 583418 542352 583654
rect 542588 583418 571532 583654
rect 571768 583418 571852 583654
rect 572088 583418 586302 583654
rect 586538 583418 586622 583654
rect 586858 583418 586890 583654
rect -2966 583334 586890 583418
rect -2966 583098 -2934 583334
rect -2698 583098 -2614 583334
rect -2378 583098 7876 583334
rect 8112 583098 8196 583334
rect 8432 583098 38032 583334
rect 38268 583098 38352 583334
rect 38588 583098 74032 583334
rect 74268 583098 74352 583334
rect 74588 583098 110032 583334
rect 110268 583098 110352 583334
rect 110588 583098 146032 583334
rect 146268 583098 146352 583334
rect 146588 583098 182032 583334
rect 182268 583098 182352 583334
rect 182588 583098 218032 583334
rect 218268 583098 218352 583334
rect 218588 583098 254032 583334
rect 254268 583098 254352 583334
rect 254588 583098 290032 583334
rect 290268 583098 290352 583334
rect 290588 583098 326032 583334
rect 326268 583098 326352 583334
rect 326588 583098 362032 583334
rect 362268 583098 362352 583334
rect 362588 583098 398032 583334
rect 398268 583098 398352 583334
rect 398588 583098 434032 583334
rect 434268 583098 434352 583334
rect 434588 583098 470032 583334
rect 470268 583098 470352 583334
rect 470588 583098 506032 583334
rect 506268 583098 506352 583334
rect 506588 583098 542032 583334
rect 542268 583098 542352 583334
rect 542588 583098 571532 583334
rect 571768 583098 571852 583334
rect 572088 583098 586302 583334
rect 586538 583098 586622 583334
rect 586858 583098 586890 583334
rect -2966 583066 586890 583098
rect -8726 574814 592650 574846
rect -8726 574578 -7734 574814
rect -7498 574578 -7414 574814
rect -7178 574578 591102 574814
rect 591338 574578 591422 574814
rect 591658 574578 592650 574814
rect -8726 574494 592650 574578
rect -8726 574258 -7734 574494
rect -7498 574258 -7414 574494
rect -7178 574258 591102 574494
rect 591338 574258 591422 574494
rect 591658 574258 592650 574494
rect -8726 574226 592650 574258
rect -6806 571094 590730 571126
rect -6806 570858 -5814 571094
rect -5578 570858 -5494 571094
rect -5258 570858 589182 571094
rect 589418 570858 589502 571094
rect 589738 570858 590730 571094
rect -6806 570774 590730 570858
rect -6806 570538 -5814 570774
rect -5578 570538 -5494 570774
rect -5258 570538 589182 570774
rect 589418 570538 589502 570774
rect 589738 570538 590730 570774
rect -6806 570506 590730 570538
rect -4886 567374 588810 567406
rect -4886 567138 -3894 567374
rect -3658 567138 -3574 567374
rect -3338 567138 587262 567374
rect 587498 567138 587582 567374
rect 587818 567138 588810 567374
rect -4886 567054 588810 567138
rect -4886 566818 -3894 567054
rect -3658 566818 -3574 567054
rect -3338 566818 587262 567054
rect 587498 566818 587582 567054
rect 587818 566818 588810 567054
rect -4886 566786 588810 566818
rect -2966 563654 586890 563686
rect -2966 563418 -1974 563654
rect -1738 563418 -1654 563654
rect -1418 563418 9116 563654
rect 9352 563418 9436 563654
rect 9672 563418 56652 563654
rect 56888 563418 56972 563654
rect 57208 563418 92652 563654
rect 92888 563418 92972 563654
rect 93208 563418 128652 563654
rect 128888 563418 128972 563654
rect 129208 563418 164652 563654
rect 164888 563418 164972 563654
rect 165208 563418 200652 563654
rect 200888 563418 200972 563654
rect 201208 563418 236652 563654
rect 236888 563418 236972 563654
rect 237208 563418 272652 563654
rect 272888 563418 272972 563654
rect 273208 563418 308652 563654
rect 308888 563418 308972 563654
rect 309208 563418 344652 563654
rect 344888 563418 344972 563654
rect 345208 563418 380652 563654
rect 380888 563418 380972 563654
rect 381208 563418 416652 563654
rect 416888 563418 416972 563654
rect 417208 563418 452652 563654
rect 452888 563418 452972 563654
rect 453208 563418 488652 563654
rect 488888 563418 488972 563654
rect 489208 563418 524652 563654
rect 524888 563418 524972 563654
rect 525208 563418 560652 563654
rect 560888 563418 560972 563654
rect 561208 563418 570292 563654
rect 570528 563418 570612 563654
rect 570848 563418 585342 563654
rect 585578 563418 585662 563654
rect 585898 563418 586890 563654
rect -2966 563334 586890 563418
rect -2966 563098 -1974 563334
rect -1738 563098 -1654 563334
rect -1418 563098 9116 563334
rect 9352 563098 9436 563334
rect 9672 563098 56652 563334
rect 56888 563098 56972 563334
rect 57208 563098 92652 563334
rect 92888 563098 92972 563334
rect 93208 563098 128652 563334
rect 128888 563098 128972 563334
rect 129208 563098 164652 563334
rect 164888 563098 164972 563334
rect 165208 563098 200652 563334
rect 200888 563098 200972 563334
rect 201208 563098 236652 563334
rect 236888 563098 236972 563334
rect 237208 563098 272652 563334
rect 272888 563098 272972 563334
rect 273208 563098 308652 563334
rect 308888 563098 308972 563334
rect 309208 563098 344652 563334
rect 344888 563098 344972 563334
rect 345208 563098 380652 563334
rect 380888 563098 380972 563334
rect 381208 563098 416652 563334
rect 416888 563098 416972 563334
rect 417208 563098 452652 563334
rect 452888 563098 452972 563334
rect 453208 563098 488652 563334
rect 488888 563098 488972 563334
rect 489208 563098 524652 563334
rect 524888 563098 524972 563334
rect 525208 563098 560652 563334
rect 560888 563098 560972 563334
rect 561208 563098 570292 563334
rect 570528 563098 570612 563334
rect 570848 563098 585342 563334
rect 585578 563098 585662 563334
rect 585898 563098 586890 563334
rect -2966 563066 586890 563098
rect -8726 554814 592650 554846
rect -8726 554578 -8694 554814
rect -8458 554578 -8374 554814
rect -8138 554578 592062 554814
rect 592298 554578 592382 554814
rect 592618 554578 592650 554814
rect -8726 554494 592650 554578
rect -8726 554258 -8694 554494
rect -8458 554258 -8374 554494
rect -8138 554258 592062 554494
rect 592298 554258 592382 554494
rect 592618 554258 592650 554494
rect -8726 554226 592650 554258
rect -6806 551094 590730 551126
rect -6806 550858 -6774 551094
rect -6538 550858 -6454 551094
rect -6218 550858 590142 551094
rect 590378 550858 590462 551094
rect 590698 550858 590730 551094
rect -6806 550774 590730 550858
rect -6806 550538 -6774 550774
rect -6538 550538 -6454 550774
rect -6218 550538 590142 550774
rect 590378 550538 590462 550774
rect 590698 550538 590730 550774
rect -6806 550506 590730 550538
rect -4886 547374 588810 547406
rect -4886 547138 -4854 547374
rect -4618 547138 -4534 547374
rect -4298 547138 588222 547374
rect 588458 547138 588542 547374
rect 588778 547138 588810 547374
rect -4886 547054 588810 547138
rect -4886 546818 -4854 547054
rect -4618 546818 -4534 547054
rect -4298 546818 588222 547054
rect 588458 546818 588542 547054
rect 588778 546818 588810 547054
rect -4886 546786 588810 546818
rect -2966 543654 586890 543686
rect -2966 543418 -2934 543654
rect -2698 543418 -2614 543654
rect -2378 543418 7876 543654
rect 8112 543418 8196 543654
rect 8432 543418 38032 543654
rect 38268 543418 38352 543654
rect 38588 543418 74032 543654
rect 74268 543418 74352 543654
rect 74588 543418 110032 543654
rect 110268 543418 110352 543654
rect 110588 543418 146032 543654
rect 146268 543418 146352 543654
rect 146588 543418 182032 543654
rect 182268 543418 182352 543654
rect 182588 543418 218032 543654
rect 218268 543418 218352 543654
rect 218588 543418 254032 543654
rect 254268 543418 254352 543654
rect 254588 543418 290032 543654
rect 290268 543418 290352 543654
rect 290588 543418 326032 543654
rect 326268 543418 326352 543654
rect 326588 543418 362032 543654
rect 362268 543418 362352 543654
rect 362588 543418 398032 543654
rect 398268 543418 398352 543654
rect 398588 543418 434032 543654
rect 434268 543418 434352 543654
rect 434588 543418 470032 543654
rect 470268 543418 470352 543654
rect 470588 543418 506032 543654
rect 506268 543418 506352 543654
rect 506588 543418 542032 543654
rect 542268 543418 542352 543654
rect 542588 543418 571532 543654
rect 571768 543418 571852 543654
rect 572088 543418 586302 543654
rect 586538 543418 586622 543654
rect 586858 543418 586890 543654
rect -2966 543334 586890 543418
rect -2966 543098 -2934 543334
rect -2698 543098 -2614 543334
rect -2378 543098 7876 543334
rect 8112 543098 8196 543334
rect 8432 543098 38032 543334
rect 38268 543098 38352 543334
rect 38588 543098 74032 543334
rect 74268 543098 74352 543334
rect 74588 543098 110032 543334
rect 110268 543098 110352 543334
rect 110588 543098 146032 543334
rect 146268 543098 146352 543334
rect 146588 543098 182032 543334
rect 182268 543098 182352 543334
rect 182588 543098 218032 543334
rect 218268 543098 218352 543334
rect 218588 543098 254032 543334
rect 254268 543098 254352 543334
rect 254588 543098 290032 543334
rect 290268 543098 290352 543334
rect 290588 543098 326032 543334
rect 326268 543098 326352 543334
rect 326588 543098 362032 543334
rect 362268 543098 362352 543334
rect 362588 543098 398032 543334
rect 398268 543098 398352 543334
rect 398588 543098 434032 543334
rect 434268 543098 434352 543334
rect 434588 543098 470032 543334
rect 470268 543098 470352 543334
rect 470588 543098 506032 543334
rect 506268 543098 506352 543334
rect 506588 543098 542032 543334
rect 542268 543098 542352 543334
rect 542588 543098 571532 543334
rect 571768 543098 571852 543334
rect 572088 543098 586302 543334
rect 586538 543098 586622 543334
rect 586858 543098 586890 543334
rect -2966 543066 586890 543098
rect -8726 534814 592650 534846
rect -8726 534578 -7734 534814
rect -7498 534578 -7414 534814
rect -7178 534578 591102 534814
rect 591338 534578 591422 534814
rect 591658 534578 592650 534814
rect -8726 534494 592650 534578
rect -8726 534258 -7734 534494
rect -7498 534258 -7414 534494
rect -7178 534258 591102 534494
rect 591338 534258 591422 534494
rect 591658 534258 592650 534494
rect -8726 534226 592650 534258
rect -6806 531094 590730 531126
rect -6806 530858 -5814 531094
rect -5578 530858 -5494 531094
rect -5258 530858 589182 531094
rect 589418 530858 589502 531094
rect 589738 530858 590730 531094
rect -6806 530774 590730 530858
rect -6806 530538 -5814 530774
rect -5578 530538 -5494 530774
rect -5258 530538 589182 530774
rect 589418 530538 589502 530774
rect 589738 530538 590730 530774
rect -6806 530506 590730 530538
rect -4886 527374 588810 527406
rect -4886 527138 -3894 527374
rect -3658 527138 -3574 527374
rect -3338 527138 587262 527374
rect 587498 527138 587582 527374
rect 587818 527138 588810 527374
rect -4886 527054 588810 527138
rect -4886 526818 -3894 527054
rect -3658 526818 -3574 527054
rect -3338 526818 587262 527054
rect 587498 526818 587582 527054
rect 587818 526818 588810 527054
rect -4886 526786 588810 526818
rect -2966 523654 586890 523686
rect -2966 523418 -1974 523654
rect -1738 523418 -1654 523654
rect -1418 523418 9116 523654
rect 9352 523418 9436 523654
rect 9672 523418 56652 523654
rect 56888 523418 56972 523654
rect 57208 523418 92652 523654
rect 92888 523418 92972 523654
rect 93208 523418 128652 523654
rect 128888 523418 128972 523654
rect 129208 523418 164652 523654
rect 164888 523418 164972 523654
rect 165208 523418 200652 523654
rect 200888 523418 200972 523654
rect 201208 523418 236652 523654
rect 236888 523418 236972 523654
rect 237208 523418 272652 523654
rect 272888 523418 272972 523654
rect 273208 523418 308652 523654
rect 308888 523418 308972 523654
rect 309208 523418 344652 523654
rect 344888 523418 344972 523654
rect 345208 523418 380652 523654
rect 380888 523418 380972 523654
rect 381208 523418 416652 523654
rect 416888 523418 416972 523654
rect 417208 523418 452652 523654
rect 452888 523418 452972 523654
rect 453208 523418 488652 523654
rect 488888 523418 488972 523654
rect 489208 523418 524652 523654
rect 524888 523418 524972 523654
rect 525208 523418 560652 523654
rect 560888 523418 560972 523654
rect 561208 523418 570292 523654
rect 570528 523418 570612 523654
rect 570848 523418 585342 523654
rect 585578 523418 585662 523654
rect 585898 523418 586890 523654
rect -2966 523334 586890 523418
rect -2966 523098 -1974 523334
rect -1738 523098 -1654 523334
rect -1418 523098 9116 523334
rect 9352 523098 9436 523334
rect 9672 523098 56652 523334
rect 56888 523098 56972 523334
rect 57208 523098 92652 523334
rect 92888 523098 92972 523334
rect 93208 523098 128652 523334
rect 128888 523098 128972 523334
rect 129208 523098 164652 523334
rect 164888 523098 164972 523334
rect 165208 523098 200652 523334
rect 200888 523098 200972 523334
rect 201208 523098 236652 523334
rect 236888 523098 236972 523334
rect 237208 523098 272652 523334
rect 272888 523098 272972 523334
rect 273208 523098 308652 523334
rect 308888 523098 308972 523334
rect 309208 523098 344652 523334
rect 344888 523098 344972 523334
rect 345208 523098 380652 523334
rect 380888 523098 380972 523334
rect 381208 523098 416652 523334
rect 416888 523098 416972 523334
rect 417208 523098 452652 523334
rect 452888 523098 452972 523334
rect 453208 523098 488652 523334
rect 488888 523098 488972 523334
rect 489208 523098 524652 523334
rect 524888 523098 524972 523334
rect 525208 523098 560652 523334
rect 560888 523098 560972 523334
rect 561208 523098 570292 523334
rect 570528 523098 570612 523334
rect 570848 523098 585342 523334
rect 585578 523098 585662 523334
rect 585898 523098 586890 523334
rect -2966 523066 586890 523098
rect -8726 514814 592650 514846
rect -8726 514578 -8694 514814
rect -8458 514578 -8374 514814
rect -8138 514578 592062 514814
rect 592298 514578 592382 514814
rect 592618 514578 592650 514814
rect -8726 514494 592650 514578
rect -8726 514258 -8694 514494
rect -8458 514258 -8374 514494
rect -8138 514258 592062 514494
rect 592298 514258 592382 514494
rect 592618 514258 592650 514494
rect -8726 514226 592650 514258
rect -6806 511094 590730 511126
rect -6806 510858 -6774 511094
rect -6538 510858 -6454 511094
rect -6218 510858 590142 511094
rect 590378 510858 590462 511094
rect 590698 510858 590730 511094
rect -6806 510774 590730 510858
rect -6806 510538 -6774 510774
rect -6538 510538 -6454 510774
rect -6218 510538 590142 510774
rect 590378 510538 590462 510774
rect 590698 510538 590730 510774
rect -6806 510506 590730 510538
rect -4886 507374 588810 507406
rect -4886 507138 -4854 507374
rect -4618 507138 -4534 507374
rect -4298 507138 588222 507374
rect 588458 507138 588542 507374
rect 588778 507138 588810 507374
rect -4886 507054 588810 507138
rect -4886 506818 -4854 507054
rect -4618 506818 -4534 507054
rect -4298 506818 588222 507054
rect 588458 506818 588542 507054
rect 588778 506818 588810 507054
rect -4886 506786 588810 506818
rect -2966 503654 586890 503686
rect -2966 503418 -2934 503654
rect -2698 503418 -2614 503654
rect -2378 503418 7876 503654
rect 8112 503418 8196 503654
rect 8432 503418 38032 503654
rect 38268 503418 38352 503654
rect 38588 503418 60622 503654
rect 60858 503418 159098 503654
rect 159334 503418 182032 503654
rect 182268 503418 182352 503654
rect 182588 503418 185622 503654
rect 185858 503418 284098 503654
rect 284334 503418 290032 503654
rect 290268 503418 290352 503654
rect 290588 503418 310622 503654
rect 310858 503418 409098 503654
rect 409334 503418 434032 503654
rect 434268 503418 434352 503654
rect 434588 503418 436622 503654
rect 436858 503418 535098 503654
rect 535334 503418 542032 503654
rect 542268 503418 542352 503654
rect 542588 503418 571532 503654
rect 571768 503418 571852 503654
rect 572088 503418 586302 503654
rect 586538 503418 586622 503654
rect 586858 503418 586890 503654
rect -2966 503334 586890 503418
rect -2966 503098 -2934 503334
rect -2698 503098 -2614 503334
rect -2378 503098 7876 503334
rect 8112 503098 8196 503334
rect 8432 503098 38032 503334
rect 38268 503098 38352 503334
rect 38588 503098 60622 503334
rect 60858 503098 159098 503334
rect 159334 503098 182032 503334
rect 182268 503098 182352 503334
rect 182588 503098 185622 503334
rect 185858 503098 284098 503334
rect 284334 503098 290032 503334
rect 290268 503098 290352 503334
rect 290588 503098 310622 503334
rect 310858 503098 409098 503334
rect 409334 503098 434032 503334
rect 434268 503098 434352 503334
rect 434588 503098 436622 503334
rect 436858 503098 535098 503334
rect 535334 503098 542032 503334
rect 542268 503098 542352 503334
rect 542588 503098 571532 503334
rect 571768 503098 571852 503334
rect 572088 503098 586302 503334
rect 586538 503098 586622 503334
rect 586858 503098 586890 503334
rect -2966 503066 586890 503098
rect -8726 494814 592650 494846
rect -8726 494578 -7734 494814
rect -7498 494578 -7414 494814
rect -7178 494578 591102 494814
rect 591338 494578 591422 494814
rect 591658 494578 592650 494814
rect -8726 494494 592650 494578
rect -8726 494258 -7734 494494
rect -7498 494258 -7414 494494
rect -7178 494258 591102 494494
rect 591338 494258 591422 494494
rect 591658 494258 592650 494494
rect -8726 494226 592650 494258
rect -6806 491094 590730 491126
rect -6806 490858 -5814 491094
rect -5578 490858 -5494 491094
rect -5258 490858 589182 491094
rect 589418 490858 589502 491094
rect 589738 490858 590730 491094
rect -6806 490774 590730 490858
rect -6806 490538 -5814 490774
rect -5578 490538 -5494 490774
rect -5258 490538 589182 490774
rect 589418 490538 589502 490774
rect 589738 490538 590730 490774
rect -6806 490506 590730 490538
rect -4886 487374 588810 487406
rect -4886 487138 -3894 487374
rect -3658 487138 -3574 487374
rect -3338 487138 587262 487374
rect 587498 487138 587582 487374
rect 587818 487138 588810 487374
rect -4886 487054 588810 487138
rect -4886 486818 -3894 487054
rect -3658 486818 -3574 487054
rect -3338 486818 587262 487054
rect 587498 486818 587582 487054
rect 587818 486818 588810 487054
rect -4886 486786 588810 486818
rect -2966 483654 586890 483686
rect -2966 483418 -1974 483654
rect -1738 483418 -1654 483654
rect -1418 483418 9116 483654
rect 9352 483418 9436 483654
rect 9672 483418 56652 483654
rect 56888 483418 56972 483654
rect 57208 483418 61342 483654
rect 61578 483418 158378 483654
rect 158614 483418 164652 483654
rect 164888 483418 164972 483654
rect 165208 483418 186342 483654
rect 186578 483418 283378 483654
rect 283614 483418 308652 483654
rect 308888 483418 308972 483654
rect 309208 483418 311342 483654
rect 311578 483418 408378 483654
rect 408614 483418 416652 483654
rect 416888 483418 416972 483654
rect 417208 483418 437342 483654
rect 437578 483418 534378 483654
rect 534614 483418 560652 483654
rect 560888 483418 560972 483654
rect 561208 483418 570292 483654
rect 570528 483418 570612 483654
rect 570848 483418 585342 483654
rect 585578 483418 585662 483654
rect 585898 483418 586890 483654
rect -2966 483334 586890 483418
rect -2966 483098 -1974 483334
rect -1738 483098 -1654 483334
rect -1418 483098 9116 483334
rect 9352 483098 9436 483334
rect 9672 483098 56652 483334
rect 56888 483098 56972 483334
rect 57208 483098 61342 483334
rect 61578 483098 158378 483334
rect 158614 483098 164652 483334
rect 164888 483098 164972 483334
rect 165208 483098 186342 483334
rect 186578 483098 283378 483334
rect 283614 483098 308652 483334
rect 308888 483098 308972 483334
rect 309208 483098 311342 483334
rect 311578 483098 408378 483334
rect 408614 483098 416652 483334
rect 416888 483098 416972 483334
rect 417208 483098 437342 483334
rect 437578 483098 534378 483334
rect 534614 483098 560652 483334
rect 560888 483098 560972 483334
rect 561208 483098 570292 483334
rect 570528 483098 570612 483334
rect 570848 483098 585342 483334
rect 585578 483098 585662 483334
rect 585898 483098 586890 483334
rect -2966 483066 586890 483098
rect -8726 474814 592650 474846
rect -8726 474578 -8694 474814
rect -8458 474578 -8374 474814
rect -8138 474578 592062 474814
rect 592298 474578 592382 474814
rect 592618 474578 592650 474814
rect -8726 474494 592650 474578
rect -8726 474258 -8694 474494
rect -8458 474258 -8374 474494
rect -8138 474258 592062 474494
rect 592298 474258 592382 474494
rect 592618 474258 592650 474494
rect -8726 474226 592650 474258
rect -6806 471094 590730 471126
rect -6806 470858 -6774 471094
rect -6538 470858 -6454 471094
rect -6218 470858 590142 471094
rect 590378 470858 590462 471094
rect 590698 470858 590730 471094
rect -6806 470774 590730 470858
rect -6806 470538 -6774 470774
rect -6538 470538 -6454 470774
rect -6218 470538 590142 470774
rect 590378 470538 590462 470774
rect 590698 470538 590730 470774
rect -6806 470506 590730 470538
rect -4886 467374 588810 467406
rect -4886 467138 -4854 467374
rect -4618 467138 -4534 467374
rect -4298 467138 588222 467374
rect 588458 467138 588542 467374
rect 588778 467138 588810 467374
rect -4886 467054 588810 467138
rect -4886 466818 -4854 467054
rect -4618 466818 -4534 467054
rect -4298 466818 588222 467054
rect 588458 466818 588542 467054
rect 588778 466818 588810 467054
rect -4886 466786 588810 466818
rect -2966 463654 586890 463686
rect -2966 463418 -2934 463654
rect -2698 463418 -2614 463654
rect -2378 463418 7876 463654
rect 8112 463418 8196 463654
rect 8432 463418 38032 463654
rect 38268 463418 38352 463654
rect 38588 463418 60622 463654
rect 60858 463418 159098 463654
rect 159334 463418 182032 463654
rect 182268 463418 182352 463654
rect 182588 463418 185622 463654
rect 185858 463418 284098 463654
rect 284334 463418 290032 463654
rect 290268 463418 290352 463654
rect 290588 463418 310622 463654
rect 310858 463418 409098 463654
rect 409334 463418 434032 463654
rect 434268 463418 434352 463654
rect 434588 463418 436622 463654
rect 436858 463418 535098 463654
rect 535334 463418 542032 463654
rect 542268 463418 542352 463654
rect 542588 463418 571532 463654
rect 571768 463418 571852 463654
rect 572088 463418 586302 463654
rect 586538 463418 586622 463654
rect 586858 463418 586890 463654
rect -2966 463334 586890 463418
rect -2966 463098 -2934 463334
rect -2698 463098 -2614 463334
rect -2378 463098 7876 463334
rect 8112 463098 8196 463334
rect 8432 463098 38032 463334
rect 38268 463098 38352 463334
rect 38588 463098 60622 463334
rect 60858 463098 159098 463334
rect 159334 463098 182032 463334
rect 182268 463098 182352 463334
rect 182588 463098 185622 463334
rect 185858 463098 284098 463334
rect 284334 463098 290032 463334
rect 290268 463098 290352 463334
rect 290588 463098 310622 463334
rect 310858 463098 409098 463334
rect 409334 463098 434032 463334
rect 434268 463098 434352 463334
rect 434588 463098 436622 463334
rect 436858 463098 535098 463334
rect 535334 463098 542032 463334
rect 542268 463098 542352 463334
rect 542588 463098 571532 463334
rect 571768 463098 571852 463334
rect 572088 463098 586302 463334
rect 586538 463098 586622 463334
rect 586858 463098 586890 463334
rect -2966 463066 586890 463098
rect -8726 454814 592650 454846
rect -8726 454578 -7734 454814
rect -7498 454578 -7414 454814
rect -7178 454578 591102 454814
rect 591338 454578 591422 454814
rect 591658 454578 592650 454814
rect -8726 454494 592650 454578
rect -8726 454258 -7734 454494
rect -7498 454258 -7414 454494
rect -7178 454258 591102 454494
rect 591338 454258 591422 454494
rect 591658 454258 592650 454494
rect -8726 454226 592650 454258
rect -6806 451094 590730 451126
rect -6806 450858 -5814 451094
rect -5578 450858 -5494 451094
rect -5258 450858 589182 451094
rect 589418 450858 589502 451094
rect 589738 450858 590730 451094
rect -6806 450774 590730 450858
rect -6806 450538 -5814 450774
rect -5578 450538 -5494 450774
rect -5258 450538 589182 450774
rect 589418 450538 589502 450774
rect 589738 450538 590730 450774
rect -6806 450506 590730 450538
rect -4886 447374 588810 447406
rect -4886 447138 -3894 447374
rect -3658 447138 -3574 447374
rect -3338 447138 587262 447374
rect 587498 447138 587582 447374
rect 587818 447138 588810 447374
rect -4886 447054 588810 447138
rect -4886 446818 -3894 447054
rect -3658 446818 -3574 447054
rect -3338 446818 587262 447054
rect 587498 446818 587582 447054
rect 587818 446818 588810 447054
rect -4886 446786 588810 446818
rect -2966 443654 586890 443686
rect -2966 443418 -1974 443654
rect -1738 443418 -1654 443654
rect -1418 443418 9116 443654
rect 9352 443418 9436 443654
rect 9672 443418 56652 443654
rect 56888 443418 56972 443654
rect 57208 443418 61342 443654
rect 61578 443418 158378 443654
rect 158614 443418 164652 443654
rect 164888 443418 164972 443654
rect 165208 443418 186342 443654
rect 186578 443418 283378 443654
rect 283614 443418 308652 443654
rect 308888 443418 308972 443654
rect 309208 443418 311342 443654
rect 311578 443418 408378 443654
rect 408614 443418 416652 443654
rect 416888 443418 416972 443654
rect 417208 443418 437342 443654
rect 437578 443418 534378 443654
rect 534614 443418 560652 443654
rect 560888 443418 560972 443654
rect 561208 443418 570292 443654
rect 570528 443418 570612 443654
rect 570848 443418 585342 443654
rect 585578 443418 585662 443654
rect 585898 443418 586890 443654
rect -2966 443334 586890 443418
rect -2966 443098 -1974 443334
rect -1738 443098 -1654 443334
rect -1418 443098 9116 443334
rect 9352 443098 9436 443334
rect 9672 443098 56652 443334
rect 56888 443098 56972 443334
rect 57208 443098 61342 443334
rect 61578 443098 158378 443334
rect 158614 443098 164652 443334
rect 164888 443098 164972 443334
rect 165208 443098 186342 443334
rect 186578 443098 283378 443334
rect 283614 443098 308652 443334
rect 308888 443098 308972 443334
rect 309208 443098 311342 443334
rect 311578 443098 408378 443334
rect 408614 443098 416652 443334
rect 416888 443098 416972 443334
rect 417208 443098 437342 443334
rect 437578 443098 534378 443334
rect 534614 443098 560652 443334
rect 560888 443098 560972 443334
rect 561208 443098 570292 443334
rect 570528 443098 570612 443334
rect 570848 443098 585342 443334
rect 585578 443098 585662 443334
rect 585898 443098 586890 443334
rect -2966 443066 586890 443098
rect -8726 434814 592650 434846
rect -8726 434578 -8694 434814
rect -8458 434578 -8374 434814
rect -8138 434578 592062 434814
rect 592298 434578 592382 434814
rect 592618 434578 592650 434814
rect -8726 434494 592650 434578
rect -8726 434258 -8694 434494
rect -8458 434258 -8374 434494
rect -8138 434258 592062 434494
rect 592298 434258 592382 434494
rect 592618 434258 592650 434494
rect -8726 434226 592650 434258
rect -6806 431094 590730 431126
rect -6806 430858 -6774 431094
rect -6538 430858 -6454 431094
rect -6218 430858 590142 431094
rect 590378 430858 590462 431094
rect 590698 430858 590730 431094
rect -6806 430774 590730 430858
rect -6806 430538 -6774 430774
rect -6538 430538 -6454 430774
rect -6218 430538 590142 430774
rect 590378 430538 590462 430774
rect 590698 430538 590730 430774
rect -6806 430506 590730 430538
rect -4886 427374 588810 427406
rect -4886 427138 -4854 427374
rect -4618 427138 -4534 427374
rect -4298 427138 588222 427374
rect 588458 427138 588542 427374
rect 588778 427138 588810 427374
rect -4886 427054 588810 427138
rect -4886 426818 -4854 427054
rect -4618 426818 -4534 427054
rect -4298 426818 588222 427054
rect 588458 426818 588542 427054
rect 588778 426818 588810 427054
rect -4886 426786 588810 426818
rect -2966 423654 586890 423686
rect -2966 423418 -2934 423654
rect -2698 423418 -2614 423654
rect -2378 423418 7876 423654
rect 8112 423418 8196 423654
rect 8432 423418 38032 423654
rect 38268 423418 38352 423654
rect 38588 423418 74032 423654
rect 74268 423418 74352 423654
rect 74588 423418 110032 423654
rect 110268 423418 110352 423654
rect 110588 423418 146032 423654
rect 146268 423418 146352 423654
rect 146588 423418 182032 423654
rect 182268 423418 182352 423654
rect 182588 423418 218032 423654
rect 218268 423418 218352 423654
rect 218588 423418 254032 423654
rect 254268 423418 254352 423654
rect 254588 423418 290032 423654
rect 290268 423418 290352 423654
rect 290588 423418 326032 423654
rect 326268 423418 326352 423654
rect 326588 423418 362032 423654
rect 362268 423418 362352 423654
rect 362588 423418 398032 423654
rect 398268 423418 398352 423654
rect 398588 423418 434032 423654
rect 434268 423418 434352 423654
rect 434588 423418 470032 423654
rect 470268 423418 470352 423654
rect 470588 423418 506032 423654
rect 506268 423418 506352 423654
rect 506588 423418 542032 423654
rect 542268 423418 542352 423654
rect 542588 423418 571532 423654
rect 571768 423418 571852 423654
rect 572088 423418 586302 423654
rect 586538 423418 586622 423654
rect 586858 423418 586890 423654
rect -2966 423334 586890 423418
rect -2966 423098 -2934 423334
rect -2698 423098 -2614 423334
rect -2378 423098 7876 423334
rect 8112 423098 8196 423334
rect 8432 423098 38032 423334
rect 38268 423098 38352 423334
rect 38588 423098 74032 423334
rect 74268 423098 74352 423334
rect 74588 423098 110032 423334
rect 110268 423098 110352 423334
rect 110588 423098 146032 423334
rect 146268 423098 146352 423334
rect 146588 423098 182032 423334
rect 182268 423098 182352 423334
rect 182588 423098 218032 423334
rect 218268 423098 218352 423334
rect 218588 423098 254032 423334
rect 254268 423098 254352 423334
rect 254588 423098 290032 423334
rect 290268 423098 290352 423334
rect 290588 423098 326032 423334
rect 326268 423098 326352 423334
rect 326588 423098 362032 423334
rect 362268 423098 362352 423334
rect 362588 423098 398032 423334
rect 398268 423098 398352 423334
rect 398588 423098 434032 423334
rect 434268 423098 434352 423334
rect 434588 423098 470032 423334
rect 470268 423098 470352 423334
rect 470588 423098 506032 423334
rect 506268 423098 506352 423334
rect 506588 423098 542032 423334
rect 542268 423098 542352 423334
rect 542588 423098 571532 423334
rect 571768 423098 571852 423334
rect 572088 423098 586302 423334
rect 586538 423098 586622 423334
rect 586858 423098 586890 423334
rect -2966 423066 586890 423098
rect -8726 414814 592650 414846
rect -8726 414578 -7734 414814
rect -7498 414578 -7414 414814
rect -7178 414578 591102 414814
rect 591338 414578 591422 414814
rect 591658 414578 592650 414814
rect -8726 414494 592650 414578
rect -8726 414258 -7734 414494
rect -7498 414258 -7414 414494
rect -7178 414258 591102 414494
rect 591338 414258 591422 414494
rect 591658 414258 592650 414494
rect -8726 414226 592650 414258
rect -6806 411094 590730 411126
rect -6806 410858 -5814 411094
rect -5578 410858 -5494 411094
rect -5258 410858 589182 411094
rect 589418 410858 589502 411094
rect 589738 410858 590730 411094
rect -6806 410774 590730 410858
rect -6806 410538 -5814 410774
rect -5578 410538 -5494 410774
rect -5258 410538 589182 410774
rect 589418 410538 589502 410774
rect 589738 410538 590730 410774
rect -6806 410506 590730 410538
rect -4886 407374 588810 407406
rect -4886 407138 -3894 407374
rect -3658 407138 -3574 407374
rect -3338 407138 587262 407374
rect 587498 407138 587582 407374
rect 587818 407138 588810 407374
rect -4886 407054 588810 407138
rect -4886 406818 -3894 407054
rect -3658 406818 -3574 407054
rect -3338 406818 587262 407054
rect 587498 406818 587582 407054
rect 587818 406818 588810 407054
rect -4886 406786 588810 406818
rect -2966 403654 586890 403686
rect -2966 403418 -1974 403654
rect -1738 403418 -1654 403654
rect -1418 403418 9116 403654
rect 9352 403418 9436 403654
rect 9672 403418 56652 403654
rect 56888 403418 56972 403654
rect 57208 403418 92652 403654
rect 92888 403418 92972 403654
rect 93208 403418 128652 403654
rect 128888 403418 128972 403654
rect 129208 403418 164652 403654
rect 164888 403418 164972 403654
rect 165208 403418 200652 403654
rect 200888 403418 200972 403654
rect 201208 403418 236652 403654
rect 236888 403418 236972 403654
rect 237208 403418 272652 403654
rect 272888 403418 272972 403654
rect 273208 403418 308652 403654
rect 308888 403418 308972 403654
rect 309208 403418 344652 403654
rect 344888 403418 344972 403654
rect 345208 403418 380652 403654
rect 380888 403418 380972 403654
rect 381208 403418 416652 403654
rect 416888 403418 416972 403654
rect 417208 403418 452652 403654
rect 452888 403418 452972 403654
rect 453208 403418 488652 403654
rect 488888 403418 488972 403654
rect 489208 403418 524652 403654
rect 524888 403418 524972 403654
rect 525208 403418 560652 403654
rect 560888 403418 560972 403654
rect 561208 403418 570292 403654
rect 570528 403418 570612 403654
rect 570848 403418 585342 403654
rect 585578 403418 585662 403654
rect 585898 403418 586890 403654
rect -2966 403334 586890 403418
rect -2966 403098 -1974 403334
rect -1738 403098 -1654 403334
rect -1418 403098 9116 403334
rect 9352 403098 9436 403334
rect 9672 403098 56652 403334
rect 56888 403098 56972 403334
rect 57208 403098 92652 403334
rect 92888 403098 92972 403334
rect 93208 403098 128652 403334
rect 128888 403098 128972 403334
rect 129208 403098 164652 403334
rect 164888 403098 164972 403334
rect 165208 403098 200652 403334
rect 200888 403098 200972 403334
rect 201208 403098 236652 403334
rect 236888 403098 236972 403334
rect 237208 403098 272652 403334
rect 272888 403098 272972 403334
rect 273208 403098 308652 403334
rect 308888 403098 308972 403334
rect 309208 403098 344652 403334
rect 344888 403098 344972 403334
rect 345208 403098 380652 403334
rect 380888 403098 380972 403334
rect 381208 403098 416652 403334
rect 416888 403098 416972 403334
rect 417208 403098 452652 403334
rect 452888 403098 452972 403334
rect 453208 403098 488652 403334
rect 488888 403098 488972 403334
rect 489208 403098 524652 403334
rect 524888 403098 524972 403334
rect 525208 403098 560652 403334
rect 560888 403098 560972 403334
rect 561208 403098 570292 403334
rect 570528 403098 570612 403334
rect 570848 403098 585342 403334
rect 585578 403098 585662 403334
rect 585898 403098 586890 403334
rect -2966 403066 586890 403098
rect -8726 394814 592650 394846
rect -8726 394578 -8694 394814
rect -8458 394578 -8374 394814
rect -8138 394578 592062 394814
rect 592298 394578 592382 394814
rect 592618 394578 592650 394814
rect -8726 394494 592650 394578
rect -8726 394258 -8694 394494
rect -8458 394258 -8374 394494
rect -8138 394258 592062 394494
rect 592298 394258 592382 394494
rect 592618 394258 592650 394494
rect -8726 394226 592650 394258
rect -6806 391094 590730 391126
rect -6806 390858 -6774 391094
rect -6538 390858 -6454 391094
rect -6218 390858 590142 391094
rect 590378 390858 590462 391094
rect 590698 390858 590730 391094
rect -6806 390774 590730 390858
rect -6806 390538 -6774 390774
rect -6538 390538 -6454 390774
rect -6218 390538 590142 390774
rect 590378 390538 590462 390774
rect 590698 390538 590730 390774
rect -6806 390506 590730 390538
rect -4886 387374 588810 387406
rect -4886 387138 -4854 387374
rect -4618 387138 -4534 387374
rect -4298 387138 588222 387374
rect 588458 387138 588542 387374
rect 588778 387138 588810 387374
rect -4886 387054 588810 387138
rect -4886 386818 -4854 387054
rect -4618 386818 -4534 387054
rect -4298 386818 588222 387054
rect 588458 386818 588542 387054
rect 588778 386818 588810 387054
rect -4886 386786 588810 386818
rect -2966 383654 586890 383686
rect -2966 383418 -2934 383654
rect -2698 383418 -2614 383654
rect -2378 383418 7876 383654
rect 8112 383418 8196 383654
rect 8432 383418 38032 383654
rect 38268 383418 38352 383654
rect 38588 383418 74032 383654
rect 74268 383418 74352 383654
rect 74588 383418 110032 383654
rect 110268 383418 110352 383654
rect 110588 383418 146032 383654
rect 146268 383418 146352 383654
rect 146588 383418 182032 383654
rect 182268 383418 182352 383654
rect 182588 383418 218032 383654
rect 218268 383418 218352 383654
rect 218588 383418 254032 383654
rect 254268 383418 254352 383654
rect 254588 383418 290032 383654
rect 290268 383418 290352 383654
rect 290588 383418 326032 383654
rect 326268 383418 326352 383654
rect 326588 383418 362032 383654
rect 362268 383418 362352 383654
rect 362588 383418 398032 383654
rect 398268 383418 398352 383654
rect 398588 383418 434032 383654
rect 434268 383418 434352 383654
rect 434588 383418 470032 383654
rect 470268 383418 470352 383654
rect 470588 383418 506032 383654
rect 506268 383418 506352 383654
rect 506588 383418 542032 383654
rect 542268 383418 542352 383654
rect 542588 383418 571532 383654
rect 571768 383418 571852 383654
rect 572088 383418 586302 383654
rect 586538 383418 586622 383654
rect 586858 383418 586890 383654
rect -2966 383334 586890 383418
rect -2966 383098 -2934 383334
rect -2698 383098 -2614 383334
rect -2378 383098 7876 383334
rect 8112 383098 8196 383334
rect 8432 383098 38032 383334
rect 38268 383098 38352 383334
rect 38588 383098 74032 383334
rect 74268 383098 74352 383334
rect 74588 383098 110032 383334
rect 110268 383098 110352 383334
rect 110588 383098 146032 383334
rect 146268 383098 146352 383334
rect 146588 383098 182032 383334
rect 182268 383098 182352 383334
rect 182588 383098 218032 383334
rect 218268 383098 218352 383334
rect 218588 383098 254032 383334
rect 254268 383098 254352 383334
rect 254588 383098 290032 383334
rect 290268 383098 290352 383334
rect 290588 383098 326032 383334
rect 326268 383098 326352 383334
rect 326588 383098 362032 383334
rect 362268 383098 362352 383334
rect 362588 383098 398032 383334
rect 398268 383098 398352 383334
rect 398588 383098 434032 383334
rect 434268 383098 434352 383334
rect 434588 383098 470032 383334
rect 470268 383098 470352 383334
rect 470588 383098 506032 383334
rect 506268 383098 506352 383334
rect 506588 383098 542032 383334
rect 542268 383098 542352 383334
rect 542588 383098 571532 383334
rect 571768 383098 571852 383334
rect 572088 383098 586302 383334
rect 586538 383098 586622 383334
rect 586858 383098 586890 383334
rect -2966 383066 586890 383098
rect -8726 374814 592650 374846
rect -8726 374578 -7734 374814
rect -7498 374578 -7414 374814
rect -7178 374578 591102 374814
rect 591338 374578 591422 374814
rect 591658 374578 592650 374814
rect -8726 374494 592650 374578
rect -8726 374258 -7734 374494
rect -7498 374258 -7414 374494
rect -7178 374258 591102 374494
rect 591338 374258 591422 374494
rect 591658 374258 592650 374494
rect -8726 374226 592650 374258
rect -6806 371094 590730 371126
rect -6806 370858 -5814 371094
rect -5578 370858 -5494 371094
rect -5258 370858 589182 371094
rect 589418 370858 589502 371094
rect 589738 370858 590730 371094
rect -6806 370774 590730 370858
rect -6806 370538 -5814 370774
rect -5578 370538 -5494 370774
rect -5258 370538 589182 370774
rect 589418 370538 589502 370774
rect 589738 370538 590730 370774
rect -6806 370506 590730 370538
rect -4886 367374 588810 367406
rect -4886 367138 -3894 367374
rect -3658 367138 -3574 367374
rect -3338 367138 587262 367374
rect 587498 367138 587582 367374
rect 587818 367138 588810 367374
rect -4886 367054 588810 367138
rect -4886 366818 -3894 367054
rect -3658 366818 -3574 367054
rect -3338 366818 587262 367054
rect 587498 366818 587582 367054
rect 587818 366818 588810 367054
rect -4886 366786 588810 366818
rect -2966 363654 586890 363686
rect -2966 363418 -1974 363654
rect -1738 363418 -1654 363654
rect -1418 363418 9116 363654
rect 9352 363418 9436 363654
rect 9672 363418 56652 363654
rect 56888 363418 56972 363654
rect 57208 363418 92652 363654
rect 92888 363418 92972 363654
rect 93208 363418 128652 363654
rect 128888 363418 128972 363654
rect 129208 363418 164652 363654
rect 164888 363418 164972 363654
rect 165208 363418 200652 363654
rect 200888 363418 200972 363654
rect 201208 363418 236652 363654
rect 236888 363418 236972 363654
rect 237208 363418 272652 363654
rect 272888 363418 272972 363654
rect 273208 363418 308652 363654
rect 308888 363418 308972 363654
rect 309208 363418 344652 363654
rect 344888 363418 344972 363654
rect 345208 363418 380652 363654
rect 380888 363418 380972 363654
rect 381208 363418 416652 363654
rect 416888 363418 416972 363654
rect 417208 363418 452652 363654
rect 452888 363418 452972 363654
rect 453208 363418 488652 363654
rect 488888 363418 488972 363654
rect 489208 363418 524652 363654
rect 524888 363418 524972 363654
rect 525208 363418 560652 363654
rect 560888 363418 560972 363654
rect 561208 363418 570292 363654
rect 570528 363418 570612 363654
rect 570848 363418 585342 363654
rect 585578 363418 585662 363654
rect 585898 363418 586890 363654
rect -2966 363334 586890 363418
rect -2966 363098 -1974 363334
rect -1738 363098 -1654 363334
rect -1418 363098 9116 363334
rect 9352 363098 9436 363334
rect 9672 363098 56652 363334
rect 56888 363098 56972 363334
rect 57208 363098 92652 363334
rect 92888 363098 92972 363334
rect 93208 363098 128652 363334
rect 128888 363098 128972 363334
rect 129208 363098 164652 363334
rect 164888 363098 164972 363334
rect 165208 363098 200652 363334
rect 200888 363098 200972 363334
rect 201208 363098 236652 363334
rect 236888 363098 236972 363334
rect 237208 363098 272652 363334
rect 272888 363098 272972 363334
rect 273208 363098 308652 363334
rect 308888 363098 308972 363334
rect 309208 363098 344652 363334
rect 344888 363098 344972 363334
rect 345208 363098 380652 363334
rect 380888 363098 380972 363334
rect 381208 363098 416652 363334
rect 416888 363098 416972 363334
rect 417208 363098 452652 363334
rect 452888 363098 452972 363334
rect 453208 363098 488652 363334
rect 488888 363098 488972 363334
rect 489208 363098 524652 363334
rect 524888 363098 524972 363334
rect 525208 363098 560652 363334
rect 560888 363098 560972 363334
rect 561208 363098 570292 363334
rect 570528 363098 570612 363334
rect 570848 363098 585342 363334
rect 585578 363098 585662 363334
rect 585898 363098 586890 363334
rect -2966 363066 586890 363098
rect -8726 354814 592650 354846
rect -8726 354578 -8694 354814
rect -8458 354578 -8374 354814
rect -8138 354578 592062 354814
rect 592298 354578 592382 354814
rect 592618 354578 592650 354814
rect -8726 354494 592650 354578
rect -8726 354258 -8694 354494
rect -8458 354258 -8374 354494
rect -8138 354258 592062 354494
rect 592298 354258 592382 354494
rect 592618 354258 592650 354494
rect -8726 354226 592650 354258
rect -6806 351094 590730 351126
rect -6806 350858 -6774 351094
rect -6538 350858 -6454 351094
rect -6218 350858 590142 351094
rect 590378 350858 590462 351094
rect 590698 350858 590730 351094
rect -6806 350774 590730 350858
rect -6806 350538 -6774 350774
rect -6538 350538 -6454 350774
rect -6218 350538 590142 350774
rect 590378 350538 590462 350774
rect 590698 350538 590730 350774
rect -6806 350506 590730 350538
rect -4886 347374 588810 347406
rect -4886 347138 -4854 347374
rect -4618 347138 -4534 347374
rect -4298 347138 588222 347374
rect 588458 347138 588542 347374
rect 588778 347138 588810 347374
rect -4886 347054 588810 347138
rect -4886 346818 -4854 347054
rect -4618 346818 -4534 347054
rect -4298 346818 588222 347054
rect 588458 346818 588542 347054
rect 588778 346818 588810 347054
rect -4886 346786 588810 346818
rect -2966 343654 586890 343686
rect -2966 343418 -2934 343654
rect -2698 343418 -2614 343654
rect -2378 343418 7876 343654
rect 8112 343418 8196 343654
rect 8432 343418 38032 343654
rect 38268 343418 38352 343654
rect 38588 343418 74032 343654
rect 74268 343418 74352 343654
rect 74588 343418 110032 343654
rect 110268 343418 110352 343654
rect 110588 343418 146032 343654
rect 146268 343418 146352 343654
rect 146588 343418 182032 343654
rect 182268 343418 182352 343654
rect 182588 343418 218032 343654
rect 218268 343418 218352 343654
rect 218588 343418 254032 343654
rect 254268 343418 254352 343654
rect 254588 343418 290032 343654
rect 290268 343418 290352 343654
rect 290588 343418 326032 343654
rect 326268 343418 326352 343654
rect 326588 343418 362032 343654
rect 362268 343418 362352 343654
rect 362588 343418 398032 343654
rect 398268 343418 398352 343654
rect 398588 343418 434032 343654
rect 434268 343418 434352 343654
rect 434588 343418 470032 343654
rect 470268 343418 470352 343654
rect 470588 343418 506032 343654
rect 506268 343418 506352 343654
rect 506588 343418 542032 343654
rect 542268 343418 542352 343654
rect 542588 343418 571532 343654
rect 571768 343418 571852 343654
rect 572088 343418 586302 343654
rect 586538 343418 586622 343654
rect 586858 343418 586890 343654
rect -2966 343334 586890 343418
rect -2966 343098 -2934 343334
rect -2698 343098 -2614 343334
rect -2378 343098 7876 343334
rect 8112 343098 8196 343334
rect 8432 343098 38032 343334
rect 38268 343098 38352 343334
rect 38588 343098 74032 343334
rect 74268 343098 74352 343334
rect 74588 343098 110032 343334
rect 110268 343098 110352 343334
rect 110588 343098 146032 343334
rect 146268 343098 146352 343334
rect 146588 343098 182032 343334
rect 182268 343098 182352 343334
rect 182588 343098 218032 343334
rect 218268 343098 218352 343334
rect 218588 343098 254032 343334
rect 254268 343098 254352 343334
rect 254588 343098 290032 343334
rect 290268 343098 290352 343334
rect 290588 343098 326032 343334
rect 326268 343098 326352 343334
rect 326588 343098 362032 343334
rect 362268 343098 362352 343334
rect 362588 343098 398032 343334
rect 398268 343098 398352 343334
rect 398588 343098 434032 343334
rect 434268 343098 434352 343334
rect 434588 343098 470032 343334
rect 470268 343098 470352 343334
rect 470588 343098 506032 343334
rect 506268 343098 506352 343334
rect 506588 343098 542032 343334
rect 542268 343098 542352 343334
rect 542588 343098 571532 343334
rect 571768 343098 571852 343334
rect 572088 343098 586302 343334
rect 586538 343098 586622 343334
rect 586858 343098 586890 343334
rect -2966 343066 586890 343098
rect -8726 334814 592650 334846
rect -8726 334578 -7734 334814
rect -7498 334578 -7414 334814
rect -7178 334578 591102 334814
rect 591338 334578 591422 334814
rect 591658 334578 592650 334814
rect -8726 334494 592650 334578
rect -8726 334258 -7734 334494
rect -7498 334258 -7414 334494
rect -7178 334258 591102 334494
rect 591338 334258 591422 334494
rect 591658 334258 592650 334494
rect -8726 334226 592650 334258
rect -6806 331094 590730 331126
rect -6806 330858 -5814 331094
rect -5578 330858 -5494 331094
rect -5258 330858 589182 331094
rect 589418 330858 589502 331094
rect 589738 330858 590730 331094
rect -6806 330774 590730 330858
rect -6806 330538 -5814 330774
rect -5578 330538 -5494 330774
rect -5258 330538 589182 330774
rect 589418 330538 589502 330774
rect 589738 330538 590730 330774
rect -6806 330506 590730 330538
rect -4886 327374 588810 327406
rect -4886 327138 -3894 327374
rect -3658 327138 -3574 327374
rect -3338 327138 587262 327374
rect 587498 327138 587582 327374
rect 587818 327138 588810 327374
rect -4886 327054 588810 327138
rect -4886 326818 -3894 327054
rect -3658 326818 -3574 327054
rect -3338 326818 587262 327054
rect 587498 326818 587582 327054
rect 587818 326818 588810 327054
rect -4886 326786 588810 326818
rect -2966 323654 586890 323686
rect -2966 323418 -1974 323654
rect -1738 323418 -1654 323654
rect -1418 323418 9116 323654
rect 9352 323418 9436 323654
rect 9672 323418 56652 323654
rect 56888 323418 56972 323654
rect 57208 323418 92652 323654
rect 92888 323418 92972 323654
rect 93208 323418 128652 323654
rect 128888 323418 128972 323654
rect 129208 323418 164652 323654
rect 164888 323418 164972 323654
rect 165208 323418 200652 323654
rect 200888 323418 200972 323654
rect 201208 323418 236652 323654
rect 236888 323418 236972 323654
rect 237208 323418 272652 323654
rect 272888 323418 272972 323654
rect 273208 323418 308652 323654
rect 308888 323418 308972 323654
rect 309208 323418 344652 323654
rect 344888 323418 344972 323654
rect 345208 323418 380652 323654
rect 380888 323418 380972 323654
rect 381208 323418 416652 323654
rect 416888 323418 416972 323654
rect 417208 323418 452652 323654
rect 452888 323418 452972 323654
rect 453208 323418 488652 323654
rect 488888 323418 488972 323654
rect 489208 323418 524652 323654
rect 524888 323418 524972 323654
rect 525208 323418 560652 323654
rect 560888 323418 560972 323654
rect 561208 323418 570292 323654
rect 570528 323418 570612 323654
rect 570848 323418 585342 323654
rect 585578 323418 585662 323654
rect 585898 323418 586890 323654
rect -2966 323334 586890 323418
rect -2966 323098 -1974 323334
rect -1738 323098 -1654 323334
rect -1418 323098 9116 323334
rect 9352 323098 9436 323334
rect 9672 323098 56652 323334
rect 56888 323098 56972 323334
rect 57208 323098 92652 323334
rect 92888 323098 92972 323334
rect 93208 323098 128652 323334
rect 128888 323098 128972 323334
rect 129208 323098 164652 323334
rect 164888 323098 164972 323334
rect 165208 323098 200652 323334
rect 200888 323098 200972 323334
rect 201208 323098 236652 323334
rect 236888 323098 236972 323334
rect 237208 323098 272652 323334
rect 272888 323098 272972 323334
rect 273208 323098 308652 323334
rect 308888 323098 308972 323334
rect 309208 323098 344652 323334
rect 344888 323098 344972 323334
rect 345208 323098 380652 323334
rect 380888 323098 380972 323334
rect 381208 323098 416652 323334
rect 416888 323098 416972 323334
rect 417208 323098 452652 323334
rect 452888 323098 452972 323334
rect 453208 323098 488652 323334
rect 488888 323098 488972 323334
rect 489208 323098 524652 323334
rect 524888 323098 524972 323334
rect 525208 323098 560652 323334
rect 560888 323098 560972 323334
rect 561208 323098 570292 323334
rect 570528 323098 570612 323334
rect 570848 323098 585342 323334
rect 585578 323098 585662 323334
rect 585898 323098 586890 323334
rect -2966 323066 586890 323098
rect -8726 314814 592650 314846
rect -8726 314578 -8694 314814
rect -8458 314578 -8374 314814
rect -8138 314578 592062 314814
rect 592298 314578 592382 314814
rect 592618 314578 592650 314814
rect -8726 314494 592650 314578
rect -8726 314258 -8694 314494
rect -8458 314258 -8374 314494
rect -8138 314258 592062 314494
rect 592298 314258 592382 314494
rect 592618 314258 592650 314494
rect -8726 314226 592650 314258
rect -6806 311094 590730 311126
rect -6806 310858 -6774 311094
rect -6538 310858 -6454 311094
rect -6218 310858 590142 311094
rect 590378 310858 590462 311094
rect 590698 310858 590730 311094
rect -6806 310774 590730 310858
rect -6806 310538 -6774 310774
rect -6538 310538 -6454 310774
rect -6218 310538 590142 310774
rect 590378 310538 590462 310774
rect 590698 310538 590730 310774
rect -6806 310506 590730 310538
rect -4886 307374 588810 307406
rect -4886 307138 -4854 307374
rect -4618 307138 -4534 307374
rect -4298 307138 588222 307374
rect 588458 307138 588542 307374
rect 588778 307138 588810 307374
rect -4886 307054 588810 307138
rect -4886 306818 -4854 307054
rect -4618 306818 -4534 307054
rect -4298 306818 588222 307054
rect 588458 306818 588542 307054
rect 588778 306818 588810 307054
rect -4886 306786 588810 306818
rect -2966 303654 586890 303686
rect -2966 303418 -2934 303654
rect -2698 303418 -2614 303654
rect -2378 303418 7876 303654
rect 8112 303418 8196 303654
rect 8432 303418 38032 303654
rect 38268 303418 38352 303654
rect 38588 303418 74032 303654
rect 74268 303418 74352 303654
rect 74588 303418 110032 303654
rect 110268 303418 110352 303654
rect 110588 303418 146032 303654
rect 146268 303418 146352 303654
rect 146588 303418 182032 303654
rect 182268 303418 182352 303654
rect 182588 303418 218032 303654
rect 218268 303418 218352 303654
rect 218588 303418 254032 303654
rect 254268 303418 254352 303654
rect 254588 303418 290032 303654
rect 290268 303418 290352 303654
rect 290588 303418 326032 303654
rect 326268 303418 326352 303654
rect 326588 303418 362032 303654
rect 362268 303418 362352 303654
rect 362588 303418 398032 303654
rect 398268 303418 398352 303654
rect 398588 303418 434032 303654
rect 434268 303418 434352 303654
rect 434588 303418 470032 303654
rect 470268 303418 470352 303654
rect 470588 303418 506032 303654
rect 506268 303418 506352 303654
rect 506588 303418 542032 303654
rect 542268 303418 542352 303654
rect 542588 303418 571532 303654
rect 571768 303418 571852 303654
rect 572088 303418 586302 303654
rect 586538 303418 586622 303654
rect 586858 303418 586890 303654
rect -2966 303334 586890 303418
rect -2966 303098 -2934 303334
rect -2698 303098 -2614 303334
rect -2378 303098 7876 303334
rect 8112 303098 8196 303334
rect 8432 303098 38032 303334
rect 38268 303098 38352 303334
rect 38588 303098 74032 303334
rect 74268 303098 74352 303334
rect 74588 303098 110032 303334
rect 110268 303098 110352 303334
rect 110588 303098 146032 303334
rect 146268 303098 146352 303334
rect 146588 303098 182032 303334
rect 182268 303098 182352 303334
rect 182588 303098 218032 303334
rect 218268 303098 218352 303334
rect 218588 303098 254032 303334
rect 254268 303098 254352 303334
rect 254588 303098 290032 303334
rect 290268 303098 290352 303334
rect 290588 303098 326032 303334
rect 326268 303098 326352 303334
rect 326588 303098 362032 303334
rect 362268 303098 362352 303334
rect 362588 303098 398032 303334
rect 398268 303098 398352 303334
rect 398588 303098 434032 303334
rect 434268 303098 434352 303334
rect 434588 303098 470032 303334
rect 470268 303098 470352 303334
rect 470588 303098 506032 303334
rect 506268 303098 506352 303334
rect 506588 303098 542032 303334
rect 542268 303098 542352 303334
rect 542588 303098 571532 303334
rect 571768 303098 571852 303334
rect 572088 303098 586302 303334
rect 586538 303098 586622 303334
rect 586858 303098 586890 303334
rect -2966 303066 586890 303098
rect -8726 294814 592650 294846
rect -8726 294578 -7734 294814
rect -7498 294578 -7414 294814
rect -7178 294578 591102 294814
rect 591338 294578 591422 294814
rect 591658 294578 592650 294814
rect -8726 294494 592650 294578
rect -8726 294258 -7734 294494
rect -7498 294258 -7414 294494
rect -7178 294258 591102 294494
rect 591338 294258 591422 294494
rect 591658 294258 592650 294494
rect -8726 294226 592650 294258
rect -6806 291094 590730 291126
rect -6806 290858 -5814 291094
rect -5578 290858 -5494 291094
rect -5258 290858 589182 291094
rect 589418 290858 589502 291094
rect 589738 290858 590730 291094
rect -6806 290774 590730 290858
rect -6806 290538 -5814 290774
rect -5578 290538 -5494 290774
rect -5258 290538 589182 290774
rect 589418 290538 589502 290774
rect 589738 290538 590730 290774
rect -6806 290506 590730 290538
rect -4886 287374 588810 287406
rect -4886 287138 -3894 287374
rect -3658 287138 -3574 287374
rect -3338 287138 587262 287374
rect 587498 287138 587582 287374
rect 587818 287138 588810 287374
rect -4886 287054 588810 287138
rect -4886 286818 -3894 287054
rect -3658 286818 -3574 287054
rect -3338 286818 587262 287054
rect 587498 286818 587582 287054
rect 587818 286818 588810 287054
rect -4886 286786 588810 286818
rect -2966 283654 586890 283686
rect -2966 283418 -1974 283654
rect -1738 283418 -1654 283654
rect -1418 283418 9116 283654
rect 9352 283418 9436 283654
rect 9672 283418 56652 283654
rect 56888 283418 56972 283654
rect 57208 283418 92652 283654
rect 92888 283418 92972 283654
rect 93208 283418 128652 283654
rect 128888 283418 128972 283654
rect 129208 283418 164652 283654
rect 164888 283418 164972 283654
rect 165208 283418 200652 283654
rect 200888 283418 200972 283654
rect 201208 283418 236652 283654
rect 236888 283418 236972 283654
rect 237208 283418 272652 283654
rect 272888 283418 272972 283654
rect 273208 283418 308652 283654
rect 308888 283418 308972 283654
rect 309208 283418 344652 283654
rect 344888 283418 344972 283654
rect 345208 283418 380652 283654
rect 380888 283418 380972 283654
rect 381208 283418 416652 283654
rect 416888 283418 416972 283654
rect 417208 283418 452652 283654
rect 452888 283418 452972 283654
rect 453208 283418 488652 283654
rect 488888 283418 488972 283654
rect 489208 283418 524652 283654
rect 524888 283418 524972 283654
rect 525208 283418 560652 283654
rect 560888 283418 560972 283654
rect 561208 283418 570292 283654
rect 570528 283418 570612 283654
rect 570848 283418 585342 283654
rect 585578 283418 585662 283654
rect 585898 283418 586890 283654
rect -2966 283334 586890 283418
rect -2966 283098 -1974 283334
rect -1738 283098 -1654 283334
rect -1418 283098 9116 283334
rect 9352 283098 9436 283334
rect 9672 283098 56652 283334
rect 56888 283098 56972 283334
rect 57208 283098 92652 283334
rect 92888 283098 92972 283334
rect 93208 283098 128652 283334
rect 128888 283098 128972 283334
rect 129208 283098 164652 283334
rect 164888 283098 164972 283334
rect 165208 283098 200652 283334
rect 200888 283098 200972 283334
rect 201208 283098 236652 283334
rect 236888 283098 236972 283334
rect 237208 283098 272652 283334
rect 272888 283098 272972 283334
rect 273208 283098 308652 283334
rect 308888 283098 308972 283334
rect 309208 283098 344652 283334
rect 344888 283098 344972 283334
rect 345208 283098 380652 283334
rect 380888 283098 380972 283334
rect 381208 283098 416652 283334
rect 416888 283098 416972 283334
rect 417208 283098 452652 283334
rect 452888 283098 452972 283334
rect 453208 283098 488652 283334
rect 488888 283098 488972 283334
rect 489208 283098 524652 283334
rect 524888 283098 524972 283334
rect 525208 283098 560652 283334
rect 560888 283098 560972 283334
rect 561208 283098 570292 283334
rect 570528 283098 570612 283334
rect 570848 283098 585342 283334
rect 585578 283098 585662 283334
rect 585898 283098 586890 283334
rect -2966 283066 586890 283098
rect -8726 274814 592650 274846
rect -8726 274578 -8694 274814
rect -8458 274578 -8374 274814
rect -8138 274578 592062 274814
rect 592298 274578 592382 274814
rect 592618 274578 592650 274814
rect -8726 274494 592650 274578
rect -8726 274258 -8694 274494
rect -8458 274258 -8374 274494
rect -8138 274258 592062 274494
rect 592298 274258 592382 274494
rect 592618 274258 592650 274494
rect -8726 274226 592650 274258
rect -6806 271094 590730 271126
rect -6806 270858 -6774 271094
rect -6538 270858 -6454 271094
rect -6218 270858 590142 271094
rect 590378 270858 590462 271094
rect 590698 270858 590730 271094
rect -6806 270774 590730 270858
rect -6806 270538 -6774 270774
rect -6538 270538 -6454 270774
rect -6218 270538 590142 270774
rect 590378 270538 590462 270774
rect 590698 270538 590730 270774
rect -6806 270506 590730 270538
rect -4886 267374 588810 267406
rect -4886 267138 -4854 267374
rect -4618 267138 -4534 267374
rect -4298 267138 588222 267374
rect 588458 267138 588542 267374
rect 588778 267138 588810 267374
rect -4886 267054 588810 267138
rect -4886 266818 -4854 267054
rect -4618 266818 -4534 267054
rect -4298 266818 588222 267054
rect 588458 266818 588542 267054
rect 588778 266818 588810 267054
rect -4886 266786 588810 266818
rect -2966 263654 586890 263686
rect -2966 263418 -2934 263654
rect -2698 263418 -2614 263654
rect -2378 263418 7876 263654
rect 8112 263418 8196 263654
rect 8432 263418 38032 263654
rect 38268 263418 38352 263654
rect 38588 263418 74032 263654
rect 74268 263418 74352 263654
rect 74588 263418 110032 263654
rect 110268 263418 110352 263654
rect 110588 263418 146032 263654
rect 146268 263418 146352 263654
rect 146588 263418 182032 263654
rect 182268 263418 182352 263654
rect 182588 263418 218032 263654
rect 218268 263418 218352 263654
rect 218588 263418 254032 263654
rect 254268 263418 254352 263654
rect 254588 263418 290032 263654
rect 290268 263418 290352 263654
rect 290588 263418 326032 263654
rect 326268 263418 326352 263654
rect 326588 263418 362032 263654
rect 362268 263418 362352 263654
rect 362588 263418 398032 263654
rect 398268 263418 398352 263654
rect 398588 263418 434032 263654
rect 434268 263418 434352 263654
rect 434588 263418 470032 263654
rect 470268 263418 470352 263654
rect 470588 263418 506032 263654
rect 506268 263418 506352 263654
rect 506588 263418 542032 263654
rect 542268 263418 542352 263654
rect 542588 263418 571532 263654
rect 571768 263418 571852 263654
rect 572088 263418 586302 263654
rect 586538 263418 586622 263654
rect 586858 263418 586890 263654
rect -2966 263334 586890 263418
rect -2966 263098 -2934 263334
rect -2698 263098 -2614 263334
rect -2378 263098 7876 263334
rect 8112 263098 8196 263334
rect 8432 263098 38032 263334
rect 38268 263098 38352 263334
rect 38588 263098 74032 263334
rect 74268 263098 74352 263334
rect 74588 263098 110032 263334
rect 110268 263098 110352 263334
rect 110588 263098 146032 263334
rect 146268 263098 146352 263334
rect 146588 263098 182032 263334
rect 182268 263098 182352 263334
rect 182588 263098 218032 263334
rect 218268 263098 218352 263334
rect 218588 263098 254032 263334
rect 254268 263098 254352 263334
rect 254588 263098 290032 263334
rect 290268 263098 290352 263334
rect 290588 263098 326032 263334
rect 326268 263098 326352 263334
rect 326588 263098 362032 263334
rect 362268 263098 362352 263334
rect 362588 263098 398032 263334
rect 398268 263098 398352 263334
rect 398588 263098 434032 263334
rect 434268 263098 434352 263334
rect 434588 263098 470032 263334
rect 470268 263098 470352 263334
rect 470588 263098 506032 263334
rect 506268 263098 506352 263334
rect 506588 263098 542032 263334
rect 542268 263098 542352 263334
rect 542588 263098 571532 263334
rect 571768 263098 571852 263334
rect 572088 263098 586302 263334
rect 586538 263098 586622 263334
rect 586858 263098 586890 263334
rect -2966 263066 586890 263098
rect -8726 254814 592650 254846
rect -8726 254578 -7734 254814
rect -7498 254578 -7414 254814
rect -7178 254578 591102 254814
rect 591338 254578 591422 254814
rect 591658 254578 592650 254814
rect -8726 254494 592650 254578
rect -8726 254258 -7734 254494
rect -7498 254258 -7414 254494
rect -7178 254258 591102 254494
rect 591338 254258 591422 254494
rect 591658 254258 592650 254494
rect -8726 254226 592650 254258
rect -6806 251094 590730 251126
rect -6806 250858 -5814 251094
rect -5578 250858 -5494 251094
rect -5258 250858 589182 251094
rect 589418 250858 589502 251094
rect 589738 250858 590730 251094
rect -6806 250774 590730 250858
rect -6806 250538 -5814 250774
rect -5578 250538 -5494 250774
rect -5258 250538 589182 250774
rect 589418 250538 589502 250774
rect 589738 250538 590730 250774
rect -6806 250506 590730 250538
rect -4886 247374 588810 247406
rect -4886 247138 -3894 247374
rect -3658 247138 -3574 247374
rect -3338 247138 587262 247374
rect 587498 247138 587582 247374
rect 587818 247138 588810 247374
rect -4886 247054 588810 247138
rect -4886 246818 -3894 247054
rect -3658 246818 -3574 247054
rect -3338 246818 587262 247054
rect 587498 246818 587582 247054
rect 587818 246818 588810 247054
rect -4886 246786 588810 246818
rect -2966 243654 586890 243686
rect -2966 243418 -1974 243654
rect -1738 243418 -1654 243654
rect -1418 243418 9116 243654
rect 9352 243418 9436 243654
rect 9672 243418 56652 243654
rect 56888 243418 56972 243654
rect 57208 243418 92652 243654
rect 92888 243418 92972 243654
rect 93208 243418 128652 243654
rect 128888 243418 128972 243654
rect 129208 243418 164652 243654
rect 164888 243418 164972 243654
rect 165208 243418 200652 243654
rect 200888 243418 200972 243654
rect 201208 243418 236652 243654
rect 236888 243418 236972 243654
rect 237208 243418 272652 243654
rect 272888 243418 272972 243654
rect 273208 243418 308652 243654
rect 308888 243418 308972 243654
rect 309208 243418 344652 243654
rect 344888 243418 344972 243654
rect 345208 243418 380652 243654
rect 380888 243418 380972 243654
rect 381208 243418 416652 243654
rect 416888 243418 416972 243654
rect 417208 243418 452652 243654
rect 452888 243418 452972 243654
rect 453208 243418 488652 243654
rect 488888 243418 488972 243654
rect 489208 243418 524652 243654
rect 524888 243418 524972 243654
rect 525208 243418 560652 243654
rect 560888 243418 560972 243654
rect 561208 243418 570292 243654
rect 570528 243418 570612 243654
rect 570848 243418 585342 243654
rect 585578 243418 585662 243654
rect 585898 243418 586890 243654
rect -2966 243334 586890 243418
rect -2966 243098 -1974 243334
rect -1738 243098 -1654 243334
rect -1418 243098 9116 243334
rect 9352 243098 9436 243334
rect 9672 243098 56652 243334
rect 56888 243098 56972 243334
rect 57208 243098 92652 243334
rect 92888 243098 92972 243334
rect 93208 243098 128652 243334
rect 128888 243098 128972 243334
rect 129208 243098 164652 243334
rect 164888 243098 164972 243334
rect 165208 243098 200652 243334
rect 200888 243098 200972 243334
rect 201208 243098 236652 243334
rect 236888 243098 236972 243334
rect 237208 243098 272652 243334
rect 272888 243098 272972 243334
rect 273208 243098 308652 243334
rect 308888 243098 308972 243334
rect 309208 243098 344652 243334
rect 344888 243098 344972 243334
rect 345208 243098 380652 243334
rect 380888 243098 380972 243334
rect 381208 243098 416652 243334
rect 416888 243098 416972 243334
rect 417208 243098 452652 243334
rect 452888 243098 452972 243334
rect 453208 243098 488652 243334
rect 488888 243098 488972 243334
rect 489208 243098 524652 243334
rect 524888 243098 524972 243334
rect 525208 243098 560652 243334
rect 560888 243098 560972 243334
rect 561208 243098 570292 243334
rect 570528 243098 570612 243334
rect 570848 243098 585342 243334
rect 585578 243098 585662 243334
rect 585898 243098 586890 243334
rect -2966 243066 586890 243098
rect -8726 234814 592650 234846
rect -8726 234578 -8694 234814
rect -8458 234578 -8374 234814
rect -8138 234578 592062 234814
rect 592298 234578 592382 234814
rect 592618 234578 592650 234814
rect -8726 234494 592650 234578
rect -8726 234258 -8694 234494
rect -8458 234258 -8374 234494
rect -8138 234258 592062 234494
rect 592298 234258 592382 234494
rect 592618 234258 592650 234494
rect -8726 234226 592650 234258
rect -6806 231094 590730 231126
rect -6806 230858 -6774 231094
rect -6538 230858 -6454 231094
rect -6218 230858 590142 231094
rect 590378 230858 590462 231094
rect 590698 230858 590730 231094
rect -6806 230774 590730 230858
rect -6806 230538 -6774 230774
rect -6538 230538 -6454 230774
rect -6218 230538 590142 230774
rect 590378 230538 590462 230774
rect 590698 230538 590730 230774
rect -6806 230506 590730 230538
rect -4886 227374 588810 227406
rect -4886 227138 -4854 227374
rect -4618 227138 -4534 227374
rect -4298 227138 588222 227374
rect 588458 227138 588542 227374
rect 588778 227138 588810 227374
rect -4886 227054 588810 227138
rect -4886 226818 -4854 227054
rect -4618 226818 -4534 227054
rect -4298 226818 588222 227054
rect 588458 226818 588542 227054
rect 588778 226818 588810 227054
rect -4886 226786 588810 226818
rect -2966 223654 586890 223686
rect -2966 223418 -2934 223654
rect -2698 223418 -2614 223654
rect -2378 223418 7876 223654
rect 8112 223418 8196 223654
rect 8432 223418 38032 223654
rect 38268 223418 38352 223654
rect 38588 223418 74032 223654
rect 74268 223418 74352 223654
rect 74588 223418 110032 223654
rect 110268 223418 110352 223654
rect 110588 223418 146032 223654
rect 146268 223418 146352 223654
rect 146588 223418 182032 223654
rect 182268 223418 182352 223654
rect 182588 223418 218032 223654
rect 218268 223418 218352 223654
rect 218588 223418 254032 223654
rect 254268 223418 254352 223654
rect 254588 223418 290032 223654
rect 290268 223418 290352 223654
rect 290588 223418 326032 223654
rect 326268 223418 326352 223654
rect 326588 223418 362032 223654
rect 362268 223418 362352 223654
rect 362588 223418 398032 223654
rect 398268 223418 398352 223654
rect 398588 223418 434032 223654
rect 434268 223418 434352 223654
rect 434588 223418 470032 223654
rect 470268 223418 470352 223654
rect 470588 223418 506032 223654
rect 506268 223418 506352 223654
rect 506588 223418 542032 223654
rect 542268 223418 542352 223654
rect 542588 223418 571532 223654
rect 571768 223418 571852 223654
rect 572088 223418 586302 223654
rect 586538 223418 586622 223654
rect 586858 223418 586890 223654
rect -2966 223334 586890 223418
rect -2966 223098 -2934 223334
rect -2698 223098 -2614 223334
rect -2378 223098 7876 223334
rect 8112 223098 8196 223334
rect 8432 223098 38032 223334
rect 38268 223098 38352 223334
rect 38588 223098 74032 223334
rect 74268 223098 74352 223334
rect 74588 223098 110032 223334
rect 110268 223098 110352 223334
rect 110588 223098 146032 223334
rect 146268 223098 146352 223334
rect 146588 223098 182032 223334
rect 182268 223098 182352 223334
rect 182588 223098 218032 223334
rect 218268 223098 218352 223334
rect 218588 223098 254032 223334
rect 254268 223098 254352 223334
rect 254588 223098 290032 223334
rect 290268 223098 290352 223334
rect 290588 223098 326032 223334
rect 326268 223098 326352 223334
rect 326588 223098 362032 223334
rect 362268 223098 362352 223334
rect 362588 223098 398032 223334
rect 398268 223098 398352 223334
rect 398588 223098 434032 223334
rect 434268 223098 434352 223334
rect 434588 223098 470032 223334
rect 470268 223098 470352 223334
rect 470588 223098 506032 223334
rect 506268 223098 506352 223334
rect 506588 223098 542032 223334
rect 542268 223098 542352 223334
rect 542588 223098 571532 223334
rect 571768 223098 571852 223334
rect 572088 223098 586302 223334
rect 586538 223098 586622 223334
rect 586858 223098 586890 223334
rect -2966 223066 586890 223098
rect -8726 214814 592650 214846
rect -8726 214578 -7734 214814
rect -7498 214578 -7414 214814
rect -7178 214578 591102 214814
rect 591338 214578 591422 214814
rect 591658 214578 592650 214814
rect -8726 214494 592650 214578
rect -8726 214258 -7734 214494
rect -7498 214258 -7414 214494
rect -7178 214258 591102 214494
rect 591338 214258 591422 214494
rect 591658 214258 592650 214494
rect -8726 214226 592650 214258
rect -6806 211094 590730 211126
rect -6806 210858 -5814 211094
rect -5578 210858 -5494 211094
rect -5258 210858 589182 211094
rect 589418 210858 589502 211094
rect 589738 210858 590730 211094
rect -6806 210774 590730 210858
rect -6806 210538 -5814 210774
rect -5578 210538 -5494 210774
rect -5258 210538 589182 210774
rect 589418 210538 589502 210774
rect 589738 210538 590730 210774
rect -6806 210506 590730 210538
rect -4886 207374 588810 207406
rect -4886 207138 -3894 207374
rect -3658 207138 -3574 207374
rect -3338 207138 587262 207374
rect 587498 207138 587582 207374
rect 587818 207138 588810 207374
rect -4886 207054 588810 207138
rect -4886 206818 -3894 207054
rect -3658 206818 -3574 207054
rect -3338 206818 587262 207054
rect 587498 206818 587582 207054
rect 587818 206818 588810 207054
rect -4886 206786 588810 206818
rect -2966 203654 586890 203686
rect -2966 203418 -1974 203654
rect -1738 203418 -1654 203654
rect -1418 203418 9116 203654
rect 9352 203418 9436 203654
rect 9672 203418 56652 203654
rect 56888 203418 56972 203654
rect 57208 203418 92652 203654
rect 92888 203418 92972 203654
rect 93208 203418 128652 203654
rect 128888 203418 128972 203654
rect 129208 203418 164652 203654
rect 164888 203418 164972 203654
rect 165208 203418 200652 203654
rect 200888 203418 200972 203654
rect 201208 203418 236652 203654
rect 236888 203418 236972 203654
rect 237208 203418 272652 203654
rect 272888 203418 272972 203654
rect 273208 203418 308652 203654
rect 308888 203418 308972 203654
rect 309208 203418 344652 203654
rect 344888 203418 344972 203654
rect 345208 203418 380652 203654
rect 380888 203418 380972 203654
rect 381208 203418 416652 203654
rect 416888 203418 416972 203654
rect 417208 203418 452652 203654
rect 452888 203418 452972 203654
rect 453208 203418 488652 203654
rect 488888 203418 488972 203654
rect 489208 203418 524652 203654
rect 524888 203418 524972 203654
rect 525208 203418 560652 203654
rect 560888 203418 560972 203654
rect 561208 203418 570292 203654
rect 570528 203418 570612 203654
rect 570848 203418 585342 203654
rect 585578 203418 585662 203654
rect 585898 203418 586890 203654
rect -2966 203334 586890 203418
rect -2966 203098 -1974 203334
rect -1738 203098 -1654 203334
rect -1418 203098 9116 203334
rect 9352 203098 9436 203334
rect 9672 203098 56652 203334
rect 56888 203098 56972 203334
rect 57208 203098 92652 203334
rect 92888 203098 92972 203334
rect 93208 203098 128652 203334
rect 128888 203098 128972 203334
rect 129208 203098 164652 203334
rect 164888 203098 164972 203334
rect 165208 203098 200652 203334
rect 200888 203098 200972 203334
rect 201208 203098 236652 203334
rect 236888 203098 236972 203334
rect 237208 203098 272652 203334
rect 272888 203098 272972 203334
rect 273208 203098 308652 203334
rect 308888 203098 308972 203334
rect 309208 203098 344652 203334
rect 344888 203098 344972 203334
rect 345208 203098 380652 203334
rect 380888 203098 380972 203334
rect 381208 203098 416652 203334
rect 416888 203098 416972 203334
rect 417208 203098 452652 203334
rect 452888 203098 452972 203334
rect 453208 203098 488652 203334
rect 488888 203098 488972 203334
rect 489208 203098 524652 203334
rect 524888 203098 524972 203334
rect 525208 203098 560652 203334
rect 560888 203098 560972 203334
rect 561208 203098 570292 203334
rect 570528 203098 570612 203334
rect 570848 203098 585342 203334
rect 585578 203098 585662 203334
rect 585898 203098 586890 203334
rect -2966 203066 586890 203098
rect -8726 194814 592650 194846
rect -8726 194578 -8694 194814
rect -8458 194578 -8374 194814
rect -8138 194578 592062 194814
rect 592298 194578 592382 194814
rect 592618 194578 592650 194814
rect -8726 194494 592650 194578
rect -8726 194258 -8694 194494
rect -8458 194258 -8374 194494
rect -8138 194258 592062 194494
rect 592298 194258 592382 194494
rect 592618 194258 592650 194494
rect -8726 194226 592650 194258
rect -6806 191094 590730 191126
rect -6806 190858 -6774 191094
rect -6538 190858 -6454 191094
rect -6218 190858 590142 191094
rect 590378 190858 590462 191094
rect 590698 190858 590730 191094
rect -6806 190774 590730 190858
rect -6806 190538 -6774 190774
rect -6538 190538 -6454 190774
rect -6218 190538 590142 190774
rect 590378 190538 590462 190774
rect 590698 190538 590730 190774
rect -6806 190506 590730 190538
rect -4886 187374 588810 187406
rect -4886 187138 -4854 187374
rect -4618 187138 -4534 187374
rect -4298 187138 588222 187374
rect 588458 187138 588542 187374
rect 588778 187138 588810 187374
rect -4886 187054 588810 187138
rect -4886 186818 -4854 187054
rect -4618 186818 -4534 187054
rect -4298 186818 588222 187054
rect 588458 186818 588542 187054
rect 588778 186818 588810 187054
rect -4886 186786 588810 186818
rect -2966 183654 586890 183686
rect -2966 183418 -2934 183654
rect -2698 183418 -2614 183654
rect -2378 183418 7876 183654
rect 8112 183418 8196 183654
rect 8432 183418 38032 183654
rect 38268 183418 38352 183654
rect 38588 183418 60622 183654
rect 60858 183418 159098 183654
rect 159334 183418 182032 183654
rect 182268 183418 182352 183654
rect 182588 183418 185622 183654
rect 185858 183418 284098 183654
rect 284334 183418 290032 183654
rect 290268 183418 290352 183654
rect 290588 183418 310622 183654
rect 310858 183418 409098 183654
rect 409334 183418 434032 183654
rect 434268 183418 434352 183654
rect 434588 183418 436622 183654
rect 436858 183418 535098 183654
rect 535334 183418 542032 183654
rect 542268 183418 542352 183654
rect 542588 183418 571532 183654
rect 571768 183418 571852 183654
rect 572088 183418 586302 183654
rect 586538 183418 586622 183654
rect 586858 183418 586890 183654
rect -2966 183334 586890 183418
rect -2966 183098 -2934 183334
rect -2698 183098 -2614 183334
rect -2378 183098 7876 183334
rect 8112 183098 8196 183334
rect 8432 183098 38032 183334
rect 38268 183098 38352 183334
rect 38588 183098 60622 183334
rect 60858 183098 159098 183334
rect 159334 183098 182032 183334
rect 182268 183098 182352 183334
rect 182588 183098 185622 183334
rect 185858 183098 284098 183334
rect 284334 183098 290032 183334
rect 290268 183098 290352 183334
rect 290588 183098 310622 183334
rect 310858 183098 409098 183334
rect 409334 183098 434032 183334
rect 434268 183098 434352 183334
rect 434588 183098 436622 183334
rect 436858 183098 535098 183334
rect 535334 183098 542032 183334
rect 542268 183098 542352 183334
rect 542588 183098 571532 183334
rect 571768 183098 571852 183334
rect 572088 183098 586302 183334
rect 586538 183098 586622 183334
rect 586858 183098 586890 183334
rect -2966 183066 586890 183098
rect -8726 174814 592650 174846
rect -8726 174578 -7734 174814
rect -7498 174578 -7414 174814
rect -7178 174578 591102 174814
rect 591338 174578 591422 174814
rect 591658 174578 592650 174814
rect -8726 174494 592650 174578
rect -8726 174258 -7734 174494
rect -7498 174258 -7414 174494
rect -7178 174258 591102 174494
rect 591338 174258 591422 174494
rect 591658 174258 592650 174494
rect -8726 174226 592650 174258
rect -6806 171094 590730 171126
rect -6806 170858 -5814 171094
rect -5578 170858 -5494 171094
rect -5258 170858 589182 171094
rect 589418 170858 589502 171094
rect 589738 170858 590730 171094
rect -6806 170774 590730 170858
rect -6806 170538 -5814 170774
rect -5578 170538 -5494 170774
rect -5258 170538 589182 170774
rect 589418 170538 589502 170774
rect 589738 170538 590730 170774
rect -6806 170506 590730 170538
rect -4886 167374 588810 167406
rect -4886 167138 -3894 167374
rect -3658 167138 -3574 167374
rect -3338 167138 587262 167374
rect 587498 167138 587582 167374
rect 587818 167138 588810 167374
rect -4886 167054 588810 167138
rect -4886 166818 -3894 167054
rect -3658 166818 -3574 167054
rect -3338 166818 587262 167054
rect 587498 166818 587582 167054
rect 587818 166818 588810 167054
rect -4886 166786 588810 166818
rect -2966 163654 586890 163686
rect -2966 163418 -1974 163654
rect -1738 163418 -1654 163654
rect -1418 163418 9116 163654
rect 9352 163418 9436 163654
rect 9672 163418 56652 163654
rect 56888 163418 56972 163654
rect 57208 163418 61342 163654
rect 61578 163418 158378 163654
rect 158614 163418 164652 163654
rect 164888 163418 164972 163654
rect 165208 163418 186342 163654
rect 186578 163418 283378 163654
rect 283614 163418 308652 163654
rect 308888 163418 308972 163654
rect 309208 163418 311342 163654
rect 311578 163418 408378 163654
rect 408614 163418 416652 163654
rect 416888 163418 416972 163654
rect 417208 163418 437342 163654
rect 437578 163418 534378 163654
rect 534614 163418 560652 163654
rect 560888 163418 560972 163654
rect 561208 163418 570292 163654
rect 570528 163418 570612 163654
rect 570848 163418 585342 163654
rect 585578 163418 585662 163654
rect 585898 163418 586890 163654
rect -2966 163334 586890 163418
rect -2966 163098 -1974 163334
rect -1738 163098 -1654 163334
rect -1418 163098 9116 163334
rect 9352 163098 9436 163334
rect 9672 163098 56652 163334
rect 56888 163098 56972 163334
rect 57208 163098 61342 163334
rect 61578 163098 158378 163334
rect 158614 163098 164652 163334
rect 164888 163098 164972 163334
rect 165208 163098 186342 163334
rect 186578 163098 283378 163334
rect 283614 163098 308652 163334
rect 308888 163098 308972 163334
rect 309208 163098 311342 163334
rect 311578 163098 408378 163334
rect 408614 163098 416652 163334
rect 416888 163098 416972 163334
rect 417208 163098 437342 163334
rect 437578 163098 534378 163334
rect 534614 163098 560652 163334
rect 560888 163098 560972 163334
rect 561208 163098 570292 163334
rect 570528 163098 570612 163334
rect 570848 163098 585342 163334
rect 585578 163098 585662 163334
rect 585898 163098 586890 163334
rect -2966 163066 586890 163098
rect -8726 154814 592650 154846
rect -8726 154578 -8694 154814
rect -8458 154578 -8374 154814
rect -8138 154578 592062 154814
rect 592298 154578 592382 154814
rect 592618 154578 592650 154814
rect -8726 154494 592650 154578
rect -8726 154258 -8694 154494
rect -8458 154258 -8374 154494
rect -8138 154258 592062 154494
rect 592298 154258 592382 154494
rect 592618 154258 592650 154494
rect -8726 154226 592650 154258
rect -6806 151094 590730 151126
rect -6806 150858 -6774 151094
rect -6538 150858 -6454 151094
rect -6218 150858 590142 151094
rect 590378 150858 590462 151094
rect 590698 150858 590730 151094
rect -6806 150774 590730 150858
rect -6806 150538 -6774 150774
rect -6538 150538 -6454 150774
rect -6218 150538 590142 150774
rect 590378 150538 590462 150774
rect 590698 150538 590730 150774
rect -6806 150506 590730 150538
rect -4886 147374 588810 147406
rect -4886 147138 -4854 147374
rect -4618 147138 -4534 147374
rect -4298 147138 588222 147374
rect 588458 147138 588542 147374
rect 588778 147138 588810 147374
rect -4886 147054 588810 147138
rect -4886 146818 -4854 147054
rect -4618 146818 -4534 147054
rect -4298 146818 588222 147054
rect 588458 146818 588542 147054
rect 588778 146818 588810 147054
rect -4886 146786 588810 146818
rect -2966 143654 586890 143686
rect -2966 143418 -2934 143654
rect -2698 143418 -2614 143654
rect -2378 143418 7876 143654
rect 8112 143418 8196 143654
rect 8432 143418 38032 143654
rect 38268 143418 38352 143654
rect 38588 143418 60622 143654
rect 60858 143418 159098 143654
rect 159334 143418 182032 143654
rect 182268 143418 182352 143654
rect 182588 143418 185622 143654
rect 185858 143418 284098 143654
rect 284334 143418 290032 143654
rect 290268 143418 290352 143654
rect 290588 143418 310622 143654
rect 310858 143418 409098 143654
rect 409334 143418 434032 143654
rect 434268 143418 434352 143654
rect 434588 143418 436622 143654
rect 436858 143418 535098 143654
rect 535334 143418 542032 143654
rect 542268 143418 542352 143654
rect 542588 143418 571532 143654
rect 571768 143418 571852 143654
rect 572088 143418 586302 143654
rect 586538 143418 586622 143654
rect 586858 143418 586890 143654
rect -2966 143334 586890 143418
rect -2966 143098 -2934 143334
rect -2698 143098 -2614 143334
rect -2378 143098 7876 143334
rect 8112 143098 8196 143334
rect 8432 143098 38032 143334
rect 38268 143098 38352 143334
rect 38588 143098 60622 143334
rect 60858 143098 159098 143334
rect 159334 143098 182032 143334
rect 182268 143098 182352 143334
rect 182588 143098 185622 143334
rect 185858 143098 284098 143334
rect 284334 143098 290032 143334
rect 290268 143098 290352 143334
rect 290588 143098 310622 143334
rect 310858 143098 409098 143334
rect 409334 143098 434032 143334
rect 434268 143098 434352 143334
rect 434588 143098 436622 143334
rect 436858 143098 535098 143334
rect 535334 143098 542032 143334
rect 542268 143098 542352 143334
rect 542588 143098 571532 143334
rect 571768 143098 571852 143334
rect 572088 143098 586302 143334
rect 586538 143098 586622 143334
rect 586858 143098 586890 143334
rect -2966 143066 586890 143098
rect -8726 134814 592650 134846
rect -8726 134578 -7734 134814
rect -7498 134578 -7414 134814
rect -7178 134578 591102 134814
rect 591338 134578 591422 134814
rect 591658 134578 592650 134814
rect -8726 134494 592650 134578
rect -8726 134258 -7734 134494
rect -7498 134258 -7414 134494
rect -7178 134258 591102 134494
rect 591338 134258 591422 134494
rect 591658 134258 592650 134494
rect -8726 134226 592650 134258
rect -6806 131094 590730 131126
rect -6806 130858 -5814 131094
rect -5578 130858 -5494 131094
rect -5258 130858 589182 131094
rect 589418 130858 589502 131094
rect 589738 130858 590730 131094
rect -6806 130774 590730 130858
rect -6806 130538 -5814 130774
rect -5578 130538 -5494 130774
rect -5258 130538 589182 130774
rect 589418 130538 589502 130774
rect 589738 130538 590730 130774
rect -6806 130506 590730 130538
rect -4886 127374 588810 127406
rect -4886 127138 -3894 127374
rect -3658 127138 -3574 127374
rect -3338 127138 587262 127374
rect 587498 127138 587582 127374
rect 587818 127138 588810 127374
rect -4886 127054 588810 127138
rect -4886 126818 -3894 127054
rect -3658 126818 -3574 127054
rect -3338 126818 587262 127054
rect 587498 126818 587582 127054
rect 587818 126818 588810 127054
rect -4886 126786 588810 126818
rect -2966 123654 586890 123686
rect -2966 123418 -1974 123654
rect -1738 123418 -1654 123654
rect -1418 123418 9116 123654
rect 9352 123418 9436 123654
rect 9672 123418 56652 123654
rect 56888 123418 56972 123654
rect 57208 123418 61342 123654
rect 61578 123418 158378 123654
rect 158614 123418 164652 123654
rect 164888 123418 164972 123654
rect 165208 123418 186342 123654
rect 186578 123418 283378 123654
rect 283614 123418 308652 123654
rect 308888 123418 308972 123654
rect 309208 123418 311342 123654
rect 311578 123418 408378 123654
rect 408614 123418 416652 123654
rect 416888 123418 416972 123654
rect 417208 123418 437342 123654
rect 437578 123418 534378 123654
rect 534614 123418 560652 123654
rect 560888 123418 560972 123654
rect 561208 123418 570292 123654
rect 570528 123418 570612 123654
rect 570848 123418 585342 123654
rect 585578 123418 585662 123654
rect 585898 123418 586890 123654
rect -2966 123334 586890 123418
rect -2966 123098 -1974 123334
rect -1738 123098 -1654 123334
rect -1418 123098 9116 123334
rect 9352 123098 9436 123334
rect 9672 123098 56652 123334
rect 56888 123098 56972 123334
rect 57208 123098 61342 123334
rect 61578 123098 158378 123334
rect 158614 123098 164652 123334
rect 164888 123098 164972 123334
rect 165208 123098 186342 123334
rect 186578 123098 283378 123334
rect 283614 123098 308652 123334
rect 308888 123098 308972 123334
rect 309208 123098 311342 123334
rect 311578 123098 408378 123334
rect 408614 123098 416652 123334
rect 416888 123098 416972 123334
rect 417208 123098 437342 123334
rect 437578 123098 534378 123334
rect 534614 123098 560652 123334
rect 560888 123098 560972 123334
rect 561208 123098 570292 123334
rect 570528 123098 570612 123334
rect 570848 123098 585342 123334
rect 585578 123098 585662 123334
rect 585898 123098 586890 123334
rect -2966 123066 586890 123098
rect -8726 114814 592650 114846
rect -8726 114578 -8694 114814
rect -8458 114578 -8374 114814
rect -8138 114578 592062 114814
rect 592298 114578 592382 114814
rect 592618 114578 592650 114814
rect -8726 114494 592650 114578
rect -8726 114258 -8694 114494
rect -8458 114258 -8374 114494
rect -8138 114258 592062 114494
rect 592298 114258 592382 114494
rect 592618 114258 592650 114494
rect -8726 114226 592650 114258
rect -6806 111094 590730 111126
rect -6806 110858 -6774 111094
rect -6538 110858 -6454 111094
rect -6218 110858 590142 111094
rect 590378 110858 590462 111094
rect 590698 110858 590730 111094
rect -6806 110774 590730 110858
rect -6806 110538 -6774 110774
rect -6538 110538 -6454 110774
rect -6218 110538 590142 110774
rect 590378 110538 590462 110774
rect 590698 110538 590730 110774
rect -6806 110506 590730 110538
rect -4886 107374 588810 107406
rect -4886 107138 -4854 107374
rect -4618 107138 -4534 107374
rect -4298 107138 588222 107374
rect 588458 107138 588542 107374
rect 588778 107138 588810 107374
rect -4886 107054 588810 107138
rect -4886 106818 -4854 107054
rect -4618 106818 -4534 107054
rect -4298 106818 588222 107054
rect 588458 106818 588542 107054
rect 588778 106818 588810 107054
rect -4886 106786 588810 106818
rect -2966 103654 586890 103686
rect -2966 103418 -2934 103654
rect -2698 103418 -2614 103654
rect -2378 103418 7876 103654
rect 8112 103418 8196 103654
rect 8432 103418 38032 103654
rect 38268 103418 38352 103654
rect 38588 103418 74032 103654
rect 74268 103418 74352 103654
rect 74588 103418 110032 103654
rect 110268 103418 110352 103654
rect 110588 103418 146032 103654
rect 146268 103418 146352 103654
rect 146588 103418 182032 103654
rect 182268 103418 182352 103654
rect 182588 103418 218032 103654
rect 218268 103418 218352 103654
rect 218588 103418 254032 103654
rect 254268 103418 254352 103654
rect 254588 103418 290032 103654
rect 290268 103418 290352 103654
rect 290588 103418 326032 103654
rect 326268 103418 326352 103654
rect 326588 103418 362032 103654
rect 362268 103418 362352 103654
rect 362588 103418 398032 103654
rect 398268 103418 398352 103654
rect 398588 103418 434032 103654
rect 434268 103418 434352 103654
rect 434588 103418 470032 103654
rect 470268 103418 470352 103654
rect 470588 103418 506032 103654
rect 506268 103418 506352 103654
rect 506588 103418 542032 103654
rect 542268 103418 542352 103654
rect 542588 103418 571532 103654
rect 571768 103418 571852 103654
rect 572088 103418 586302 103654
rect 586538 103418 586622 103654
rect 586858 103418 586890 103654
rect -2966 103334 586890 103418
rect -2966 103098 -2934 103334
rect -2698 103098 -2614 103334
rect -2378 103098 7876 103334
rect 8112 103098 8196 103334
rect 8432 103098 38032 103334
rect 38268 103098 38352 103334
rect 38588 103098 74032 103334
rect 74268 103098 74352 103334
rect 74588 103098 110032 103334
rect 110268 103098 110352 103334
rect 110588 103098 146032 103334
rect 146268 103098 146352 103334
rect 146588 103098 182032 103334
rect 182268 103098 182352 103334
rect 182588 103098 218032 103334
rect 218268 103098 218352 103334
rect 218588 103098 254032 103334
rect 254268 103098 254352 103334
rect 254588 103098 290032 103334
rect 290268 103098 290352 103334
rect 290588 103098 326032 103334
rect 326268 103098 326352 103334
rect 326588 103098 362032 103334
rect 362268 103098 362352 103334
rect 362588 103098 398032 103334
rect 398268 103098 398352 103334
rect 398588 103098 434032 103334
rect 434268 103098 434352 103334
rect 434588 103098 470032 103334
rect 470268 103098 470352 103334
rect 470588 103098 506032 103334
rect 506268 103098 506352 103334
rect 506588 103098 542032 103334
rect 542268 103098 542352 103334
rect 542588 103098 571532 103334
rect 571768 103098 571852 103334
rect 572088 103098 586302 103334
rect 586538 103098 586622 103334
rect 586858 103098 586890 103334
rect -2966 103066 586890 103098
rect -8726 94814 592650 94846
rect -8726 94578 -7734 94814
rect -7498 94578 -7414 94814
rect -7178 94578 591102 94814
rect 591338 94578 591422 94814
rect 591658 94578 592650 94814
rect -8726 94494 592650 94578
rect -8726 94258 -7734 94494
rect -7498 94258 -7414 94494
rect -7178 94258 591102 94494
rect 591338 94258 591422 94494
rect 591658 94258 592650 94494
rect -8726 94226 592650 94258
rect -6806 91094 590730 91126
rect -6806 90858 -5814 91094
rect -5578 90858 -5494 91094
rect -5258 90858 589182 91094
rect 589418 90858 589502 91094
rect 589738 90858 590730 91094
rect -6806 90774 590730 90858
rect -6806 90538 -5814 90774
rect -5578 90538 -5494 90774
rect -5258 90538 589182 90774
rect 589418 90538 589502 90774
rect 589738 90538 590730 90774
rect -6806 90506 590730 90538
rect -4886 87374 588810 87406
rect -4886 87138 -3894 87374
rect -3658 87138 -3574 87374
rect -3338 87138 587262 87374
rect 587498 87138 587582 87374
rect 587818 87138 588810 87374
rect -4886 87054 588810 87138
rect -4886 86818 -3894 87054
rect -3658 86818 -3574 87054
rect -3338 86818 587262 87054
rect 587498 86818 587582 87054
rect 587818 86818 588810 87054
rect -4886 86786 588810 86818
rect -2966 83654 586890 83686
rect -2966 83418 -1974 83654
rect -1738 83418 -1654 83654
rect -1418 83418 9116 83654
rect 9352 83418 9436 83654
rect 9672 83418 56652 83654
rect 56888 83418 56972 83654
rect 57208 83418 61342 83654
rect 61578 83418 158378 83654
rect 158614 83418 164652 83654
rect 164888 83418 164972 83654
rect 165208 83418 186342 83654
rect 186578 83418 283378 83654
rect 283614 83418 308652 83654
rect 308888 83418 308972 83654
rect 309208 83418 311342 83654
rect 311578 83418 408378 83654
rect 408614 83418 416652 83654
rect 416888 83418 416972 83654
rect 417208 83418 437342 83654
rect 437578 83418 534378 83654
rect 534614 83418 560652 83654
rect 560888 83418 560972 83654
rect 561208 83418 570292 83654
rect 570528 83418 570612 83654
rect 570848 83418 585342 83654
rect 585578 83418 585662 83654
rect 585898 83418 586890 83654
rect -2966 83334 586890 83418
rect -2966 83098 -1974 83334
rect -1738 83098 -1654 83334
rect -1418 83098 9116 83334
rect 9352 83098 9436 83334
rect 9672 83098 56652 83334
rect 56888 83098 56972 83334
rect 57208 83098 61342 83334
rect 61578 83098 158378 83334
rect 158614 83098 164652 83334
rect 164888 83098 164972 83334
rect 165208 83098 186342 83334
rect 186578 83098 283378 83334
rect 283614 83098 308652 83334
rect 308888 83098 308972 83334
rect 309208 83098 311342 83334
rect 311578 83098 408378 83334
rect 408614 83098 416652 83334
rect 416888 83098 416972 83334
rect 417208 83098 437342 83334
rect 437578 83098 534378 83334
rect 534614 83098 560652 83334
rect 560888 83098 560972 83334
rect 561208 83098 570292 83334
rect 570528 83098 570612 83334
rect 570848 83098 585342 83334
rect 585578 83098 585662 83334
rect 585898 83098 586890 83334
rect -2966 83066 586890 83098
rect -8726 74814 592650 74846
rect -8726 74578 -8694 74814
rect -8458 74578 -8374 74814
rect -8138 74578 592062 74814
rect 592298 74578 592382 74814
rect 592618 74578 592650 74814
rect -8726 74494 592650 74578
rect -8726 74258 -8694 74494
rect -8458 74258 -8374 74494
rect -8138 74258 592062 74494
rect 592298 74258 592382 74494
rect 592618 74258 592650 74494
rect -8726 74226 592650 74258
rect -6806 71094 590730 71126
rect -6806 70858 -6774 71094
rect -6538 70858 -6454 71094
rect -6218 70858 590142 71094
rect 590378 70858 590462 71094
rect 590698 70858 590730 71094
rect -6806 70774 590730 70858
rect -6806 70538 -6774 70774
rect -6538 70538 -6454 70774
rect -6218 70538 590142 70774
rect 590378 70538 590462 70774
rect 590698 70538 590730 70774
rect -6806 70506 590730 70538
rect -4886 67374 588810 67406
rect -4886 67138 -4854 67374
rect -4618 67138 -4534 67374
rect -4298 67138 588222 67374
rect 588458 67138 588542 67374
rect 588778 67138 588810 67374
rect -4886 67054 588810 67138
rect -4886 66818 -4854 67054
rect -4618 66818 -4534 67054
rect -4298 66818 588222 67054
rect 588458 66818 588542 67054
rect 588778 66818 588810 67054
rect -4886 66786 588810 66818
rect -2966 63654 586890 63686
rect -2966 63418 -2934 63654
rect -2698 63418 -2614 63654
rect -2378 63418 7876 63654
rect 8112 63418 8196 63654
rect 8432 63418 38032 63654
rect 38268 63418 38352 63654
rect 38588 63418 60622 63654
rect 60858 63418 159098 63654
rect 159334 63418 182032 63654
rect 182268 63418 182352 63654
rect 182588 63418 185622 63654
rect 185858 63418 284098 63654
rect 284334 63418 290032 63654
rect 290268 63418 290352 63654
rect 290588 63418 310622 63654
rect 310858 63418 409098 63654
rect 409334 63418 434032 63654
rect 434268 63418 434352 63654
rect 434588 63418 436622 63654
rect 436858 63418 535098 63654
rect 535334 63418 542032 63654
rect 542268 63418 542352 63654
rect 542588 63418 571532 63654
rect 571768 63418 571852 63654
rect 572088 63418 586302 63654
rect 586538 63418 586622 63654
rect 586858 63418 586890 63654
rect -2966 63334 586890 63418
rect -2966 63098 -2934 63334
rect -2698 63098 -2614 63334
rect -2378 63098 7876 63334
rect 8112 63098 8196 63334
rect 8432 63098 38032 63334
rect 38268 63098 38352 63334
rect 38588 63098 60622 63334
rect 60858 63098 159098 63334
rect 159334 63098 182032 63334
rect 182268 63098 182352 63334
rect 182588 63098 185622 63334
rect 185858 63098 284098 63334
rect 284334 63098 290032 63334
rect 290268 63098 290352 63334
rect 290588 63098 310622 63334
rect 310858 63098 409098 63334
rect 409334 63098 434032 63334
rect 434268 63098 434352 63334
rect 434588 63098 436622 63334
rect 436858 63098 535098 63334
rect 535334 63098 542032 63334
rect 542268 63098 542352 63334
rect 542588 63098 571532 63334
rect 571768 63098 571852 63334
rect 572088 63098 586302 63334
rect 586538 63098 586622 63334
rect 586858 63098 586890 63334
rect -2966 63066 586890 63098
rect -8726 54814 592650 54846
rect -8726 54578 -7734 54814
rect -7498 54578 -7414 54814
rect -7178 54578 591102 54814
rect 591338 54578 591422 54814
rect 591658 54578 592650 54814
rect -8726 54494 592650 54578
rect -8726 54258 -7734 54494
rect -7498 54258 -7414 54494
rect -7178 54258 591102 54494
rect 591338 54258 591422 54494
rect 591658 54258 592650 54494
rect -8726 54226 592650 54258
rect -6806 51094 590730 51126
rect -6806 50858 -5814 51094
rect -5578 50858 -5494 51094
rect -5258 50858 589182 51094
rect 589418 50858 589502 51094
rect 589738 50858 590730 51094
rect -6806 50774 590730 50858
rect -6806 50538 -5814 50774
rect -5578 50538 -5494 50774
rect -5258 50538 589182 50774
rect 589418 50538 589502 50774
rect 589738 50538 590730 50774
rect -6806 50506 590730 50538
rect -4886 47374 588810 47406
rect -4886 47138 -3894 47374
rect -3658 47138 -3574 47374
rect -3338 47138 587262 47374
rect 587498 47138 587582 47374
rect 587818 47138 588810 47374
rect -4886 47054 588810 47138
rect -4886 46818 -3894 47054
rect -3658 46818 -3574 47054
rect -3338 46818 587262 47054
rect 587498 46818 587582 47054
rect 587818 46818 588810 47054
rect -4886 46786 588810 46818
rect -2966 43654 586890 43686
rect -2966 43418 -1974 43654
rect -1738 43418 -1654 43654
rect -1418 43418 9116 43654
rect 9352 43418 9436 43654
rect 9672 43418 56652 43654
rect 56888 43418 56972 43654
rect 57208 43418 61342 43654
rect 61578 43418 158378 43654
rect 158614 43418 164652 43654
rect 164888 43418 164972 43654
rect 165208 43418 186342 43654
rect 186578 43418 283378 43654
rect 283614 43418 308652 43654
rect 308888 43418 308972 43654
rect 309208 43418 311342 43654
rect 311578 43418 408378 43654
rect 408614 43418 416652 43654
rect 416888 43418 416972 43654
rect 417208 43418 437342 43654
rect 437578 43418 534378 43654
rect 534614 43418 560652 43654
rect 560888 43418 560972 43654
rect 561208 43418 570292 43654
rect 570528 43418 570612 43654
rect 570848 43418 585342 43654
rect 585578 43418 585662 43654
rect 585898 43418 586890 43654
rect -2966 43334 586890 43418
rect -2966 43098 -1974 43334
rect -1738 43098 -1654 43334
rect -1418 43098 9116 43334
rect 9352 43098 9436 43334
rect 9672 43098 56652 43334
rect 56888 43098 56972 43334
rect 57208 43098 61342 43334
rect 61578 43098 158378 43334
rect 158614 43098 164652 43334
rect 164888 43098 164972 43334
rect 165208 43098 186342 43334
rect 186578 43098 283378 43334
rect 283614 43098 308652 43334
rect 308888 43098 308972 43334
rect 309208 43098 311342 43334
rect 311578 43098 408378 43334
rect 408614 43098 416652 43334
rect 416888 43098 416972 43334
rect 417208 43098 437342 43334
rect 437578 43098 534378 43334
rect 534614 43098 560652 43334
rect 560888 43098 560972 43334
rect 561208 43098 570292 43334
rect 570528 43098 570612 43334
rect 570848 43098 585342 43334
rect 585578 43098 585662 43334
rect 585898 43098 586890 43334
rect -2966 43066 586890 43098
rect -8726 34814 592650 34846
rect -8726 34578 -8694 34814
rect -8458 34578 -8374 34814
rect -8138 34578 592062 34814
rect 592298 34578 592382 34814
rect 592618 34578 592650 34814
rect -8726 34494 592650 34578
rect -8726 34258 -8694 34494
rect -8458 34258 -8374 34494
rect -8138 34258 592062 34494
rect 592298 34258 592382 34494
rect 592618 34258 592650 34494
rect -8726 34226 592650 34258
rect -6806 31094 590730 31126
rect -6806 30858 -6774 31094
rect -6538 30858 -6454 31094
rect -6218 30858 590142 31094
rect 590378 30858 590462 31094
rect 590698 30858 590730 31094
rect -6806 30774 590730 30858
rect -6806 30538 -6774 30774
rect -6538 30538 -6454 30774
rect -6218 30538 590142 30774
rect 590378 30538 590462 30774
rect 590698 30538 590730 30774
rect -6806 30506 590730 30538
rect -4886 27374 588810 27406
rect -4886 27138 -4854 27374
rect -4618 27138 -4534 27374
rect -4298 27138 588222 27374
rect 588458 27138 588542 27374
rect 588778 27138 588810 27374
rect -4886 27054 588810 27138
rect -4886 26818 -4854 27054
rect -4618 26818 -4534 27054
rect -4298 26818 588222 27054
rect 588458 26818 588542 27054
rect 588778 26818 588810 27054
rect -4886 26786 588810 26818
rect -2966 23654 586890 23686
rect -2966 23418 -2934 23654
rect -2698 23418 -2614 23654
rect -2378 23418 7876 23654
rect 8112 23418 8196 23654
rect 8432 23418 38032 23654
rect 38268 23418 38352 23654
rect 38588 23418 60622 23654
rect 60858 23418 159098 23654
rect 159334 23418 182032 23654
rect 182268 23418 182352 23654
rect 182588 23418 185622 23654
rect 185858 23418 284098 23654
rect 284334 23418 290032 23654
rect 290268 23418 290352 23654
rect 290588 23418 310622 23654
rect 310858 23418 409098 23654
rect 409334 23418 434032 23654
rect 434268 23418 434352 23654
rect 434588 23418 436622 23654
rect 436858 23418 535098 23654
rect 535334 23418 542032 23654
rect 542268 23418 542352 23654
rect 542588 23418 571532 23654
rect 571768 23418 571852 23654
rect 572088 23418 586302 23654
rect 586538 23418 586622 23654
rect 586858 23418 586890 23654
rect -2966 23334 586890 23418
rect -2966 23098 -2934 23334
rect -2698 23098 -2614 23334
rect -2378 23098 7876 23334
rect 8112 23098 8196 23334
rect 8432 23098 38032 23334
rect 38268 23098 38352 23334
rect 38588 23098 60622 23334
rect 60858 23098 159098 23334
rect 159334 23098 182032 23334
rect 182268 23098 182352 23334
rect 182588 23098 185622 23334
rect 185858 23098 284098 23334
rect 284334 23098 290032 23334
rect 290268 23098 290352 23334
rect 290588 23098 310622 23334
rect 310858 23098 409098 23334
rect 409334 23098 434032 23334
rect 434268 23098 434352 23334
rect 434588 23098 436622 23334
rect 436858 23098 535098 23334
rect 535334 23098 542032 23334
rect 542268 23098 542352 23334
rect 542588 23098 571532 23334
rect 571768 23098 571852 23334
rect 572088 23098 586302 23334
rect 586538 23098 586622 23334
rect 586858 23098 586890 23334
rect -2966 23066 586890 23098
rect -8726 14814 592650 14846
rect -8726 14578 -7734 14814
rect -7498 14578 -7414 14814
rect -7178 14578 591102 14814
rect 591338 14578 591422 14814
rect 591658 14578 592650 14814
rect -8726 14494 592650 14578
rect -8726 14258 -7734 14494
rect -7498 14258 -7414 14494
rect -7178 14258 591102 14494
rect 591338 14258 591422 14494
rect 591658 14258 592650 14494
rect -8726 14226 592650 14258
rect -6806 11094 590730 11126
rect -6806 10858 -5814 11094
rect -5578 10858 -5494 11094
rect -5258 10858 589182 11094
rect 589418 10858 589502 11094
rect 589738 10858 590730 11094
rect -6806 10774 590730 10858
rect -6806 10538 -5814 10774
rect -5578 10538 -5494 10774
rect -5258 10538 589182 10774
rect 589418 10538 589502 10774
rect 589738 10538 590730 10774
rect -6806 10506 590730 10538
rect -4886 7374 588810 7406
rect -4886 7138 -3894 7374
rect -3658 7138 -3574 7374
rect -3338 7138 587262 7374
rect 587498 7138 587582 7374
rect 587818 7138 588810 7374
rect -4886 7054 588810 7138
rect -4886 6818 -3894 7054
rect -3658 6818 -3574 7054
rect -3338 6818 587262 7054
rect 587498 6818 587582 7054
rect 587818 6818 588810 7054
rect -4886 6786 588810 6818
rect -2966 3654 586890 3686
rect -2966 3418 -1974 3654
rect -1738 3418 -1654 3654
rect -1418 3418 585342 3654
rect 585578 3418 585662 3654
rect 585898 3418 586890 3654
rect -2966 3334 586890 3418
rect -2966 3098 -1974 3334
rect -1738 3098 -1654 3334
rect -1418 3098 585342 3334
rect 585578 3098 585662 3334
rect 585898 3098 586890 3334
rect -2966 3066 586890 3098
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 2026 -346
rect 2262 -582 2346 -346
rect 2582 -582 42026 -346
rect 42262 -582 42346 -346
rect 42582 -582 82026 -346
rect 82262 -582 82346 -346
rect 82582 -582 122026 -346
rect 122262 -582 122346 -346
rect 122582 -582 162026 -346
rect 162262 -582 162346 -346
rect 162582 -582 202026 -346
rect 202262 -582 202346 -346
rect 202582 -582 242026 -346
rect 242262 -582 242346 -346
rect 242582 -582 282026 -346
rect 282262 -582 282346 -346
rect 282582 -582 322026 -346
rect 322262 -582 322346 -346
rect 322582 -582 362026 -346
rect 362262 -582 362346 -346
rect 362582 -582 402026 -346
rect 402262 -582 402346 -346
rect 402582 -582 442026 -346
rect 442262 -582 442346 -346
rect 442582 -582 482026 -346
rect 482262 -582 482346 -346
rect 482582 -582 522026 -346
rect 522262 -582 522346 -346
rect 522582 -582 562026 -346
rect 562262 -582 562346 -346
rect 562582 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 2026 -666
rect 2262 -902 2346 -666
rect 2582 -902 42026 -666
rect 42262 -902 42346 -666
rect 42582 -902 82026 -666
rect 82262 -902 82346 -666
rect 82582 -902 122026 -666
rect 122262 -902 122346 -666
rect 122582 -902 162026 -666
rect 162262 -902 162346 -666
rect 162582 -902 202026 -666
rect 202262 -902 202346 -666
rect 202582 -902 242026 -666
rect 242262 -902 242346 -666
rect 242582 -902 282026 -666
rect 282262 -902 282346 -666
rect 282582 -902 322026 -666
rect 322262 -902 322346 -666
rect 322582 -902 362026 -666
rect 362262 -902 362346 -666
rect 362582 -902 402026 -666
rect 402262 -902 402346 -666
rect 402582 -902 442026 -666
rect 442262 -902 442346 -666
rect 442582 -902 482026 -666
rect 482262 -902 482346 -666
rect 482582 -902 522026 -666
rect 522262 -902 522346 -666
rect 522582 -902 562026 -666
rect 562262 -902 562346 -666
rect 562582 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 22026 -1306
rect 22262 -1542 22346 -1306
rect 22582 -1542 62026 -1306
rect 62262 -1542 62346 -1306
rect 62582 -1542 102026 -1306
rect 102262 -1542 102346 -1306
rect 102582 -1542 142026 -1306
rect 142262 -1542 142346 -1306
rect 142582 -1542 182026 -1306
rect 182262 -1542 182346 -1306
rect 182582 -1542 222026 -1306
rect 222262 -1542 222346 -1306
rect 222582 -1542 262026 -1306
rect 262262 -1542 262346 -1306
rect 262582 -1542 302026 -1306
rect 302262 -1542 302346 -1306
rect 302582 -1542 342026 -1306
rect 342262 -1542 342346 -1306
rect 342582 -1542 382026 -1306
rect 382262 -1542 382346 -1306
rect 382582 -1542 422026 -1306
rect 422262 -1542 422346 -1306
rect 422582 -1542 462026 -1306
rect 462262 -1542 462346 -1306
rect 462582 -1542 502026 -1306
rect 502262 -1542 502346 -1306
rect 502582 -1542 542026 -1306
rect 542262 -1542 542346 -1306
rect 542582 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 22026 -1626
rect 22262 -1862 22346 -1626
rect 22582 -1862 62026 -1626
rect 62262 -1862 62346 -1626
rect 62582 -1862 102026 -1626
rect 102262 -1862 102346 -1626
rect 102582 -1862 142026 -1626
rect 142262 -1862 142346 -1626
rect 142582 -1862 182026 -1626
rect 182262 -1862 182346 -1626
rect 182582 -1862 222026 -1626
rect 222262 -1862 222346 -1626
rect 222582 -1862 262026 -1626
rect 262262 -1862 262346 -1626
rect 262582 -1862 302026 -1626
rect 302262 -1862 302346 -1626
rect 302582 -1862 342026 -1626
rect 342262 -1862 342346 -1626
rect 342582 -1862 382026 -1626
rect 382262 -1862 382346 -1626
rect 382582 -1862 422026 -1626
rect 422262 -1862 422346 -1626
rect 422582 -1862 462026 -1626
rect 462262 -1862 462346 -1626
rect 462582 -1862 502026 -1626
rect 502262 -1862 502346 -1626
rect 502582 -1862 542026 -1626
rect 542262 -1862 542346 -1626
rect 542582 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5746 -2266
rect 5982 -2502 6066 -2266
rect 6302 -2502 45746 -2266
rect 45982 -2502 46066 -2266
rect 46302 -2502 85746 -2266
rect 85982 -2502 86066 -2266
rect 86302 -2502 125746 -2266
rect 125982 -2502 126066 -2266
rect 126302 -2502 165746 -2266
rect 165982 -2502 166066 -2266
rect 166302 -2502 205746 -2266
rect 205982 -2502 206066 -2266
rect 206302 -2502 245746 -2266
rect 245982 -2502 246066 -2266
rect 246302 -2502 285746 -2266
rect 285982 -2502 286066 -2266
rect 286302 -2502 325746 -2266
rect 325982 -2502 326066 -2266
rect 326302 -2502 365746 -2266
rect 365982 -2502 366066 -2266
rect 366302 -2502 405746 -2266
rect 405982 -2502 406066 -2266
rect 406302 -2502 445746 -2266
rect 445982 -2502 446066 -2266
rect 446302 -2502 485746 -2266
rect 485982 -2502 486066 -2266
rect 486302 -2502 525746 -2266
rect 525982 -2502 526066 -2266
rect 526302 -2502 565746 -2266
rect 565982 -2502 566066 -2266
rect 566302 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5746 -2586
rect 5982 -2822 6066 -2586
rect 6302 -2822 45746 -2586
rect 45982 -2822 46066 -2586
rect 46302 -2822 85746 -2586
rect 85982 -2822 86066 -2586
rect 86302 -2822 125746 -2586
rect 125982 -2822 126066 -2586
rect 126302 -2822 165746 -2586
rect 165982 -2822 166066 -2586
rect 166302 -2822 205746 -2586
rect 205982 -2822 206066 -2586
rect 206302 -2822 245746 -2586
rect 245982 -2822 246066 -2586
rect 246302 -2822 285746 -2586
rect 285982 -2822 286066 -2586
rect 286302 -2822 325746 -2586
rect 325982 -2822 326066 -2586
rect 326302 -2822 365746 -2586
rect 365982 -2822 366066 -2586
rect 366302 -2822 405746 -2586
rect 405982 -2822 406066 -2586
rect 406302 -2822 445746 -2586
rect 445982 -2822 446066 -2586
rect 446302 -2822 485746 -2586
rect 485982 -2822 486066 -2586
rect 486302 -2822 525746 -2586
rect 525982 -2822 526066 -2586
rect 526302 -2822 565746 -2586
rect 565982 -2822 566066 -2586
rect 566302 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 25746 -3226
rect 25982 -3462 26066 -3226
rect 26302 -3462 65746 -3226
rect 65982 -3462 66066 -3226
rect 66302 -3462 105746 -3226
rect 105982 -3462 106066 -3226
rect 106302 -3462 145746 -3226
rect 145982 -3462 146066 -3226
rect 146302 -3462 185746 -3226
rect 185982 -3462 186066 -3226
rect 186302 -3462 225746 -3226
rect 225982 -3462 226066 -3226
rect 226302 -3462 265746 -3226
rect 265982 -3462 266066 -3226
rect 266302 -3462 305746 -3226
rect 305982 -3462 306066 -3226
rect 306302 -3462 345746 -3226
rect 345982 -3462 346066 -3226
rect 346302 -3462 385746 -3226
rect 385982 -3462 386066 -3226
rect 386302 -3462 425746 -3226
rect 425982 -3462 426066 -3226
rect 426302 -3462 465746 -3226
rect 465982 -3462 466066 -3226
rect 466302 -3462 505746 -3226
rect 505982 -3462 506066 -3226
rect 506302 -3462 545746 -3226
rect 545982 -3462 546066 -3226
rect 546302 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 25746 -3546
rect 25982 -3782 26066 -3546
rect 26302 -3782 65746 -3546
rect 65982 -3782 66066 -3546
rect 66302 -3782 105746 -3546
rect 105982 -3782 106066 -3546
rect 106302 -3782 145746 -3546
rect 145982 -3782 146066 -3546
rect 146302 -3782 185746 -3546
rect 185982 -3782 186066 -3546
rect 186302 -3782 225746 -3546
rect 225982 -3782 226066 -3546
rect 226302 -3782 265746 -3546
rect 265982 -3782 266066 -3546
rect 266302 -3782 305746 -3546
rect 305982 -3782 306066 -3546
rect 306302 -3782 345746 -3546
rect 345982 -3782 346066 -3546
rect 346302 -3782 385746 -3546
rect 385982 -3782 386066 -3546
rect 386302 -3782 425746 -3546
rect 425982 -3782 426066 -3546
rect 426302 -3782 465746 -3546
rect 465982 -3782 466066 -3546
rect 466302 -3782 505746 -3546
rect 505982 -3782 506066 -3546
rect 506302 -3782 545746 -3546
rect 545982 -3782 546066 -3546
rect 546302 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9466 -4186
rect 9702 -4422 9786 -4186
rect 10022 -4422 49466 -4186
rect 49702 -4422 49786 -4186
rect 50022 -4422 89466 -4186
rect 89702 -4422 89786 -4186
rect 90022 -4422 129466 -4186
rect 129702 -4422 129786 -4186
rect 130022 -4422 169466 -4186
rect 169702 -4422 169786 -4186
rect 170022 -4422 209466 -4186
rect 209702 -4422 209786 -4186
rect 210022 -4422 249466 -4186
rect 249702 -4422 249786 -4186
rect 250022 -4422 289466 -4186
rect 289702 -4422 289786 -4186
rect 290022 -4422 329466 -4186
rect 329702 -4422 329786 -4186
rect 330022 -4422 369466 -4186
rect 369702 -4422 369786 -4186
rect 370022 -4422 409466 -4186
rect 409702 -4422 409786 -4186
rect 410022 -4422 449466 -4186
rect 449702 -4422 449786 -4186
rect 450022 -4422 489466 -4186
rect 489702 -4422 489786 -4186
rect 490022 -4422 529466 -4186
rect 529702 -4422 529786 -4186
rect 530022 -4422 569466 -4186
rect 569702 -4422 569786 -4186
rect 570022 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9466 -4506
rect 9702 -4742 9786 -4506
rect 10022 -4742 49466 -4506
rect 49702 -4742 49786 -4506
rect 50022 -4742 89466 -4506
rect 89702 -4742 89786 -4506
rect 90022 -4742 129466 -4506
rect 129702 -4742 129786 -4506
rect 130022 -4742 169466 -4506
rect 169702 -4742 169786 -4506
rect 170022 -4742 209466 -4506
rect 209702 -4742 209786 -4506
rect 210022 -4742 249466 -4506
rect 249702 -4742 249786 -4506
rect 250022 -4742 289466 -4506
rect 289702 -4742 289786 -4506
rect 290022 -4742 329466 -4506
rect 329702 -4742 329786 -4506
rect 330022 -4742 369466 -4506
rect 369702 -4742 369786 -4506
rect 370022 -4742 409466 -4506
rect 409702 -4742 409786 -4506
rect 410022 -4742 449466 -4506
rect 449702 -4742 449786 -4506
rect 450022 -4742 489466 -4506
rect 489702 -4742 489786 -4506
rect 490022 -4742 529466 -4506
rect 529702 -4742 529786 -4506
rect 530022 -4742 569466 -4506
rect 569702 -4742 569786 -4506
rect 570022 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 29466 -5146
rect 29702 -5382 29786 -5146
rect 30022 -5382 69466 -5146
rect 69702 -5382 69786 -5146
rect 70022 -5382 109466 -5146
rect 109702 -5382 109786 -5146
rect 110022 -5382 149466 -5146
rect 149702 -5382 149786 -5146
rect 150022 -5382 189466 -5146
rect 189702 -5382 189786 -5146
rect 190022 -5382 229466 -5146
rect 229702 -5382 229786 -5146
rect 230022 -5382 269466 -5146
rect 269702 -5382 269786 -5146
rect 270022 -5382 309466 -5146
rect 309702 -5382 309786 -5146
rect 310022 -5382 349466 -5146
rect 349702 -5382 349786 -5146
rect 350022 -5382 389466 -5146
rect 389702 -5382 389786 -5146
rect 390022 -5382 429466 -5146
rect 429702 -5382 429786 -5146
rect 430022 -5382 469466 -5146
rect 469702 -5382 469786 -5146
rect 470022 -5382 509466 -5146
rect 509702 -5382 509786 -5146
rect 510022 -5382 549466 -5146
rect 549702 -5382 549786 -5146
rect 550022 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 29466 -5466
rect 29702 -5702 29786 -5466
rect 30022 -5702 69466 -5466
rect 69702 -5702 69786 -5466
rect 70022 -5702 109466 -5466
rect 109702 -5702 109786 -5466
rect 110022 -5702 149466 -5466
rect 149702 -5702 149786 -5466
rect 150022 -5702 189466 -5466
rect 189702 -5702 189786 -5466
rect 190022 -5702 229466 -5466
rect 229702 -5702 229786 -5466
rect 230022 -5702 269466 -5466
rect 269702 -5702 269786 -5466
rect 270022 -5702 309466 -5466
rect 309702 -5702 309786 -5466
rect 310022 -5702 349466 -5466
rect 349702 -5702 349786 -5466
rect 350022 -5702 389466 -5466
rect 389702 -5702 389786 -5466
rect 390022 -5702 429466 -5466
rect 429702 -5702 429786 -5466
rect 430022 -5702 469466 -5466
rect 469702 -5702 469786 -5466
rect 470022 -5702 509466 -5466
rect 509702 -5702 509786 -5466
rect 510022 -5702 549466 -5466
rect 549702 -5702 549786 -5466
rect 550022 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 13186 -6106
rect 13422 -6342 13506 -6106
rect 13742 -6342 53186 -6106
rect 53422 -6342 53506 -6106
rect 53742 -6342 93186 -6106
rect 93422 -6342 93506 -6106
rect 93742 -6342 133186 -6106
rect 133422 -6342 133506 -6106
rect 133742 -6342 173186 -6106
rect 173422 -6342 173506 -6106
rect 173742 -6342 213186 -6106
rect 213422 -6342 213506 -6106
rect 213742 -6342 253186 -6106
rect 253422 -6342 253506 -6106
rect 253742 -6342 293186 -6106
rect 293422 -6342 293506 -6106
rect 293742 -6342 333186 -6106
rect 333422 -6342 333506 -6106
rect 333742 -6342 373186 -6106
rect 373422 -6342 373506 -6106
rect 373742 -6342 413186 -6106
rect 413422 -6342 413506 -6106
rect 413742 -6342 453186 -6106
rect 453422 -6342 453506 -6106
rect 453742 -6342 493186 -6106
rect 493422 -6342 493506 -6106
rect 493742 -6342 533186 -6106
rect 533422 -6342 533506 -6106
rect 533742 -6342 573186 -6106
rect 573422 -6342 573506 -6106
rect 573742 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 13186 -6426
rect 13422 -6662 13506 -6426
rect 13742 -6662 53186 -6426
rect 53422 -6662 53506 -6426
rect 53742 -6662 93186 -6426
rect 93422 -6662 93506 -6426
rect 93742 -6662 133186 -6426
rect 133422 -6662 133506 -6426
rect 133742 -6662 173186 -6426
rect 173422 -6662 173506 -6426
rect 173742 -6662 213186 -6426
rect 213422 -6662 213506 -6426
rect 213742 -6662 253186 -6426
rect 253422 -6662 253506 -6426
rect 253742 -6662 293186 -6426
rect 293422 -6662 293506 -6426
rect 293742 -6662 333186 -6426
rect 333422 -6662 333506 -6426
rect 333742 -6662 373186 -6426
rect 373422 -6662 373506 -6426
rect 373742 -6662 413186 -6426
rect 413422 -6662 413506 -6426
rect 413742 -6662 453186 -6426
rect 453422 -6662 453506 -6426
rect 453742 -6662 493186 -6426
rect 493422 -6662 493506 -6426
rect 493742 -6662 533186 -6426
rect 533422 -6662 533506 -6426
rect 533742 -6662 573186 -6426
rect 573422 -6662 573506 -6426
rect 573742 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33186 -7066
rect 33422 -7302 33506 -7066
rect 33742 -7302 73186 -7066
rect 73422 -7302 73506 -7066
rect 73742 -7302 113186 -7066
rect 113422 -7302 113506 -7066
rect 113742 -7302 153186 -7066
rect 153422 -7302 153506 -7066
rect 153742 -7302 193186 -7066
rect 193422 -7302 193506 -7066
rect 193742 -7302 233186 -7066
rect 233422 -7302 233506 -7066
rect 233742 -7302 273186 -7066
rect 273422 -7302 273506 -7066
rect 273742 -7302 313186 -7066
rect 313422 -7302 313506 -7066
rect 313742 -7302 353186 -7066
rect 353422 -7302 353506 -7066
rect 353742 -7302 393186 -7066
rect 393422 -7302 393506 -7066
rect 393742 -7302 433186 -7066
rect 433422 -7302 433506 -7066
rect 433742 -7302 473186 -7066
rect 473422 -7302 473506 -7066
rect 473742 -7302 513186 -7066
rect 513422 -7302 513506 -7066
rect 513742 -7302 553186 -7066
rect 553422 -7302 553506 -7066
rect 553742 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33186 -7386
rect 33422 -7622 33506 -7386
rect 33742 -7622 73186 -7386
rect 73422 -7622 73506 -7386
rect 73742 -7622 113186 -7386
rect 113422 -7622 113506 -7386
rect 113742 -7622 153186 -7386
rect 153422 -7622 153506 -7386
rect 153742 -7622 193186 -7386
rect 193422 -7622 193506 -7386
rect 193742 -7622 233186 -7386
rect 233422 -7622 233506 -7386
rect 233742 -7622 273186 -7386
rect 273422 -7622 273506 -7386
rect 273742 -7622 313186 -7386
rect 313422 -7622 313506 -7386
rect 313742 -7622 353186 -7386
rect 353422 -7622 353506 -7386
rect 353742 -7622 393186 -7386
rect 393422 -7622 393506 -7386
rect 393742 -7622 433186 -7386
rect 433422 -7622 433506 -7386
rect 433742 -7622 473186 -7386
rect 473422 -7622 473506 -7386
rect 473742 -7622 513186 -7386
rect 513422 -7622 513506 -7386
rect 513742 -7622 553186 -7386
rect 553422 -7622 553506 -7386
rect 553742 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_proj_example  mprj
timestamp 0
transform 1 0 4000 0 1 4000
box 0 0 571964 694008
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 3066 586890 3686 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 43066 586890 43686 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 83066 586890 83686 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 123066 586890 123686 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 163066 586890 163686 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 203066 586890 203686 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 243066 586890 243686 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 283066 586890 283686 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 323066 586890 323686 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 363066 586890 363686 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 403066 586890 403686 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 443066 586890 443686 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 483066 586890 483686 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 523066 586890 523686 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 563066 586890 563686 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 603066 586890 603686 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 643066 586890 643686 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 683066 586890 683686 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1994 -1894 2614 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 41994 -1894 42614 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 81994 -1894 82614 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 121994 -1894 122614 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 161994 -1894 162614 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 201994 -1894 202614 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 241994 -1894 242614 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 281994 -1894 282614 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 321994 -1894 322614 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361994 -1894 362614 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 401994 -1894 402614 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 441994 -1894 442614 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 481994 -1894 482614 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 521994 -1894 522614 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 561994 -1894 562614 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1994 700008 2614 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 41994 700008 42614 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 81994 700008 82614 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 121994 700008 122614 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 161994 700008 162614 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 201994 700008 202614 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 241994 700008 242614 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 281994 700008 282614 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 321994 700008 322614 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361994 700008 362614 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 401994 700008 402614 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 441994 700008 442614 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 481994 700008 482614 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 521994 700008 522614 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 561994 700008 562614 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6786 588810 7406 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 46786 588810 47406 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 86786 588810 87406 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 126786 588810 127406 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 166786 588810 167406 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 206786 588810 207406 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 246786 588810 247406 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 286786 588810 287406 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 326786 588810 327406 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366786 588810 367406 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 406786 588810 407406 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 446786 588810 447406 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 486786 588810 487406 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 526786 588810 527406 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 566786 588810 567406 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 606786 588810 607406 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 646786 588810 647406 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 686786 588810 687406 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5714 -3814 6334 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 45714 -3814 46334 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 85714 -3814 86334 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 125714 -3814 126334 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 165714 -3814 166334 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 205714 -3814 206334 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 245714 -3814 246334 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 285714 -3814 286334 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 325714 -3814 326334 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 365714 -3814 366334 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 405714 -3814 406334 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 445714 -3814 446334 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 485714 -3814 486334 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 525714 -3814 526334 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 565714 -3814 566334 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5714 700008 6334 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 45714 700008 46334 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 85714 700008 86334 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 125714 700008 126334 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 165714 700008 166334 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 205714 700008 206334 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 245714 700008 246334 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 285714 700008 286334 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 325714 700008 326334 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365714 700008 366334 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 405714 700008 406334 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 445714 700008 446334 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 485714 700008 486334 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 525714 700008 526334 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 565714 700008 566334 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10506 590730 11126 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 50506 590730 51126 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 90506 590730 91126 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 130506 590730 131126 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 170506 590730 171126 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 210506 590730 211126 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 250506 590730 251126 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 290506 590730 291126 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 330506 590730 331126 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370506 590730 371126 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 410506 590730 411126 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 450506 590730 451126 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 490506 590730 491126 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 530506 590730 531126 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 570506 590730 571126 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 610506 590730 611126 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 650506 590730 651126 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 690506 590730 691126 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9434 -5734 10054 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 49434 -5734 50054 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 89434 -5734 90054 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 129434 -5734 130054 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 169434 -5734 170054 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 209434 -5734 210054 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 249434 -5734 250054 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 289434 -5734 290054 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 329434 -5734 330054 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 369434 -5734 370054 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 409434 -5734 410054 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 449434 -5734 450054 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 489434 -5734 490054 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 529434 -5734 530054 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 569434 -5734 570054 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9434 700008 10054 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 49434 700008 50054 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 89434 700008 90054 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 129434 700008 130054 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 169434 700008 170054 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 209434 700008 210054 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 249434 700008 250054 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 289434 700008 290054 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 329434 700008 330054 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369434 700008 370054 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 409434 700008 410054 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 449434 700008 450054 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 489434 700008 490054 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 529434 700008 530054 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 569434 700008 570054 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14226 592650 14846 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 54226 592650 54846 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 94226 592650 94846 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 134226 592650 134846 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 174226 592650 174846 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 214226 592650 214846 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 254226 592650 254846 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 294226 592650 294846 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 334226 592650 334846 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374226 592650 374846 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 414226 592650 414846 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 454226 592650 454846 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 494226 592650 494846 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 534226 592650 534846 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 574226 592650 574846 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 614226 592650 614846 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 654226 592650 654846 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 694226 592650 694846 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 13154 -7654 13774 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 53154 -7654 53774 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 93154 -7654 93774 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 133154 -7654 133774 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 173154 -7654 173774 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 213154 -7654 213774 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 253154 -7654 253774 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 293154 -7654 293774 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 333154 -7654 333774 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 373154 -7654 373774 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 413154 -7654 413774 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 453154 -7654 453774 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 493154 -7654 493774 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 533154 -7654 533774 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 573154 -7654 573774 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 13154 700008 13774 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 53154 700008 53774 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 93154 700008 93774 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 133154 700008 133774 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 173154 700008 173774 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 213154 700008 213774 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 253154 700008 253774 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 293154 700008 293774 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 333154 700008 333774 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 373154 700008 373774 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 413154 700008 413774 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 453154 700008 453774 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 493154 700008 493774 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 533154 700008 533774 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 573154 700008 573774 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 30506 590730 31126 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 70506 590730 71126 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 110506 590730 111126 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 150506 590730 151126 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 190506 590730 191126 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 230506 590730 231126 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 270506 590730 271126 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 310506 590730 311126 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 350506 590730 351126 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 390506 590730 391126 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 430506 590730 431126 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 470506 590730 471126 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 510506 590730 511126 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 550506 590730 551126 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 590506 590730 591126 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 630506 590730 631126 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 670506 590730 671126 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 29434 -5734 30054 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 69434 -5734 70054 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 109434 -5734 110054 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 149434 -5734 150054 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 189434 -5734 190054 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 229434 -5734 230054 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 269434 -5734 270054 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 309434 -5734 310054 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 349434 -5734 350054 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 389434 -5734 390054 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 429434 -5734 430054 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 469434 -5734 470054 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 509434 -5734 510054 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 549434 -5734 550054 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 29434 700008 30054 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 69434 700008 70054 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 109434 700008 110054 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 149434 700008 150054 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 189434 700008 190054 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 229434 700008 230054 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 269434 700008 270054 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 309434 700008 310054 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 349434 700008 350054 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 389434 700008 390054 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 429434 700008 430054 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 469434 700008 470054 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 509434 700008 510054 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 549434 700008 550054 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 34226 592650 34846 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 74226 592650 74846 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 114226 592650 114846 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 154226 592650 154846 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 194226 592650 194846 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 234226 592650 234846 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 274226 592650 274846 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 314226 592650 314846 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 354226 592650 354846 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 394226 592650 394846 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 434226 592650 434846 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 474226 592650 474846 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 514226 592650 514846 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 554226 592650 554846 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 594226 592650 594846 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 634226 592650 634846 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 674226 592650 674846 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 33154 -7654 33774 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 73154 -7654 73774 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 113154 -7654 113774 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 153154 -7654 153774 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 193154 -7654 193774 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 233154 -7654 233774 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 273154 -7654 273774 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 313154 -7654 313774 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 353154 -7654 353774 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 393154 -7654 393774 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 433154 -7654 433774 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 473154 -7654 473774 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 513154 -7654 513774 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 553154 -7654 553774 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 33154 700008 33774 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 73154 700008 73774 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 113154 700008 113774 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 153154 700008 153774 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 193154 700008 193774 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 233154 700008 233774 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 273154 700008 273774 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 313154 700008 313774 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 353154 700008 353774 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 393154 700008 393774 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 433154 700008 433774 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 473154 700008 473774 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 513154 700008 513774 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 553154 700008 553774 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 23066 586890 23686 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 63066 586890 63686 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 103066 586890 103686 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 143066 586890 143686 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 183066 586890 183686 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 223066 586890 223686 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 263066 586890 263686 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 303066 586890 303686 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 343066 586890 343686 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 383066 586890 383686 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 423066 586890 423686 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 463066 586890 463686 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 503066 586890 503686 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 543066 586890 543686 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 583066 586890 583686 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 623066 586890 623686 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 663066 586890 663686 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 21994 -1894 22614 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 61994 -1894 62614 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 101994 -1894 102614 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 141994 -1894 142614 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 181994 -1894 182614 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 221994 -1894 222614 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 261994 -1894 262614 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 301994 -1894 302614 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 341994 -1894 342614 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 381994 -1894 382614 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 421994 -1894 422614 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 461994 -1894 462614 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 501994 -1894 502614 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 541994 -1894 542614 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 21994 700008 22614 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 61994 700008 62614 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 101994 700008 102614 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 141994 700008 142614 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 181994 700008 182614 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 221994 700008 222614 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 261994 700008 262614 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 301994 700008 302614 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 341994 700008 342614 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 381994 700008 382614 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 421994 700008 422614 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 461994 700008 462614 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 501994 700008 502614 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 541994 700008 542614 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 26786 588810 27406 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 66786 588810 67406 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 106786 588810 107406 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 146786 588810 147406 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 186786 588810 187406 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 226786 588810 227406 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 266786 588810 267406 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 306786 588810 307406 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 346786 588810 347406 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 386786 588810 387406 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 426786 588810 427406 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 466786 588810 467406 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 506786 588810 507406 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 546786 588810 547406 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 586786 588810 587406 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 626786 588810 627406 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 666786 588810 667406 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 25714 -3814 26334 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 65714 -3814 66334 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 105714 -3814 106334 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 145714 -3814 146334 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 185714 -3814 186334 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 225714 -3814 226334 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 265714 -3814 266334 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 305714 -3814 306334 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 345714 -3814 346334 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 385714 -3814 386334 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 425714 -3814 426334 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 465714 -3814 466334 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 505714 -3814 506334 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 545714 -3814 546334 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 25714 700008 26334 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 65714 700008 66334 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 105714 700008 106334 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 145714 700008 146334 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 185714 700008 186334 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 225714 700008 226334 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 265714 700008 266334 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 305714 700008 306334 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 345714 700008 346334 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 385714 700008 386334 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 425714 700008 426334 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 465714 700008 466334 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 505714 700008 506334 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 545714 700008 546334 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
